magic
tech sky130A
magscale 1 2
timestamp 1696522064
<< metal1 >>
rect 10830 20044 11030 20046
rect 10830 19846 11634 20044
rect 12710 19832 13632 20026
rect 14684 19974 15582 20016
rect 14684 19862 14968 19974
rect 15100 19862 15582 19974
rect 14684 19814 15582 19862
rect 25932 11604 26514 11606
rect 25868 11404 26514 11604
rect 25932 11402 26514 11404
rect 7812 6804 8012 6826
rect 7812 6650 7832 6804
rect 7992 6650 8012 6804
rect 7812 6626 8012 6650
rect 39776 5826 39976 6026
<< via1 >>
rect 14968 19862 15100 19974
rect 16658 19842 16786 19978
rect 7832 6650 7992 6804
<< metal2 >>
rect 14926 19988 15148 20006
rect 14926 19850 14946 19988
rect 15118 19850 15148 19988
rect 14926 19836 15148 19850
rect 16642 19980 16798 19988
rect 16642 19840 16654 19980
rect 16786 19840 16798 19980
rect 16642 19830 16798 19840
rect 7774 6836 8046 6856
rect 7774 6614 7800 6836
rect 8024 6614 8046 6836
rect 7774 6598 8046 6614
<< via2 >>
rect 14946 19974 15118 19988
rect 14946 19862 14968 19974
rect 14968 19862 15100 19974
rect 15100 19862 15118 19974
rect 14946 19850 15118 19862
rect 16654 19978 16786 19980
rect 16654 19842 16658 19978
rect 16658 19842 16786 19978
rect 16654 19840 16786 19842
rect 22378 17494 22560 17662
rect 26816 17436 27132 17736
rect 33716 17482 33844 17620
rect 35284 17486 35462 17638
rect 39800 17508 39966 17676
rect 30800 9584 30918 9698
rect 7800 6804 8024 6836
rect 7800 6650 7832 6804
rect 7832 6650 7992 6804
rect 7992 6650 8024 6804
rect 7800 6614 8024 6650
rect 12458 6600 12712 6860
<< metal3 >>
rect 14886 21134 35636 21536
rect 14896 19988 15170 21134
rect 14896 19850 14946 19988
rect 15118 19850 15170 19988
rect 14896 18414 15170 19850
rect 16626 19980 22636 20010
rect 16626 19840 16654 19980
rect 16786 19840 22636 19980
rect 16626 19802 22636 19840
rect 7660 18158 15170 18414
rect 7660 18156 15128 18158
rect 7662 8644 8016 18156
rect 22308 17662 22636 19802
rect 22308 17494 22378 17662
rect 22560 17494 22636 17662
rect 22308 17474 22636 17494
rect 26768 17756 27182 17794
rect 26768 17406 26798 17756
rect 27148 17406 27182 17756
rect 35170 17638 35636 21134
rect 33706 17622 33856 17628
rect 33706 17482 33710 17622
rect 33850 17482 33856 17622
rect 33706 17476 33856 17482
rect 35170 17486 35284 17638
rect 35462 17486 35636 17638
rect 26768 17376 27182 17406
rect 35170 17382 35636 17486
rect 39756 17706 40018 17728
rect 39756 17470 39774 17706
rect 40004 17470 40018 17706
rect 39756 17456 40018 17470
rect 30790 9698 30940 9716
rect 30790 9584 30800 9698
rect 30918 9584 30940 9698
rect 30790 9574 30940 9584
rect 7662 8080 12896 8644
rect 7722 6860 12734 6902
rect 7722 6836 12458 6860
rect 7722 6614 7800 6836
rect 8024 6614 12458 6836
rect 7722 6600 12458 6614
rect 12712 6600 12734 6860
rect 7722 6538 12734 6600
<< via3 >>
rect 26798 17736 27148 17756
rect 26798 17436 26816 17736
rect 26816 17436 27132 17736
rect 27132 17436 27148 17736
rect 26798 17406 27148 17436
rect 33710 17620 33850 17622
rect 33710 17482 33716 17620
rect 33716 17482 33844 17620
rect 33844 17482 33850 17620
rect 39774 17676 40004 17706
rect 39774 17508 39800 17676
rect 39800 17508 39966 17676
rect 39966 17508 40004 17676
rect 39774 17470 40004 17508
rect 30806 9590 30912 9692
<< metal4 >>
rect 26712 22328 27238 22358
rect 26708 22326 44074 22328
rect 26708 22024 44078 22326
rect 26712 17756 27238 22024
rect 20584 12966 21098 17736
rect 26712 17406 26798 17756
rect 27148 17406 27238 17756
rect 39654 17706 40104 17794
rect 26712 17328 27238 17406
rect 33678 17622 33890 17672
rect 33678 17482 33710 17622
rect 33850 17482 33890 17622
rect 12386 12638 21098 12966
rect 20584 10572 21098 12638
rect 24732 13026 25104 13034
rect 33678 13026 33890 17482
rect 24732 12636 33890 13026
rect 24732 12630 25104 12636
rect 33678 12634 33890 12636
rect 39654 17470 39774 17706
rect 40004 17470 40104 17706
rect 24730 10080 25104 12630
rect 39654 11626 40104 17470
rect 43562 11626 44078 22024
rect 39646 11068 44080 11626
rect 24162 9900 31140 10080
rect 24730 9884 25104 9900
rect 30988 9732 31140 9900
rect 30776 9692 31142 9732
rect 30776 9590 30806 9692
rect 30912 9590 31142 9692
rect 30776 9554 31142 9590
rect 39654 6080 40104 11068
rect 35866 5752 40110 6080
use opamp  x1
timestamp 1696521366
transform 1 0 19232 0 1 3428
box 6068 1244 19288 9014
use switch  x2
timestamp 1696147897
transform 0 1 32036 -1 0 21894
box -53 -918 8642 11418
use switch  x3
timestamp 1696147897
transform 0 1 19130 -1 0 21904
box -53 -918 8642 11418
use switch  x4
timestamp 1696147897
transform 1 0 8253 0 1 4996
box -53 -918 8642 11418
use not  x5
timestamp 1696147843
transform 1 0 10958 0 1 19770
box 476 -578 1868 990
use not  x6
timestamp 1696147843
transform 1 0 12976 0 1 19752
box 476 -578 1868 990
use not  x7
timestamp 1696147843
transform 1 0 14944 0 1 19742
box 476 -578 1868 990
use sky130_fd_pr__cap_mim_m3_1_3HBNLG  XC1
timestamp 1695395215
transform 1 0 21062 0 1 8034
box -3186 -3040 3186 3040
<< labels >>
flabel metal1 10830 19846 11030 20046 0 FreeSans 256 0 0 0 sw1
port 0 nsew
flabel metal1 39776 5826 39976 6026 0 FreeSans 256 0 0 0 shout
port 3 nsew
flabel metal1 25868 11404 26068 11604 0 FreeSans 256 0 0 0 opbias
port 1 nsew
flabel metal1 7812 6626 8012 6826 0 FreeSans 256 0 0 0 shin
port 2 nsew
<< end >>
