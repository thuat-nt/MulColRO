magic
tech sky130A
magscale 1 2
timestamp 1695461917
<< error_p >>
rect 167104 617048 167106 617098
rect 167132 617048 167134 617126
rect 166552 616808 167190 617048
rect 172318 617004 172320 617082
rect 172346 617004 172348 617054
rect 172262 616764 172900 617004
rect 167086 616502 167106 616622
rect 167114 616496 167134 616650
rect 172318 616452 172338 616606
rect 172346 616458 172366 616578
rect 189325 616416 189359 619559
rect 192071 613502 192105 619460
rect 192843 616416 192877 619559
rect 194396 616416 194430 619564
rect 197914 616416 197948 617020
rect 189325 613195 189359 613502
rect 189439 613291 189473 613325
rect 190097 613291 190131 613325
rect 190755 613291 190789 613325
rect 191413 613291 191447 613325
rect 192071 613291 192105 613325
rect 192729 613291 192783 613325
rect 189389 613257 189393 613291
rect 189405 613257 192783 613291
rect 120502 610080 120504 610130
rect 120530 610080 120532 610158
rect 119950 609840 120588 610080
rect 125716 610036 125718 610114
rect 125744 610036 125746 610086
rect 125660 609796 126298 610036
rect 120484 609534 120504 609654
rect 120512 609528 120532 609682
rect 125716 609484 125736 609638
rect 125744 609490 125764 609610
rect 112980 603945 113014 608884
rect 116416 608866 117898 608978
rect 114976 608832 121142 608866
rect 116416 608208 117898 608832
rect 114976 608174 121142 608208
rect 116416 607550 117898 608174
rect 119950 607550 120588 607648
rect 120638 607562 121186 607590
rect 120638 607556 121154 607562
rect 120638 607550 120672 607556
rect 114976 607522 121146 607550
rect 121152 607535 121154 607556
rect 121175 607551 121186 607562
rect 114976 607516 121142 607522
rect 116416 607402 117898 607516
rect 119950 607186 120588 607516
rect 120638 607274 120672 607516
rect 121000 607476 121011 607487
rect 120702 607432 120774 607470
rect 120824 607460 121011 607476
rect 121012 607460 121084 607470
rect 120812 607436 121084 607460
rect 121012 607432 121084 607436
rect 120740 607398 120774 607432
rect 120784 607408 121040 607432
rect 121000 607388 121011 607399
rect 121050 607398 121084 607432
rect 120824 607354 121011 607388
rect 121152 607274 121186 607535
rect 120638 607240 121186 607274
rect 119950 606914 120588 607172
rect 119798 606892 120588 606914
rect 114976 606858 120588 606892
rect 119798 606840 120588 606858
rect 119950 606710 120588 606840
rect 120638 607080 121186 607114
rect 120638 606892 120672 607080
rect 120702 606956 120774 606994
rect 120778 606984 120810 607004
rect 121000 607000 121011 607011
rect 120778 606956 120782 606976
rect 120824 606966 121011 607000
rect 121012 606956 121084 606994
rect 120740 606906 120774 606956
rect 121000 606912 121011 606923
rect 120824 606904 121011 606912
rect 121050 606906 121084 606956
rect 120824 606892 121000 606904
rect 121152 606893 121186 607080
rect 121192 606998 121226 607488
rect 121294 606998 121328 608884
rect 121192 606920 121328 606998
rect 120638 606858 121142 606892
rect 121152 606877 121176 606893
rect 121152 606870 121186 606877
rect 120638 606798 120672 606858
rect 121152 606854 121260 606870
rect 121152 606842 121186 606854
rect 121152 606826 121232 606842
rect 121152 606798 121186 606826
rect 120638 606764 121186 606798
rect 121192 606522 121226 606826
rect 121294 606522 121328 606920
rect 121192 606436 121328 606522
rect 121192 606326 121226 606436
rect 113055 606315 121253 606326
rect 113066 606303 121242 606315
rect 113055 606292 121253 606303
rect 113082 606246 113116 606292
rect 114096 606246 114554 606266
rect 121192 606262 121226 606292
rect 114096 606234 114594 606246
rect 113166 606188 121142 606234
rect 113166 606178 121153 606188
rect 114096 606174 114594 606178
rect 113082 605582 113116 606172
rect 114136 606154 114594 606174
rect 113746 606130 114850 606150
rect 113718 606102 114878 606122
rect 117006 605970 117454 605998
rect 117006 605786 117472 605970
rect 117024 605758 117472 605786
rect 119770 605587 120424 605600
rect 116120 605576 118252 605587
rect 118870 605576 121153 605587
rect 121192 605582 121226 606172
rect 113166 605566 121153 605576
rect 113166 605520 121142 605566
rect 119806 605502 120460 605520
rect 113082 605492 113116 605496
rect 121192 605492 121226 605496
rect 113035 605428 121273 605462
rect 121294 605350 121328 606436
rect 124920 606954 124954 608840
rect 125062 607512 125610 607546
rect 125022 606954 125056 607444
rect 125062 607230 125096 607512
rect 125576 607506 125610 607512
rect 125102 607478 125610 607506
rect 125106 607472 125130 607478
rect 125542 607472 125610 607478
rect 125424 607432 125435 607443
rect 125126 607388 125198 607426
rect 125248 607416 125435 607432
rect 125436 607416 125508 607426
rect 125236 607392 125508 607416
rect 125436 607388 125508 607392
rect 125164 607354 125198 607388
rect 125208 607364 125464 607388
rect 125424 607344 125435 607355
rect 125474 607354 125508 607388
rect 125248 607310 125435 607344
rect 125576 607230 125610 607472
rect 125062 607196 125610 607230
rect 125660 607142 126298 607604
rect 124920 606876 125056 606954
rect 125062 607036 125610 607070
rect 124920 606478 124954 606876
rect 125062 606826 125096 607036
rect 125424 606956 125435 606967
rect 125126 606912 125198 606950
rect 125248 606922 125435 606956
rect 125438 606950 125470 606960
rect 125436 606912 125508 606950
rect 125164 606888 125198 606912
rect 125474 606888 125508 606912
rect 125164 606878 125236 606888
rect 125237 606868 125435 606879
rect 125474 606878 125546 606888
rect 125248 606860 125435 606868
rect 125248 606848 125424 606860
rect 125576 606848 125610 607036
rect 124988 606810 125096 606826
rect 125106 606814 125610 606848
rect 125062 606798 125096 606810
rect 125016 606782 125096 606798
rect 125022 606478 125056 606782
rect 125062 606754 125096 606782
rect 125576 606754 125610 606814
rect 125062 606720 125610 606754
rect 125660 606870 126298 607128
rect 125660 606848 126450 606870
rect 125660 606814 133082 606848
rect 125660 606796 126450 606814
rect 125660 606666 126298 606796
rect 124920 606392 125056 606478
rect 124920 605404 124954 606392
rect 125022 606282 125056 606392
rect 131634 606282 131690 606304
rect 124995 606271 133193 606282
rect 125006 606259 133182 606271
rect 124995 606248 133193 606259
rect 125022 606218 125056 606248
rect 131694 606202 132152 606222
rect 131658 606190 132152 606202
rect 125106 606144 133082 606190
rect 125106 606134 133093 606144
rect 131658 606130 132152 606134
rect 125022 605538 125056 606128
rect 131658 606110 132112 606130
rect 131634 606086 132502 606106
rect 130622 606072 130678 606078
rect 131634 606058 132530 606078
rect 131634 606030 131690 606058
rect 128794 605926 129242 605954
rect 128776 605742 129242 605926
rect 128776 605714 129224 605742
rect 125824 605543 126478 605556
rect 125095 605532 133093 605543
rect 133132 605538 133166 606128
rect 125106 605522 133093 605532
rect 125106 605476 133082 605522
rect 125788 605458 126442 605476
rect 125022 605448 125056 605452
rect 133132 605448 133166 605452
rect 124975 605404 133213 605418
rect 133234 605404 133268 608840
rect 124920 605384 133268 605404
rect 124920 605350 124954 605384
rect 133234 605350 133268 605384
rect 117012 605114 117460 605326
rect 118844 605316 135136 605350
rect 116474 604550 117112 605012
rect 117162 604924 117710 604958
rect 117162 604896 117196 604924
rect 117676 604896 117710 604924
rect 118844 604896 118878 605316
rect 119688 605248 119726 605286
rect 120446 605248 120484 605286
rect 121192 605248 121226 605316
rect 121236 605264 121242 605306
rect 119020 605214 119726 605248
rect 119778 605214 120484 605248
rect 120536 605214 121226 605248
rect 121153 605176 121154 605177
rect 121192 605176 121226 605214
rect 121278 605204 121284 605264
rect 121294 605214 121328 605316
rect 121290 605204 121328 605214
rect 121250 605180 121328 605204
rect 121232 605178 121328 605180
rect 121232 605176 121266 605178
rect 121278 605176 121284 605178
rect 121154 605175 121155 605176
rect 118947 605164 118992 605175
rect 119705 605164 119750 605175
rect 120463 605164 120508 605175
rect 118958 604896 118992 605164
rect 119003 604908 119004 604909
rect 119704 604908 119705 604909
rect 119004 604907 119005 604908
rect 119703 604907 119704 604908
rect 119716 604896 119750 605164
rect 119761 604908 119762 604909
rect 120462 604908 120463 604909
rect 119762 604907 119763 604908
rect 120461 604907 120462 604908
rect 120474 604896 120508 605164
rect 121192 605150 121272 605176
rect 121192 604924 121266 605150
rect 120519 604908 120520 604909
rect 121198 604908 121266 604924
rect 120520 604907 120521 604908
rect 121142 604896 121153 604907
rect 117162 604862 117230 604896
rect 117310 604878 117562 604882
rect 117308 604862 117564 604878
rect 117162 604858 117196 604862
rect 117308 604858 117340 604862
rect 117162 604856 117340 604858
rect 117534 604856 117564 604862
rect 117676 604862 117744 604896
rect 118810 604862 121153 604896
rect 117162 604642 117196 604856
rect 117336 604844 117536 604850
rect 117336 604838 117340 604844
rect 117226 604830 117340 604838
rect 117212 604828 117340 604830
rect 117348 604838 117536 604844
rect 117348 604828 117646 604838
rect 117226 604806 117336 604828
rect 117348 604810 117535 604828
rect 117536 604806 117646 604828
rect 117226 604804 117646 604806
rect 117226 604800 117336 604804
rect 117536 604800 117646 604804
rect 117264 604778 117336 604800
rect 117264 604776 117564 604778
rect 117264 604766 117336 604776
rect 117337 604756 117535 604767
rect 117574 604766 117646 604800
rect 117348 604722 117535 604756
rect 117676 604642 117710 604862
rect 117162 604608 117710 604642
rect 118844 604238 118878 604862
rect 118958 604238 118992 604862
rect 119004 604850 119005 604851
rect 119703 604850 119704 604851
rect 119003 604849 119004 604850
rect 119704 604849 119705 604850
rect 119003 604250 119004 604251
rect 119704 604250 119705 604251
rect 119004 604249 119005 604250
rect 119703 604249 119704 604250
rect 119716 604238 119750 604862
rect 119762 604850 119763 604851
rect 120461 604850 120462 604851
rect 119761 604849 119762 604850
rect 120462 604849 120463 604850
rect 119786 604260 119790 604272
rect 119761 604250 119762 604251
rect 119762 604249 119763 604250
rect 119798 604238 119802 604260
rect 120462 604250 120463 604251
rect 120461 604249 120462 604250
rect 120474 604238 120508 604862
rect 120520 604850 120521 604851
rect 121154 604850 121226 604872
rect 121232 604850 121266 604908
rect 120519 604849 120520 604850
rect 121154 604834 121266 604850
rect 121192 604266 121266 604834
rect 120519 604250 120520 604251
rect 121198 604250 121266 604266
rect 120520 604249 120521 604250
rect 121142 604238 121153 604249
rect 118810 604204 121153 604238
rect 117078 604010 117210 604128
rect 117010 603945 117458 604010
rect 118844 603945 118878 604204
rect 118958 603945 118992 604204
rect 119004 604192 119005 604193
rect 119703 604192 119704 604193
rect 119003 604191 119004 604192
rect 119704 604191 119705 604192
rect 119608 604162 119668 604176
rect 119716 603945 119750 604204
rect 119762 604192 119763 604193
rect 120461 604192 120462 604193
rect 119761 604191 119762 604192
rect 120462 604191 120463 604192
rect 119792 604162 119854 604176
rect 120358 604162 120468 604176
rect 120474 603945 120508 604204
rect 120520 604192 120521 604193
rect 121154 604192 121226 604214
rect 121232 604192 121266 604250
rect 120519 604191 120520 604192
rect 121154 604176 121266 604192
rect 120514 604162 120624 604176
rect 121192 603945 121266 604176
rect 121290 603945 121328 605178
rect 112949 602738 121387 603945
rect 112985 600042 113019 602738
rect 118808 602485 121387 602738
rect 113168 602466 113468 602485
rect 114820 602466 116320 602485
rect 117888 602468 121387 602485
rect 118460 602368 118472 602434
rect 118702 602356 118718 602434
rect 113412 602340 114876 602356
rect 116510 602288 117076 602322
rect 116510 601966 116544 602288
rect 117042 602224 117076 602288
rect 117126 602224 117746 602340
rect 116694 602208 116892 602219
rect 116565 602146 116693 602193
rect 116705 602174 116892 602208
rect 116978 602193 117746 602224
rect 116893 602146 117746 602193
rect 116612 602108 116693 602146
rect 116940 602108 117746 602146
rect 116694 602080 116892 602091
rect 116950 602082 117746 602108
rect 116705 602046 116892 602080
rect 116978 602012 117746 602082
rect 117042 601966 117076 602012
rect 116510 601932 117076 601966
rect 117126 601918 117746 602012
rect 116986 601366 117434 601578
rect 117078 601356 117210 601366
rect 118808 601255 121387 602468
rect 113060 601244 121387 601255
rect 113071 601232 121387 601244
rect 113060 601221 121387 601232
rect 113087 601175 113121 601221
rect 113996 601163 114452 601182
rect 118808 601163 121387 601221
rect 113180 601107 121387 601163
rect 113087 600511 113121 601101
rect 114034 601092 114490 601107
rect 116986 600902 117434 600912
rect 116978 600700 117434 600902
rect 116978 600690 117426 600700
rect 116120 600505 118252 600516
rect 118808 600505 121387 601107
rect 121990 600616 122024 605164
rect 124264 600616 124298 605164
rect 124920 603901 124954 605316
rect 128326 605312 128612 605316
rect 125022 605282 125032 605286
rect 125046 605282 125056 605286
rect 124984 605214 125010 605248
rect 125022 605180 125056 605282
rect 125752 605248 125790 605286
rect 126510 605248 126548 605286
rect 127268 605248 127306 605286
rect 128026 605248 128064 605286
rect 128360 605248 128578 605298
rect 128784 605282 128822 605286
rect 128784 605248 129236 605282
rect 129542 605248 129580 605286
rect 129706 605248 129928 605286
rect 130300 605248 130338 605286
rect 131058 605248 131096 605286
rect 131816 605248 131854 605286
rect 132574 605248 132612 605286
rect 133132 605248 133166 605316
rect 133234 605248 133268 605316
rect 125068 605214 125790 605248
rect 125842 605214 126548 605248
rect 126600 605214 127306 605248
rect 127358 605214 128064 605248
rect 128116 605214 129580 605248
rect 129632 605214 130338 605248
rect 130390 605214 131096 605248
rect 131148 605214 131854 605248
rect 131906 605214 132612 605248
rect 132664 605214 133268 605248
rect 125022 605176 125032 605180
rect 125046 605176 125056 605180
rect 125094 605176 125095 605177
rect 125010 604864 125068 605176
rect 125093 605175 125094 605176
rect 125769 605164 125814 605175
rect 126527 605164 126572 605175
rect 127285 605164 127330 605175
rect 128043 605164 128088 605175
rect 125768 604864 125769 604865
rect 125767 604863 125768 604864
rect 125780 604852 125814 605164
rect 125825 604864 125826 604865
rect 126526 604864 126527 604865
rect 125826 604863 125827 604864
rect 126525 604863 126526 604864
rect 126538 604852 126572 605164
rect 126583 604864 126584 604865
rect 127284 604864 127285 604865
rect 126584 604863 126585 604864
rect 127283 604863 127284 604864
rect 127296 604852 127330 605164
rect 127341 604864 127342 604865
rect 128042 604864 128043 604865
rect 127342 604863 127343 604864
rect 128041 604863 128042 604864
rect 128054 604852 128088 605164
rect 128788 605070 129236 605214
rect 133093 605176 133094 605177
rect 133094 605175 133095 605176
rect 129559 605164 129604 605175
rect 130317 605164 130362 605175
rect 131075 605164 131120 605175
rect 131833 605164 131878 605175
rect 132591 605164 132636 605175
rect 128686 604914 128712 604950
rect 128714 604914 128740 604950
rect 128812 604914 128846 605070
rect 129570 604968 129604 605164
rect 128538 604880 129086 604914
rect 128099 604864 128100 604865
rect 128100 604863 128101 604864
rect 128538 604863 128572 604880
rect 128360 604852 128578 604863
rect 128686 604858 128712 604880
rect 128714 604858 128740 604880
rect 128800 604864 128801 604865
rect 128799 604863 128800 604864
rect 128812 604852 128846 604880
rect 128857 604864 128858 604865
rect 128858 604863 128859 604864
rect 129052 604852 129086 604880
rect 129136 604863 129774 604968
rect 130316 604864 130317 604865
rect 130315 604863 130316 604864
rect 129136 604852 129928 604863
rect 130328 604852 130362 605164
rect 130373 604864 130374 604865
rect 131074 604864 131075 604865
rect 130374 604863 130375 604864
rect 131073 604863 131074 604864
rect 131086 604852 131120 605164
rect 131131 604864 131132 604865
rect 131832 604864 131833 604865
rect 131132 604863 131133 604864
rect 131831 604863 131832 604864
rect 131844 604852 131878 605164
rect 131889 604864 131890 604865
rect 132590 604864 132591 604865
rect 131890 604863 131891 604864
rect 132589 604863 132590 604864
rect 132602 604852 132636 605164
rect 133132 604880 133166 605214
rect 132647 604864 132648 604865
rect 132648 604863 132649 604864
rect 133082 604852 133093 604863
rect 125106 604818 133093 604852
rect 125767 604806 125768 604807
rect 125010 604206 125068 604806
rect 125768 604805 125769 604806
rect 125780 604350 125814 604818
rect 125826 604806 125827 604807
rect 126525 604806 126526 604807
rect 125825 604805 125826 604806
rect 126526 604805 126527 604806
rect 125734 604216 125854 604350
rect 125734 604202 126450 604216
rect 126526 604206 126527 604207
rect 126525 604205 126526 604206
rect 125780 604194 126450 604202
rect 126538 604194 126572 604818
rect 126584 604806 126585 604807
rect 127283 604806 127284 604807
rect 126583 604805 126584 604806
rect 127284 604805 127285 604806
rect 126583 604206 126584 604207
rect 127284 604206 127285 604207
rect 126584 604205 126585 604206
rect 127283 604205 127284 604206
rect 127296 604194 127330 604818
rect 127342 604806 127343 604807
rect 128041 604806 128042 604807
rect 127341 604805 127342 604806
rect 128042 604805 128043 604806
rect 127341 604206 127342 604207
rect 128042 604206 128043 604207
rect 127342 604205 127343 604206
rect 128041 604205 128042 604206
rect 128054 604194 128088 604818
rect 128100 604806 128101 604807
rect 128099 604805 128100 604806
rect 128538 604598 128572 604818
rect 128712 604812 128714 604818
rect 128686 604806 128712 604812
rect 128714 604806 128740 604812
rect 128799 604806 128800 604807
rect 128712 604800 128714 604806
rect 128800 604805 128801 604806
rect 128812 604800 128846 604818
rect 128908 604814 128940 604818
rect 128908 604812 128956 604814
rect 128858 604806 128859 604807
rect 128900 604806 128911 604811
rect 128857 604805 128858 604806
rect 128900 604800 128912 604806
rect 128708 604794 128916 604800
rect 128602 604756 128674 604794
rect 128708 604784 128984 604794
rect 128724 604766 128911 604784
rect 128712 604760 128772 604762
rect 128640 604722 128674 604756
rect 128712 604732 128772 604734
rect 128812 604712 128846 604766
rect 128912 604762 128984 604784
rect 128896 604760 128984 604762
rect 128912 604756 128984 604760
rect 128896 604732 128940 604734
rect 128900 604712 128911 604723
rect 128950 604722 128984 604756
rect 128724 604678 128911 604712
rect 128812 604598 128846 604678
rect 129052 604598 129086 604818
rect 128538 604564 129086 604598
rect 128812 604408 128846 604564
rect 129136 604506 129774 604818
rect 130315 604806 130316 604807
rect 130316 604805 130317 604806
rect 128794 604402 128908 604408
rect 128099 604206 128100 604207
rect 128800 604206 128801 604207
rect 128100 604205 128101 604206
rect 128799 604205 128800 604206
rect 128812 604194 128846 604402
rect 128857 604206 128858 604207
rect 129558 604206 129559 604207
rect 128858 604205 128859 604206
rect 129557 604205 129558 604206
rect 129570 604194 129604 604506
rect 129615 604206 129616 604207
rect 130316 604206 130317 604207
rect 129616 604205 129617 604206
rect 130315 604205 130316 604206
rect 130328 604194 130362 604818
rect 130374 604806 130375 604807
rect 131073 604806 131074 604807
rect 130373 604805 130374 604806
rect 131074 604805 131075 604806
rect 130373 604206 130374 604207
rect 131074 604206 131075 604207
rect 130374 604205 130375 604206
rect 131073 604205 131074 604206
rect 131086 604194 131120 604818
rect 131132 604806 131133 604807
rect 131831 604806 131832 604807
rect 131131 604805 131132 604806
rect 131832 604805 131833 604806
rect 131131 604206 131132 604207
rect 131832 604206 131833 604207
rect 131132 604205 131133 604206
rect 131831 604205 131832 604206
rect 131844 604194 131878 604818
rect 131890 604806 131891 604807
rect 132589 604806 132590 604807
rect 131889 604805 131890 604806
rect 132590 604805 132591 604806
rect 131889 604206 131890 604207
rect 132590 604206 132591 604207
rect 131890 604205 131891 604206
rect 132589 604205 132590 604206
rect 132602 604194 132636 604818
rect 132648 604806 132649 604807
rect 132647 604805 132648 604806
rect 133094 604790 133166 604828
rect 133132 604222 133166 604790
rect 132647 604206 132648 604207
rect 132648 604205 132649 604206
rect 133082 604194 133093 604205
rect 125106 604160 133093 604194
rect 125767 604148 125768 604149
rect 125010 603901 125068 604148
rect 125768 604147 125769 604148
rect 125780 604142 126450 604160
rect 126525 604148 126526 604149
rect 126526 604147 126527 604148
rect 125682 604118 125730 604132
rect 125780 603901 125814 604142
rect 125854 604118 125926 604132
rect 126430 604118 126532 604132
rect 126538 603901 126572 604160
rect 126584 604148 126585 604149
rect 127283 604148 127284 604149
rect 126583 604147 126584 604148
rect 127284 604147 127285 604148
rect 126578 604118 126694 604132
rect 127296 603901 127330 604160
rect 127342 604148 127343 604149
rect 128041 604148 128042 604149
rect 127341 604147 127342 604148
rect 128042 604147 128043 604148
rect 128054 603901 128088 604160
rect 128100 604148 128101 604149
rect 128799 604148 128800 604149
rect 128099 604147 128100 604148
rect 128800 604147 128801 604148
rect 128812 603966 128846 604160
rect 128858 604148 128859 604149
rect 129557 604148 129558 604149
rect 128857 604147 128858 604148
rect 129558 604147 129559 604148
rect 129038 603966 129170 604084
rect 128790 603901 129238 603966
rect 129570 603901 129604 604160
rect 129616 604148 129617 604149
rect 130315 604148 130316 604149
rect 129615 604147 129616 604148
rect 130316 604147 130317 604148
rect 130328 603901 130362 604160
rect 130374 604148 130375 604149
rect 131073 604148 131074 604149
rect 130373 604147 130374 604148
rect 131074 604147 131075 604148
rect 131086 603901 131120 604160
rect 131132 604148 131133 604149
rect 131831 604148 131832 604149
rect 131131 604147 131132 604148
rect 131832 604147 131833 604148
rect 131844 603901 131878 604160
rect 131890 604148 131891 604149
rect 132589 604148 132590 604149
rect 131889 604147 131890 604148
rect 132590 604147 132591 604148
rect 132602 603901 132636 604160
rect 132648 604148 132649 604149
rect 132647 604147 132648 604148
rect 133094 604132 133166 604170
rect 133132 603901 133166 604132
rect 133234 603901 133268 605214
rect 113180 600449 121387 600505
rect 113087 600421 113121 600425
rect 118808 600394 121387 600449
rect 124861 600394 133299 603901
rect 134876 600616 134910 605164
rect 136334 604568 142254 608788
rect 136334 604548 142294 604568
rect 136294 602464 136295 602465
rect 136293 602463 136294 602464
rect 136334 602424 142254 604548
rect 142256 604129 142257 604548
rect 142294 604129 142314 604548
rect 142256 604128 142314 604129
rect 142542 602476 142606 608840
rect 142723 606227 142757 612591
rect 142887 612545 142954 612558
rect 143402 612545 143479 612558
rect 143545 612545 143612 612558
rect 144060 612545 144137 612558
rect 144203 612545 144274 612558
rect 144722 612545 144795 612558
rect 144861 612545 144944 612558
rect 145392 612545 145453 612558
rect 145519 612545 145596 612558
rect 146044 612545 146111 612558
rect 144153 610033 144187 612492
rect 145469 610033 145503 612492
rect 142825 609999 146173 610033
rect 142837 609965 142871 609999
rect 143495 609978 143529 609999
rect 144153 609978 144187 609999
rect 144811 609978 144845 609999
rect 145469 609978 145503 609999
rect 146127 609978 146161 609999
rect 143467 609965 143529 609978
rect 144125 609965 144187 609978
rect 144783 609965 144845 609978
rect 145441 609965 145503 609978
rect 142837 609863 142877 609965
rect 143467 609937 143535 609965
rect 144125 609937 144193 609965
rect 144783 609937 144851 609965
rect 145441 609937 145509 609965
rect 146099 609937 146161 609978
rect 142887 609931 142905 609937
rect 143461 609931 143535 609937
rect 143545 609931 143563 609937
rect 144119 609931 144193 609937
rect 144203 609931 144221 609937
rect 144777 609931 144851 609937
rect 144861 609931 144879 609937
rect 145435 609931 145509 609937
rect 145519 609931 145537 609937
rect 146093 609931 146161 609937
rect 142883 609897 143535 609931
rect 143541 609897 144193 609931
rect 144199 609897 144851 609931
rect 144857 609897 145509 609931
rect 145515 609897 146161 609931
rect 142887 609891 142905 609897
rect 143461 609891 143479 609897
rect 143489 609863 143535 609897
rect 143545 609891 143563 609897
rect 144119 609891 144137 609897
rect 144147 609863 144193 609897
rect 144203 609891 144221 609897
rect 144777 609891 144795 609897
rect 144805 609863 144851 609897
rect 144861 609891 144879 609897
rect 145435 609891 145453 609897
rect 145463 609863 145509 609897
rect 145519 609891 145537 609897
rect 146093 609891 146111 609897
rect 146121 609863 146161 609897
rect 142837 606323 142871 609863
rect 143396 608792 143402 609316
rect 143495 606323 143529 609863
rect 144153 608978 144187 609863
rect 144811 608978 144845 609863
rect 143816 608686 145298 608978
rect 143732 608238 145298 608686
rect 143816 608044 145298 608238
rect 145469 608044 145503 609863
rect 146084 608792 146100 609260
rect 143816 607672 145870 608044
rect 143816 607402 145298 607672
rect 144153 606323 144187 607402
rect 144811 606323 144845 607402
rect 145469 606323 145503 607672
rect 146127 606323 146161 609863
rect 142787 606289 142791 606323
rect 142825 606289 146173 606323
rect 142837 606268 142871 606289
rect 143495 606268 143529 606289
rect 144153 606268 144187 606289
rect 144811 606268 144845 606289
rect 145469 606268 145503 606289
rect 142691 605386 142757 606227
rect 142825 606221 145726 606268
rect 146067 606221 146114 606268
rect 142837 606187 143482 606221
rect 143495 606187 144140 606221
rect 144153 606187 144798 606221
rect 144811 606187 145456 606221
rect 145469 606187 146114 606221
rect 142837 606140 142883 606187
rect 142912 606181 142922 606187
rect 143402 606181 143447 606187
rect 143495 606181 143580 606187
rect 144060 606181 144105 606187
rect 142793 606128 142811 606140
rect 142837 606128 142882 606140
rect 142894 606138 142912 606181
rect 142922 606138 142940 606181
rect 143495 606140 143541 606181
rect 144112 606153 144133 606187
rect 144153 606140 144199 606187
rect 144220 606181 144242 606187
rect 144722 606181 144763 606187
rect 144811 606181 144912 606187
rect 145392 606181 145421 606187
rect 143452 606128 143483 606139
rect 143495 606128 143540 606140
rect 144110 606128 144141 606139
rect 144153 606128 144198 606140
rect 144214 606138 144220 606181
rect 144242 606138 144248 606181
rect 144811 606140 144857 606181
rect 145432 606153 145449 606187
rect 145469 606140 145515 606187
rect 145540 606181 145564 606187
rect 146044 606181 146079 606187
rect 144768 606128 144799 606139
rect 144811 606128 144856 606140
rect 145426 606128 145457 606139
rect 145469 606128 145514 606140
rect 145536 606138 145540 606181
rect 145564 606138 145568 606181
rect 146084 606128 146115 606139
rect 146127 606128 146161 606289
rect 142793 605386 142882 606128
rect 143463 605386 143540 606128
rect 144121 605386 144198 606128
rect 144779 605386 144856 606128
rect 145437 605386 145514 606128
rect 134180 600532 135136 600566
rect 121215 600391 121249 600394
rect 113049 600357 121287 600391
rect 121215 600202 121249 600357
rect 121215 600116 121304 600202
rect 121215 600042 121249 600116
rect 112949 598970 121364 600042
rect 124897 599714 124931 600394
rect 124984 600347 125604 600394
rect 125654 600347 125688 600394
rect 125788 600384 126442 600394
rect 126186 600347 126220 600384
rect 133127 600377 133161 600381
rect 124961 600313 133195 600347
rect 124984 600304 125604 600313
rect 124961 600218 125604 600304
rect 124984 600034 125604 600218
rect 125654 600086 125688 600313
rect 125694 600312 125836 600313
rect 125849 600312 126118 600313
rect 125709 600266 125790 600312
rect 125849 600294 126036 600312
rect 126037 600266 126118 600312
rect 125756 600228 125790 600266
rect 126084 600228 126118 600266
rect 126025 600200 126036 600211
rect 125849 600166 126036 600200
rect 126186 600086 126220 600313
rect 125654 600052 126220 600086
rect 125392 599880 125494 599896
rect 126032 599880 126438 599882
rect 124961 599771 124988 599828
rect 124999 599809 125026 599866
rect 125420 599852 125494 599868
rect 126032 599852 126410 599854
rect 124961 599742 124988 599757
rect 125092 599747 133068 599781
rect 124897 599684 124993 599714
rect 124999 599704 125026 599719
rect 125039 599684 125390 599714
rect 125420 599704 125694 599714
rect 124897 599668 124931 599684
rect 125039 599668 125220 599684
rect 125420 599668 125620 599704
rect 125836 599668 126410 599714
rect 131428 599698 132780 599714
rect 133229 599668 133263 600394
rect 124861 599006 133263 599668
rect 124842 598970 133263 599006
rect 112949 598936 133263 598970
rect 96481 595155 96515 597713
rect 112949 597667 121364 598936
rect 94816 595121 99255 595155
rect 96481 595041 96515 595121
rect 96583 595075 96617 595121
rect 99221 595063 99255 595121
rect 96536 595041 96617 595048
rect 96676 595041 99255 595063
rect 96447 595029 99255 595041
rect 96447 595017 99060 595029
rect 96447 595007 99071 595017
rect 96481 594383 96515 595007
rect 96536 595001 96664 595007
rect 96567 594995 96664 595001
rect 96583 594433 96617 594995
rect 99072 594979 99153 595026
rect 99119 594417 99153 594979
rect 99072 594405 99169 594417
rect 99221 594405 99255 595029
rect 112980 594971 113014 597667
rect 118920 597352 119326 597667
rect 119570 597352 121364 597667
rect 113055 597341 121364 597352
rect 113066 597329 121364 597341
rect 113055 597318 121364 597329
rect 113082 597272 113116 597318
rect 114096 597272 114554 597292
rect 114096 597260 114594 597272
rect 118920 597260 119326 597318
rect 119570 597260 121364 597318
rect 113166 597204 121364 597260
rect 114096 597200 114594 597204
rect 113082 596608 113116 597198
rect 114136 597180 114594 597200
rect 113746 597156 114850 597176
rect 113718 597128 114878 597148
rect 118762 597142 118818 597148
rect 119446 597142 119502 597148
rect 117006 596996 117454 597024
rect 117006 596812 117472 596996
rect 117024 596784 117472 596812
rect 119456 596616 119502 596640
rect 119570 596613 121364 597204
rect 116120 596602 121364 596613
rect 113166 596546 121364 596602
rect 113082 596518 113116 596522
rect 119570 596488 121364 596546
rect 113035 596454 121364 596488
rect 117012 596140 117460 596352
rect 116474 595576 117112 596038
rect 117162 595950 117710 595984
rect 117162 595922 117196 595950
rect 117676 595922 117710 595950
rect 117162 595888 117230 595922
rect 117310 595904 117562 595908
rect 117308 595888 117564 595904
rect 117162 595884 117196 595888
rect 117308 595884 117340 595888
rect 117162 595882 117340 595884
rect 117534 595882 117564 595888
rect 117676 595888 117744 595922
rect 117162 595668 117196 595882
rect 117336 595870 117536 595876
rect 117336 595864 117340 595870
rect 117226 595856 117340 595864
rect 117212 595854 117340 595856
rect 117348 595864 117536 595870
rect 117348 595854 117646 595864
rect 117226 595832 117336 595854
rect 117348 595836 117535 595854
rect 117536 595832 117646 595854
rect 117226 595830 117646 595832
rect 117226 595826 117336 595830
rect 117536 595826 117646 595830
rect 117264 595804 117336 595826
rect 117264 595802 117564 595804
rect 117264 595792 117336 595802
rect 117337 595782 117535 595793
rect 117574 595792 117646 595826
rect 117348 595748 117535 595782
rect 117676 595668 117710 595888
rect 117162 595634 117710 595668
rect 119570 595202 121364 596454
rect 119450 595188 121364 595202
rect 117078 595036 117210 595154
rect 117010 594971 117458 595036
rect 119570 594971 121364 595188
rect 96676 594383 99255 594405
rect 96481 594371 99255 594383
rect 96481 594349 99060 594371
rect 99072 594359 99200 594368
rect 96481 594291 96515 594349
rect 99119 594321 99153 594325
rect 99221 594291 99255 594371
rect 96481 594257 104751 594291
rect 99221 593342 99255 594257
rect 112949 593764 121364 594971
rect 124842 597693 133263 598936
rect 136302 600214 142254 602424
rect 124842 597623 133262 597693
rect 124842 597316 129078 597623
rect 124842 597104 129196 597316
rect 124842 596978 129078 597104
rect 124842 596967 133151 596978
rect 124842 596955 133140 596967
rect 124842 596944 133151 596955
rect 124842 596886 129078 596944
rect 131652 596898 132110 596918
rect 133090 596898 133124 596944
rect 131612 596886 132110 596898
rect 124842 596840 133040 596886
rect 124842 596830 133051 596840
rect 124842 596650 129078 596830
rect 131612 596826 132110 596830
rect 131612 596806 132070 596826
rect 131356 596782 132460 596802
rect 131328 596754 132488 596774
rect 124842 596438 129200 596650
rect 124842 596410 129182 596438
rect 124842 596228 129078 596410
rect 133040 596228 133051 596239
rect 133090 596234 133124 596824
rect 124842 596218 133051 596228
rect 124842 596172 133040 596218
rect 124842 596114 129078 596172
rect 133090 596144 133124 596148
rect 124842 596080 133158 596114
rect 124842 595978 129078 596080
rect 124842 595766 129194 595978
rect 124842 594780 129078 595766
rect 129094 595202 129732 595664
rect 133090 594918 133124 595486
rect 132448 594856 133148 594890
rect 124842 594662 129128 594780
rect 133090 594692 133124 594828
rect 133192 594692 133226 597623
rect 136262 595792 136263 595793
rect 136261 595791 136262 595792
rect 136302 595752 142222 600214
rect 142262 600174 142263 600175
rect 142261 600173 142262 600174
rect 142510 600162 142606 602476
rect 142655 605212 145672 605386
rect 142655 605018 145870 605212
rect 142655 604504 145672 605018
rect 146095 604950 146161 606128
rect 146209 606227 146227 606289
rect 146241 606227 146275 612591
rect 147106 608832 147142 608848
rect 147794 606232 147828 612596
rect 147958 612550 148040 612558
rect 148488 612550 148550 612558
rect 148616 612550 148692 612558
rect 149140 612550 149208 612558
rect 149274 612550 149350 612558
rect 149798 612550 149866 612558
rect 149932 612550 150014 612558
rect 150462 612550 150524 612558
rect 150590 612550 150666 612558
rect 151114 612550 151182 612558
rect 147896 610004 151244 610038
rect 147908 609970 147942 610004
rect 148566 609974 148600 610004
rect 149224 609974 149258 610004
rect 149882 609974 149916 610004
rect 150540 609974 150574 610004
rect 151198 609974 151232 610004
rect 148538 609970 148600 609974
rect 147908 609868 147948 609970
rect 148538 609942 148606 609970
rect 149196 609942 150204 609974
rect 150512 609970 150574 609974
rect 150512 609942 150580 609970
rect 151170 609942 151232 609974
rect 147958 609936 147976 609942
rect 148532 609936 148606 609942
rect 148616 609936 148634 609942
rect 149190 609936 150204 609942
rect 150506 609936 150580 609942
rect 150590 609936 150608 609942
rect 151164 609936 151232 609942
rect 147954 609902 148606 609936
rect 148612 609902 149264 609936
rect 147958 609896 147976 609902
rect 148532 609896 148550 609902
rect 148560 609868 148606 609902
rect 148616 609896 148634 609902
rect 149190 609896 149208 609902
rect 149218 609868 149264 609902
rect 149274 609902 149922 609936
rect 149274 609896 149292 609902
rect 149848 609896 149866 609902
rect 149876 609868 149922 609902
rect 149932 609902 150580 609936
rect 150586 609902 151232 609936
rect 149932 609896 149950 609902
rect 150506 609896 150524 609902
rect 150534 609868 150580 609902
rect 150590 609896 150608 609902
rect 151164 609896 151182 609902
rect 151192 609868 151232 609902
rect 147908 606328 147942 609868
rect 148566 606328 148600 609868
rect 149224 606328 149258 609868
rect 149882 606328 149916 609868
rect 150540 606328 150574 609868
rect 151198 606328 151232 609868
rect 147858 606294 147862 606328
rect 147896 606294 151244 606328
rect 147908 606264 147942 606294
rect 148566 606264 148600 606294
rect 149224 606264 149258 606294
rect 149882 606264 149916 606294
rect 150540 606264 150574 606294
rect 146209 605386 146275 606227
rect 146024 604504 146044 604950
rect 146052 604504 146161 604950
rect 142655 604423 146161 604504
rect 142655 604355 145672 604423
rect 146083 604407 146161 604423
rect 146089 604355 146161 604407
rect 142655 604321 146195 604355
rect 142655 603669 145672 604321
rect 146089 603976 146161 604321
rect 146095 603703 146161 603976
rect 146095 603669 146181 603703
rect 142655 603635 146181 603669
rect 142655 603567 145672 603635
rect 146095 603614 146161 603635
rect 146067 603567 146161 603614
rect 142655 603533 146161 603567
rect 142655 601803 145672 603533
rect 146024 602120 146044 602788
rect 146052 602120 146072 602788
rect 146095 601862 146161 603533
rect 146095 601850 146129 601862
rect 146083 601803 146141 601850
rect 142655 601769 146141 601803
rect 142655 601701 145672 601769
rect 146083 601753 146129 601769
rect 142655 601667 146141 601701
rect 142655 600394 145672 601667
rect 142510 595804 142574 600162
rect 142691 599555 142725 600394
rect 142805 599651 142839 600394
rect 143463 599651 143497 600394
rect 144121 599651 144155 600394
rect 144779 599651 144813 600394
rect 145042 599651 145254 599668
rect 145437 599651 145471 600394
rect 146095 599651 146129 601667
rect 146208 601631 146311 605386
rect 147762 605350 147828 606232
rect 147904 606226 148544 606264
rect 148562 606226 149202 606264
rect 149220 606226 149860 606264
rect 149878 606226 150518 606264
rect 150536 606226 151176 606264
rect 147908 606192 148544 606226
rect 148566 606222 149202 606226
rect 148566 606192 149204 606222
rect 147908 606154 147954 606192
rect 147980 606186 148008 606192
rect 148488 606186 148518 606192
rect 148566 606186 148660 606192
rect 149140 606186 149176 606192
rect 148566 606154 148612 606186
rect 149182 606158 149204 606192
rect 149224 606192 149860 606226
rect 149882 606192 150518 606226
rect 150540 606192 151176 606226
rect 149224 606154 149270 606192
rect 149290 606186 149318 606192
rect 149798 606186 149834 606192
rect 149882 606186 149982 606192
rect 150462 606186 150492 606192
rect 149882 606154 149928 606186
rect 150504 606158 150520 606186
rect 150540 606154 150586 606192
rect 150612 606186 150634 606192
rect 151114 606186 151150 606192
rect 147864 606142 147882 606154
rect 147908 606142 147953 606154
rect 148523 606142 148554 606153
rect 148566 606142 148611 606154
rect 149181 606142 149212 606153
rect 149224 606142 149269 606154
rect 149839 606142 149870 606153
rect 149882 606142 149927 606154
rect 150497 606142 150528 606153
rect 150540 606142 150585 606154
rect 147864 605350 147953 606142
rect 148534 605350 148611 606142
rect 149192 605350 149269 606142
rect 149850 605350 149927 606142
rect 150508 605350 150585 606142
rect 150606 606138 150612 606186
rect 150634 606138 150640 606186
rect 151155 606142 151186 606153
rect 151198 606142 151232 606294
rect 151166 605350 151232 606142
rect 151280 606232 151298 606294
rect 151312 606232 151346 612596
rect 189293 611385 189359 613195
rect 189435 613205 189439 613223
rect 189435 613189 189485 613205
rect 189496 613195 189514 613210
rect 189524 613195 189542 613208
rect 190037 613189 190084 613236
rect 190093 613205 190097 613223
rect 190093 613189 190143 613205
rect 190695 613195 190742 613236
rect 190686 613189 190742 613195
rect 190751 613205 190755 613223
rect 190751 613189 190801 613205
rect 190816 613195 190822 613198
rect 190844 613195 190850 613208
rect 191353 613189 191400 613236
rect 191409 613205 191413 613223
rect 191409 613189 191459 613205
rect 192011 613195 192058 613236
rect 192006 613189 192058 613195
rect 192067 613205 192071 613223
rect 192067 613189 192117 613205
rect 192669 613189 192716 613236
rect 189439 613155 190084 613189
rect 190097 613155 190742 613189
rect 190755 613155 191400 613189
rect 191413 613155 192058 613189
rect 192071 613155 192716 613189
rect 189439 613108 189485 613155
rect 189395 613096 189413 613108
rect 189439 613096 189473 613108
rect 189395 611484 189473 613096
rect 189496 611808 189514 613149
rect 189524 611780 189542 613149
rect 190097 613108 190143 613155
rect 190686 613149 190707 613155
rect 190714 613121 190735 613155
rect 190755 613108 190801 613155
rect 190054 613096 190085 613107
rect 190097 613096 190131 613108
rect 190712 613096 190743 613107
rect 190755 613096 190789 613108
rect 189293 609576 189327 611385
rect 189395 611323 189441 611484
rect 189994 611431 190004 612830
rect 190022 611459 190032 612802
rect 190065 611484 190131 613096
rect 190723 611484 190789 613096
rect 190816 611796 190822 613149
rect 190844 611768 190850 613149
rect 191413 613108 191459 613155
rect 192006 613149 192023 613155
rect 192034 613121 192051 613155
rect 192071 613108 192117 613155
rect 191370 613096 191401 613107
rect 191413 613096 191447 613108
rect 192028 613096 192059 613107
rect 192071 613096 192105 613108
rect 190065 611472 190099 611484
rect 190723 611472 190757 611484
rect 190053 611459 190112 611472
rect 190022 611450 190112 611459
rect 190119 611450 190150 611459
rect 190053 611431 190112 611450
rect 189994 611425 190112 611431
rect 189501 611391 190112 611425
rect 190147 611425 190178 611431
rect 190711 611425 190770 611472
rect 191304 611431 191324 612836
rect 191332 611459 191352 612808
rect 191381 611484 191447 613096
rect 192039 611484 192105 613096
rect 192138 611774 192142 613149
rect 192166 611746 192170 613149
rect 192686 613096 192717 613107
rect 192729 613096 192763 613257
rect 191381 611472 191415 611484
rect 192039 611472 192073 611484
rect 191369 611459 191428 611472
rect 191332 611456 191428 611459
rect 191435 611456 191460 611459
rect 191369 611431 191428 611456
rect 191304 611428 191428 611431
rect 191463 611428 191488 611431
rect 191369 611425 191428 611428
rect 192027 611425 192086 611472
rect 192626 611431 192646 612806
rect 192654 611431 192674 612778
rect 192697 611484 192763 613096
rect 192811 613195 192829 613257
rect 192843 613195 192877 613502
rect 194396 613200 194430 613502
rect 194510 613296 194544 613330
rect 195168 613296 195202 613330
rect 195826 613296 195860 613330
rect 196484 613296 196518 613330
rect 197142 613296 197176 613330
rect 197800 613296 197854 613330
rect 194460 613262 194464 613296
rect 194476 613262 197854 613296
rect 192697 611472 192731 611484
rect 192685 611425 192743 611472
rect 190147 611422 190770 611425
rect 190159 611391 190770 611422
rect 190817 611391 191428 611425
rect 191475 611391 192086 611425
rect 192133 611391 192743 611425
rect 190053 611375 190099 611391
rect 190711 611375 190757 611391
rect 191369 611375 191415 611391
rect 192027 611375 192073 611391
rect 192685 611375 192731 611391
rect 192811 611385 192877 613195
rect 194364 611408 194430 613200
rect 194506 613210 194510 613228
rect 194506 613194 194556 613210
rect 195108 613194 195146 613232
rect 195164 613210 195168 613228
rect 195164 613194 195214 613210
rect 195766 613200 195804 613232
rect 195756 613194 195804 613200
rect 195822 613210 195826 613228
rect 195822 613194 195872 613210
rect 196424 613194 196462 613232
rect 196480 613210 196484 613228
rect 196480 613194 196530 613210
rect 197082 613194 197120 613232
rect 197138 613210 197142 613228
rect 197138 613194 197188 613210
rect 197740 613194 197778 613232
rect 194510 613160 195146 613194
rect 195168 613190 195804 613194
rect 195168 613160 195806 613190
rect 194510 613122 194556 613160
rect 195168 613122 195214 613160
rect 195756 613154 195778 613160
rect 195784 613126 195806 613160
rect 195826 613160 196462 613194
rect 196484 613160 197120 613194
rect 197142 613160 197778 613194
rect 195826 613122 195872 613160
rect 196484 613122 196530 613160
rect 197078 613154 197094 613160
rect 197106 613126 197122 613154
rect 197142 613122 197188 613160
rect 194466 613110 194484 613122
rect 194510 613110 194544 613122
rect 195125 613110 195156 613121
rect 195168 613110 195202 613122
rect 195783 613110 195814 613121
rect 195826 613110 195860 613122
rect 196441 613110 196472 613121
rect 196484 613110 196518 613122
rect 197099 613110 197130 613121
rect 197142 613110 197176 613122
rect 194466 611498 194544 613110
rect 192039 611323 192073 611375
rect 189395 611289 192743 611323
rect 192039 609576 192073 611289
rect 192811 609576 192845 611385
rect 189293 609538 192845 609576
rect 167126 608678 167132 608690
rect 167318 608678 167326 608690
rect 167098 608650 167132 608662
rect 167318 608650 167354 608662
rect 166588 608226 167154 608260
rect 166588 608131 166622 608226
rect 166959 608146 166970 608157
rect 166783 608143 166970 608146
rect 166783 608131 166959 608143
rect 167120 608131 167154 608226
rect 166554 608097 167154 608131
rect 166588 607904 166622 608097
rect 166643 608085 166771 608097
rect 166971 608085 167068 608097
rect 166643 608084 166724 608085
rect 166971 608084 167052 608085
rect 166690 608046 166724 608084
rect 167018 608046 167052 608084
rect 166680 608020 166732 608032
rect 166959 608018 166970 608029
rect 166652 607992 166760 608004
rect 166783 607984 166970 608018
rect 167104 608004 167106 608091
rect 167120 607904 167154 608097
rect 166588 607870 167154 607904
rect 167204 608069 167824 608274
rect 171962 608072 172092 608093
rect 167204 607852 167851 608069
rect 171776 608047 172092 608072
rect 172278 608047 172684 608093
rect 171804 608019 172092 608044
rect 172278 608019 172628 608044
rect 167817 607798 167851 607852
rect 166588 607750 167154 607784
rect 166588 607462 166622 607750
rect 166959 607670 166970 607681
rect 166643 607608 166724 607655
rect 166783 607636 166970 607670
rect 166971 607608 167052 607655
rect 166690 607570 166724 607608
rect 167018 607570 167052 607608
rect 167120 607556 167154 607750
rect 166959 607542 166970 607553
rect 167086 607542 167106 607556
rect 166783 607508 166970 607542
rect 167010 607528 167106 607542
rect 167114 607542 167154 607556
rect 167204 607646 167851 607798
rect 167204 607560 167906 607646
rect 167204 607542 167851 607560
rect 167114 607522 167851 607542
rect 167120 607514 167154 607522
rect 167204 607514 167851 607522
rect 166982 607501 167851 607514
rect 166982 607500 167824 607501
rect 167086 607494 167824 607500
rect 166745 607470 166997 607473
rect 167120 607462 167154 607494
rect 166588 607439 167154 607462
rect 166588 607428 166622 607439
rect 167120 607428 167154 607439
rect 166588 607427 167154 607428
rect 166622 607413 167120 607427
rect 166588 607394 167154 607413
rect 167204 607376 167824 607494
rect 171586 607478 172206 607900
rect 172256 607852 172822 607886
rect 172256 607530 172290 607852
rect 172627 607772 172638 607783
rect 172311 607710 172392 607757
rect 172451 607738 172638 607772
rect 172639 607710 172720 607757
rect 172358 607672 172392 607710
rect 172686 607672 172720 607710
rect 172627 607644 172638 607655
rect 172451 607610 172638 607644
rect 172788 607530 172822 607852
rect 172256 607496 172822 607530
rect 171644 607424 171662 607463
rect 171962 607435 171992 607470
rect 172018 607435 172020 607470
rect 171678 607424 171696 607429
rect 171586 607378 172206 607424
rect 172318 607410 172760 607444
rect 172256 607383 172822 607410
rect 171586 607376 172266 607378
rect 171586 607362 172324 607376
rect 171586 607350 172206 607362
rect 171586 607348 172238 607350
rect 171586 607315 172296 607348
rect 171586 607281 175456 607315
rect 171586 607245 172206 607281
rect 172256 607148 172296 607281
rect 172304 607154 172324 607274
rect 172358 607247 172392 607250
rect 172686 607247 172720 607250
rect 172256 607116 172290 607148
rect 172788 607116 172822 607281
rect 151280 605350 151346 606232
rect 152206 605386 152446 605722
rect 151730 605350 152192 605386
rect 146340 605316 152192 605350
rect 147070 605308 147228 605316
rect 146370 605180 146388 605282
rect 147762 605248 147828 605316
rect 147864 605312 147953 605316
rect 148534 605312 148611 605316
rect 147864 605248 147942 605312
rect 148534 605264 148600 605312
rect 149192 605286 149269 605316
rect 149850 605286 149927 605316
rect 150508 605312 150585 605316
rect 148522 605248 148600 605264
rect 148604 605248 148642 605286
rect 149192 605264 149400 605286
rect 149180 605248 149400 605264
rect 149414 605248 150158 605286
rect 150508 605264 150574 605312
rect 150496 605248 150574 605264
rect 150878 605248 150916 605286
rect 151166 605279 151232 605316
rect 151166 605264 151244 605279
rect 151154 605248 151244 605264
rect 146404 605214 146422 605248
rect 147178 605214 147862 605248
rect 147864 605214 148642 605248
rect 148694 605214 149400 605248
rect 149452 605214 150158 605248
rect 150210 605214 150916 605248
rect 150968 605214 151244 605248
rect 147024 604386 147142 604488
rect 147024 604366 147190 604386
rect 147070 604238 147190 604366
rect 147762 604378 147828 605214
rect 147864 605176 147942 605214
rect 148522 605176 148600 605214
rect 147876 605164 147942 605176
rect 147874 604542 147942 605164
rect 147952 604814 147980 604950
rect 147874 604384 147948 604542
rect 147958 604480 147976 604486
rect 148534 604480 148600 605176
rect 148632 605175 148634 605180
rect 149180 605176 149269 605214
rect 149838 605176 149927 605214
rect 150496 605176 150574 605214
rect 151154 605176 151244 605214
rect 148621 605164 148666 605175
rect 148632 604518 148666 605164
rect 149192 604950 149269 605176
rect 149379 605164 149435 605175
rect 149192 604518 149298 604950
rect 149318 604518 149354 604950
rect 149390 604518 149435 605164
rect 149850 604518 149927 605176
rect 150137 605164 150193 605175
rect 150148 604518 150193 605164
rect 148632 604480 148670 604518
rect 149192 604480 150204 604518
rect 150508 604480 150574 605176
rect 150895 605164 150940 605175
rect 150906 604518 150940 605164
rect 150906 604480 150944 604518
rect 151166 604480 151232 605176
rect 147954 604446 148600 604480
rect 148612 604446 149269 604480
rect 149286 604446 149927 604480
rect 149944 604446 150574 604480
rect 150586 604446 151232 604480
rect 147958 604440 147976 604446
rect 147874 604382 147942 604384
rect 148534 604382 148600 604446
rect 148632 604382 148666 604446
rect 149192 604440 149269 604446
rect 147874 604378 147953 604382
rect 148534 604378 148611 604382
rect 148632 604378 148677 604382
rect 149192 604378 149298 604440
rect 149318 604378 149354 604440
rect 149390 604378 149435 604446
rect 149850 604378 149927 604446
rect 150148 604378 150193 604446
rect 150508 604382 150574 604446
rect 150906 604382 150940 604446
rect 151166 604382 151232 604446
rect 150508 604378 150585 604382
rect 150906 604378 150951 604382
rect 151166 604378 151243 604382
rect 151280 604378 151346 605316
rect 151382 605302 151612 605310
rect 151556 605208 151612 605216
rect 151730 605084 152192 605316
rect 152206 605084 152668 605386
rect 159582 605350 159616 606878
rect 167896 605350 167930 606878
rect 189293 606523 189327 609538
rect 192039 609520 192073 609538
rect 189362 609482 192780 609520
rect 189407 606619 189441 606653
rect 190065 606619 190099 606653
rect 190723 606619 190757 606653
rect 191381 606619 191415 606653
rect 192039 606619 192073 609482
rect 192697 606619 192731 606653
rect 189375 606585 192765 606619
rect 171480 605350 171514 606504
rect 155296 605316 173036 605350
rect 159582 605248 159616 605316
rect 159684 605248 159718 605316
rect 159974 605248 160012 605286
rect 160732 605248 160770 605286
rect 161490 605248 161528 605286
rect 162248 605248 162286 605286
rect 163006 605248 163044 605286
rect 163764 605248 163802 605286
rect 164522 605248 164560 605286
rect 165280 605248 165318 605286
rect 166038 605248 166076 605286
rect 166796 605248 166834 605286
rect 167554 605248 167592 605286
rect 167794 605248 167828 605316
rect 167896 605248 167930 605316
rect 159582 605214 160012 605248
rect 160064 605214 160770 605248
rect 160822 605214 161528 605248
rect 161580 605214 162286 605248
rect 162338 605214 163044 605248
rect 163096 605214 163802 605248
rect 163854 605214 164560 605248
rect 164612 605214 165318 605248
rect 165370 605214 166076 605248
rect 166128 605214 166834 605248
rect 166886 605214 167592 605248
rect 167644 605214 167930 605248
rect 170572 605214 170602 605248
rect 151784 605000 152134 605034
rect 151594 604960 151618 604986
rect 151622 604932 151646 604958
rect 151556 604886 151582 604912
rect 147762 604344 151346 604378
rect 147762 603674 147828 604344
rect 147874 603674 147953 604344
rect 148534 603674 148611 604344
rect 148632 603674 148677 604344
rect 149192 603976 149298 604344
rect 149318 603976 149354 604344
rect 149192 603674 149269 603976
rect 149390 603674 149435 604344
rect 149850 603674 149927 604344
rect 150148 603674 150193 604344
rect 150508 603674 150585 604344
rect 150906 603674 150951 604344
rect 151166 603708 151243 604344
rect 151166 603674 151252 603708
rect 151280 603674 151346 604344
rect 151594 604308 151606 604662
rect 151622 604308 151634 604662
rect 151784 604520 151818 605000
rect 151976 604932 152014 604970
rect 151942 604898 152014 604932
rect 151887 604848 151932 604859
rect 151975 604848 152020 604859
rect 151898 604672 151932 604848
rect 151986 604672 152020 604848
rect 151976 604622 152014 604660
rect 151942 604588 152014 604622
rect 152100 604520 152134 605000
rect 151784 604486 152134 604520
rect 152260 605000 152610 605034
rect 152260 604520 152294 605000
rect 152422 604966 152460 604970
rect 152422 604948 152486 604966
rect 152410 604898 152486 604948
rect 152410 604882 152468 604898
rect 152388 604860 152408 604864
rect 152388 604859 152414 604860
rect 152363 604848 152414 604859
rect 152374 604672 152414 604848
rect 152388 604660 152414 604672
rect 152416 604660 152456 604882
rect 152462 604859 152490 604864
rect 152462 604672 152496 604859
rect 152388 604656 152408 604660
rect 152416 604656 152460 604660
rect 152462 604656 152490 604672
rect 152416 604638 152486 604656
rect 152410 604588 152486 604638
rect 152410 604572 152468 604588
rect 152576 604520 152610 605000
rect 152260 604486 152610 604520
rect 151622 604252 151662 604308
rect 147762 603640 151346 603674
rect 146476 602254 146502 602260
rect 146504 602254 146530 602288
rect 146884 602196 147346 602834
rect 146942 602112 147292 602146
rect 146942 601632 146976 602112
rect 147062 602078 147154 602082
rect 147062 602044 147168 602078
rect 147100 602010 147168 602044
rect 147104 601972 147150 602010
rect 147045 601960 147101 601971
rect 147056 601784 147101 601960
rect 147116 601960 147150 601972
rect 147162 601960 147189 601971
rect 147116 601784 147189 601960
rect 147116 601772 147150 601784
rect 147062 601768 147154 601772
rect 147062 601734 147168 601768
rect 147100 601700 147168 601734
rect 147104 601684 147150 601700
rect 147258 601632 147292 602112
rect 146208 601606 146279 601631
rect 146942 601606 147292 601632
rect 147762 601724 147828 603640
rect 147874 603610 147953 603640
rect 148534 603610 148611 603640
rect 148632 603610 148677 603640
rect 149192 603610 149269 603640
rect 149390 603610 149435 603640
rect 149850 603610 149927 603640
rect 150148 603610 150193 603640
rect 150508 603610 150585 603640
rect 150906 603610 150951 603640
rect 151166 603610 151243 603640
rect 147874 603538 151243 603610
rect 147874 603282 147953 603538
rect 148534 603282 148611 603538
rect 148632 603282 148677 603538
rect 147874 603144 147942 603282
rect 148534 603144 148600 603282
rect 148632 603144 148666 603282
rect 149192 603220 149269 603538
rect 147874 602788 147953 603144
rect 147874 602198 147980 602788
rect 147874 602128 147953 602198
rect 147954 602160 147970 602176
rect 147970 602156 147976 602160
rect 147874 602120 147954 602128
rect 147970 602120 147982 602156
rect 147874 602104 147970 602120
rect 147874 601876 147953 602104
rect 148534 601876 148611 603144
rect 147874 601724 147910 601876
rect 147920 601724 147921 601876
rect 148534 601864 148579 601876
rect 148632 601864 148677 603144
rect 149192 603112 149280 603220
rect 148888 602788 149280 603112
rect 148888 602604 149298 602788
rect 149192 602120 149298 602604
rect 149318 602120 149354 602788
rect 149192 601876 149269 602120
rect 149192 601864 149237 601876
rect 149390 601864 149435 603538
rect 149850 601876 149927 603538
rect 149850 601864 149895 601876
rect 150148 601864 150193 603538
rect 150508 603470 150585 603538
rect 150906 603470 150951 603538
rect 150508 603212 150574 603470
rect 150508 603146 150596 603212
rect 150360 602638 150682 603146
rect 150906 603144 150940 603470
rect 150966 603454 150974 603470
rect 151166 603444 151243 603538
rect 151166 603144 151232 603444
rect 150508 602558 150596 602638
rect 150508 601876 150585 602558
rect 150508 601864 150553 601876
rect 150906 601864 150951 603144
rect 151166 601876 151243 603144
rect 151166 601864 151211 601876
rect 147932 601826 148579 601864
rect 148590 601826 149237 601864
rect 149248 601826 149895 601864
rect 149906 601826 150553 601864
rect 150564 601826 151211 601864
rect 147970 601792 148579 601826
rect 148628 601803 149237 601826
rect 148621 601792 149237 601803
rect 149286 601792 149895 601826
rect 149944 601792 150553 601826
rect 150602 601792 151211 601826
rect 148534 601724 148579 601792
rect 148632 601724 148677 601792
rect 149192 601724 149237 601792
rect 149390 601724 149435 601792
rect 149850 601724 149895 601792
rect 150148 601724 150193 601792
rect 150508 601724 150553 601792
rect 150906 601724 150951 601792
rect 151166 601724 151211 601792
rect 151280 601724 151346 603640
rect 151730 602430 152192 603068
rect 152206 602430 152668 603068
rect 151784 602346 152134 602380
rect 151556 602232 151582 602258
rect 151556 602176 151638 602202
rect 151784 601866 151818 602346
rect 151924 602318 151930 602320
rect 151994 602318 152004 602320
rect 151904 602278 152014 602316
rect 151942 602248 152014 602278
rect 151924 602246 152014 602248
rect 151942 602244 152014 602246
rect 151887 602194 151943 602205
rect 151975 602194 152031 602205
rect 151898 602018 151943 602194
rect 151986 602018 152031 602194
rect 151904 601968 152014 602006
rect 151942 601934 152014 601968
rect 152100 601866 152134 602346
rect 151784 601832 152134 601866
rect 152260 602346 152610 602380
rect 152260 601866 152294 602346
rect 152400 602318 152406 602320
rect 152380 602312 152460 602316
rect 152380 602278 152486 602312
rect 152410 602248 152486 602278
rect 152400 602246 152486 602248
rect 152410 602244 152486 602246
rect 152410 602228 152468 602244
rect 152368 602205 152414 602206
rect 152363 602202 152414 602205
rect 152360 602144 152414 602202
rect 152416 602202 152456 602228
rect 152468 602202 152507 602205
rect 152416 602144 152507 602202
rect 152374 602018 152410 602144
rect 152420 602006 152456 602144
rect 152462 602018 152507 602144
rect 152380 602002 152460 602006
rect 152380 601968 152486 602002
rect 152410 601934 152486 601968
rect 152410 601918 152468 601934
rect 152576 601866 152610 602346
rect 152260 601832 152610 601866
rect 147762 601690 151346 601724
rect 147762 601606 147796 601690
rect 147874 601606 147910 601690
rect 147920 601606 147921 601690
rect 148534 601606 148579 601690
rect 148632 601606 148677 601690
rect 149192 601606 149237 601690
rect 149390 601606 149435 601690
rect 149850 601606 149895 601690
rect 150148 601606 150193 601690
rect 150508 601606 150553 601690
rect 150906 601606 150951 601690
rect 151166 601606 151211 601690
rect 151280 601606 151314 601690
rect 158486 601606 158520 605164
rect 159582 603456 159616 605214
rect 159684 604914 159718 605214
rect 159756 605176 159757 605177
rect 167755 605176 167756 605177
rect 159755 605175 159756 605176
rect 167756 605175 167757 605176
rect 159991 605164 160036 605175
rect 160749 605164 160794 605175
rect 161507 605164 161552 605175
rect 162265 605164 162310 605175
rect 163023 605164 163068 605175
rect 163781 605164 163826 605175
rect 164539 605164 164584 605175
rect 165297 605164 165342 605175
rect 166055 605164 166100 605175
rect 166813 605164 166858 605175
rect 167571 605164 167616 605175
rect 159990 604898 159991 604899
rect 159989 604897 159990 604898
rect 160002 604886 160036 605164
rect 160047 604898 160048 604899
rect 160748 604898 160749 604899
rect 160048 604897 160049 604898
rect 160747 604897 160748 604898
rect 160760 604886 160794 605164
rect 160805 604898 160806 604899
rect 161506 604898 161507 604899
rect 160806 604897 160807 604898
rect 161505 604897 161506 604898
rect 161518 604886 161552 605164
rect 161563 604898 161564 604899
rect 162264 604898 162265 604899
rect 161564 604897 161565 604898
rect 162263 604897 162264 604898
rect 162276 604886 162310 605164
rect 162321 604898 162322 604899
rect 163022 604898 163023 604899
rect 162322 604897 162323 604898
rect 163021 604897 163022 604898
rect 163034 604886 163068 605164
rect 163718 604978 163786 604986
rect 163746 604950 163786 604958
rect 163079 604898 163080 604899
rect 163780 604898 163781 604899
rect 163080 604897 163081 604898
rect 163779 604897 163780 604898
rect 163792 604886 163826 605164
rect 163832 604978 163898 604986
rect 163832 604950 163870 604958
rect 163837 604898 163838 604899
rect 164538 604898 164539 604899
rect 163838 604897 163839 604898
rect 164537 604897 164538 604898
rect 164550 604886 164584 605164
rect 165232 604978 165302 604998
rect 165260 604950 165302 604970
rect 164595 604898 164596 604899
rect 165296 604898 165297 604899
rect 164596 604897 164597 604898
rect 165295 604897 165296 604898
rect 165308 604886 165342 605164
rect 165348 604978 165412 604998
rect 165348 604950 165384 604970
rect 165353 604898 165354 604899
rect 166054 604898 166055 604899
rect 165354 604897 165355 604898
rect 166053 604897 166054 604898
rect 166066 604886 166100 605164
rect 166111 604898 166112 604899
rect 166812 604898 166813 604899
rect 166112 604897 166113 604898
rect 166811 604897 166812 604898
rect 166824 604886 166858 605164
rect 166869 604898 166870 604899
rect 167570 604898 167571 604899
rect 166870 604897 166871 604898
rect 167569 604897 167570 604898
rect 167582 604886 167616 605164
rect 167794 604914 167828 605214
rect 167627 604898 167628 604899
rect 167628 604897 167629 604898
rect 167744 604886 167755 604897
rect 159646 604824 159718 604862
rect 159768 604852 167755 604886
rect 159989 604840 159990 604841
rect 159990 604839 159991 604840
rect 159684 604256 159718 604824
rect 159990 604240 159991 604241
rect 159989 604239 159990 604240
rect 160002 604228 160036 604852
rect 160048 604840 160049 604841
rect 160747 604840 160748 604841
rect 160047 604839 160048 604840
rect 160748 604839 160749 604840
rect 160760 604272 160794 604852
rect 160806 604840 160807 604841
rect 161505 604840 161506 604841
rect 160805 604839 160806 604840
rect 161506 604839 161507 604840
rect 160716 604266 160836 604272
rect 160047 604240 160048 604241
rect 160748 604240 160749 604241
rect 160048 604239 160049 604240
rect 160747 604239 160748 604240
rect 160760 604228 160794 604266
rect 160805 604240 160806 604241
rect 161506 604240 161507 604241
rect 160806 604239 160807 604240
rect 161505 604239 161506 604240
rect 161518 604228 161552 604852
rect 161564 604840 161565 604841
rect 162263 604840 162264 604841
rect 161563 604839 161564 604840
rect 162264 604839 162265 604840
rect 161563 604240 161564 604241
rect 162264 604240 162265 604241
rect 161564 604239 161565 604240
rect 162263 604239 162264 604240
rect 162276 604228 162310 604852
rect 162322 604840 162323 604841
rect 163021 604840 163022 604841
rect 162321 604839 162322 604840
rect 163022 604839 163023 604840
rect 162321 604240 162322 604241
rect 163022 604240 163023 604241
rect 162322 604239 162323 604240
rect 163021 604239 163022 604240
rect 163034 604228 163068 604852
rect 163080 604840 163081 604841
rect 163779 604840 163780 604841
rect 163079 604839 163080 604840
rect 163780 604839 163781 604840
rect 163079 604240 163080 604241
rect 163780 604240 163781 604241
rect 163080 604239 163081 604240
rect 163779 604239 163780 604240
rect 163792 604228 163826 604852
rect 163838 604840 163839 604841
rect 164537 604840 164538 604841
rect 163837 604839 163838 604840
rect 164538 604839 164539 604840
rect 163837 604240 163838 604241
rect 164538 604240 164539 604241
rect 163838 604239 163839 604240
rect 164537 604239 164538 604240
rect 164550 604228 164584 604852
rect 164596 604840 164597 604841
rect 165295 604840 165296 604841
rect 164595 604839 164596 604840
rect 165296 604839 165297 604840
rect 164595 604240 164596 604241
rect 165296 604240 165297 604241
rect 164596 604239 164597 604240
rect 165295 604239 165296 604240
rect 165308 604228 165342 604852
rect 165354 604840 165355 604841
rect 166053 604840 166054 604841
rect 165353 604839 165354 604840
rect 166054 604839 166055 604840
rect 165353 604240 165354 604241
rect 166054 604240 166055 604241
rect 165354 604239 165355 604240
rect 166053 604239 166054 604240
rect 166066 604228 166100 604852
rect 166112 604840 166113 604841
rect 166811 604840 166812 604841
rect 166111 604839 166112 604840
rect 166812 604839 166813 604840
rect 166111 604240 166112 604241
rect 166812 604240 166813 604241
rect 166112 604239 166113 604240
rect 166811 604239 166812 604240
rect 166824 604228 166858 604852
rect 166870 604840 166871 604841
rect 167569 604840 167570 604841
rect 166869 604839 166870 604840
rect 167570 604839 167571 604840
rect 166869 604240 166870 604241
rect 167570 604240 167571 604241
rect 166870 604239 166871 604240
rect 167569 604239 167570 604240
rect 167582 604228 167616 604852
rect 167628 604840 167629 604841
rect 167627 604839 167628 604840
rect 167756 604824 167828 604862
rect 167794 604256 167828 604824
rect 167627 604240 167628 604241
rect 167628 604239 167629 604240
rect 167744 604228 167755 604239
rect 159646 604166 159718 604204
rect 159768 604194 167755 604228
rect 159989 604182 159990 604183
rect 159990 604181 159991 604182
rect 159684 603598 159718 604166
rect 159990 603582 159991 603583
rect 159989 603581 159990 603582
rect 160002 603570 160036 604194
rect 160048 604182 160049 604183
rect 160747 604182 160748 604183
rect 160047 604181 160048 604182
rect 160748 604181 160749 604182
rect 160047 603582 160048 603583
rect 160748 603582 160749 603583
rect 160048 603581 160049 603582
rect 160747 603581 160748 603582
rect 160760 603570 160794 604194
rect 160806 604182 160807 604183
rect 161505 604182 161506 604183
rect 160805 604181 160806 604182
rect 161506 604181 161507 604182
rect 160805 603582 160806 603583
rect 161506 603582 161507 603583
rect 160806 603581 160807 603582
rect 161505 603581 161506 603582
rect 161518 603570 161552 604194
rect 161564 604182 161565 604183
rect 162263 604182 162264 604183
rect 161563 604181 161564 604182
rect 162264 604181 162265 604182
rect 161563 603582 161564 603583
rect 162264 603582 162265 603583
rect 161564 603581 161565 603582
rect 162263 603581 162264 603582
rect 162276 603570 162310 604194
rect 162322 604182 162323 604183
rect 163021 604182 163022 604183
rect 162321 604181 162322 604182
rect 163022 604181 163023 604182
rect 162321 603582 162322 603583
rect 163022 603582 163023 603583
rect 162322 603581 162323 603582
rect 163021 603581 163022 603582
rect 163034 603570 163068 604194
rect 163080 604182 163081 604183
rect 163779 604182 163780 604183
rect 163079 604181 163080 604182
rect 163780 604181 163781 604182
rect 163684 603602 163694 603668
rect 163712 603630 163722 603668
rect 163079 603582 163080 603583
rect 163780 603582 163781 603583
rect 163080 603581 163081 603582
rect 163779 603581 163780 603582
rect 163792 603570 163826 604194
rect 163838 604182 163839 604183
rect 164537 604182 164538 604183
rect 163837 604181 163838 604182
rect 164538 604181 164539 604182
rect 163837 603582 163838 603583
rect 164538 603582 164539 603583
rect 163838 603581 163839 603582
rect 164537 603581 164538 603582
rect 164550 603570 164584 604194
rect 164596 604182 164597 604183
rect 165295 604182 165296 604183
rect 164595 604181 164596 604182
rect 165296 604181 165297 604182
rect 164595 603582 164596 603583
rect 164596 603581 164597 603582
rect 165260 603580 165302 603604
rect 165232 603570 165302 603576
rect 165308 603570 165342 604194
rect 165354 604182 165355 604183
rect 166053 604182 166054 604183
rect 165353 604181 165354 604182
rect 166054 604181 166055 604182
rect 165348 603580 165384 603604
rect 166054 603582 166055 603583
rect 166053 603581 166054 603582
rect 165348 603570 165412 603576
rect 166066 603570 166100 604194
rect 166112 604182 166113 604183
rect 166811 604182 166812 604183
rect 166111 604181 166112 604182
rect 166812 604181 166813 604182
rect 166111 603582 166112 603583
rect 166812 603582 166813 603583
rect 166112 603581 166113 603582
rect 166811 603581 166812 603582
rect 166824 603570 166858 604194
rect 166870 604182 166871 604183
rect 167569 604182 167570 604183
rect 166869 604181 166870 604182
rect 167570 604181 167571 604182
rect 166869 603582 166870 603583
rect 167570 603582 167571 603583
rect 166870 603581 166871 603582
rect 167569 603581 167570 603582
rect 167582 603570 167616 604194
rect 167628 604182 167629 604183
rect 167627 604181 167628 604182
rect 167756 604166 167828 604204
rect 167794 603598 167828 604166
rect 167627 603582 167628 603583
rect 167628 603581 167629 603582
rect 167744 603570 167755 603581
rect 159768 603536 167755 603570
rect 160002 603456 160036 603536
rect 160760 603456 160794 603536
rect 161518 603456 161552 603536
rect 162276 603456 162310 603536
rect 163034 603456 163068 603536
rect 163792 603456 163826 603536
rect 164550 603456 164584 603536
rect 165308 603456 165342 603536
rect 166066 603456 166100 603536
rect 166824 603456 166858 603536
rect 167582 603456 167616 603536
rect 167896 603456 167930 605214
rect 170606 605180 170636 605282
rect 171480 605248 171514 605316
rect 171558 605268 171576 605282
rect 171530 605248 171576 605254
rect 171582 605248 171616 605316
rect 172102 605282 172140 605286
rect 172860 605282 172898 605286
rect 171622 605268 172142 605282
rect 172152 605268 172900 605282
rect 172102 605254 172140 605268
rect 172860 605254 172898 605268
rect 171622 605248 172140 605254
rect 171480 605214 172140 605248
rect 172180 605240 172898 605254
rect 172192 605214 172898 605240
rect 170632 603714 170648 604232
rect 170670 603752 170686 604194
rect 159582 603422 167930 603456
rect 163034 601939 163068 603422
rect 163668 603088 163694 603118
rect 163696 603116 163722 603118
rect 163758 603116 163782 603118
rect 163786 603088 163810 603118
rect 171480 603082 171514 605214
rect 171582 605198 171616 605214
rect 171654 605176 172118 605182
rect 172176 605176 172876 605182
rect 173002 605170 173036 605316
rect 171544 605108 171616 605146
rect 171666 605136 173036 605170
rect 172117 605124 172118 605125
rect 172118 605123 172119 605124
rect 171582 604540 171616 605108
rect 172118 604524 172119 604525
rect 172117 604523 172118 604524
rect 172130 604512 172164 605136
rect 172176 605124 172177 605125
rect 172875 605124 172876 605125
rect 172175 605123 172176 605124
rect 172876 605123 172877 605124
rect 172175 604524 172176 604525
rect 172876 604524 172877 604525
rect 172176 604523 172177 604524
rect 172875 604523 172876 604524
rect 172888 604512 172922 605136
rect 173002 604512 173036 605136
rect 171544 604450 171616 604488
rect 171666 604478 173036 604512
rect 172117 604466 172118 604467
rect 172118 604465 172119 604466
rect 171582 603882 171616 604450
rect 172118 603866 172119 603867
rect 172117 603865 172118 603866
rect 172130 603854 172164 604478
rect 172176 604466 172177 604467
rect 172875 604466 172876 604467
rect 172175 604465 172176 604466
rect 172876 604465 172877 604466
rect 172175 603866 172176 603867
rect 172876 603866 172877 603867
rect 172176 603865 172177 603866
rect 172875 603865 172876 603866
rect 172888 603854 172922 604478
rect 173002 603854 173036 604478
rect 171544 603792 171616 603830
rect 171666 603820 173036 603854
rect 172117 603808 172118 603809
rect 172118 603807 172119 603808
rect 171582 603224 171616 603792
rect 172118 603208 172119 603209
rect 172117 603207 172118 603208
rect 172130 603196 172164 603820
rect 172176 603808 172177 603809
rect 172875 603808 172876 603809
rect 172175 603807 172176 603808
rect 172876 603807 172877 603808
rect 172175 603208 172176 603209
rect 172876 603208 172877 603209
rect 172176 603207 172177 603208
rect 172875 603207 172876 603208
rect 172888 603196 172922 603820
rect 173002 603196 173036 603820
rect 171666 603178 173036 603196
rect 189279 605021 189327 606523
rect 189407 606533 189441 606585
rect 190065 606564 190099 606585
rect 190723 606564 190757 606585
rect 191381 606564 191415 606585
rect 192039 606564 192073 606585
rect 192697 606564 192731 606585
rect 190023 606533 190099 606564
rect 190681 606533 190757 606564
rect 191339 606533 191415 606564
rect 191997 606533 192073 606564
rect 189407 606436 189453 606533
rect 190023 606517 190111 606533
rect 190681 606517 190769 606533
rect 191339 606517 191427 606533
rect 191997 606517 192085 606533
rect 192655 606517 192731 606564
rect 192811 606523 192845 609538
rect 194364 609566 194398 611408
rect 194466 611346 194512 611498
rect 195064 611454 195090 612574
rect 195092 611454 195118 612546
rect 195136 611498 195202 613110
rect 195794 611498 195860 613110
rect 195136 611486 195170 611498
rect 195794 611486 195828 611498
rect 195124 611448 195174 611486
rect 195228 611454 195246 611470
rect 195782 611448 195832 611486
rect 196384 611454 196400 612556
rect 196412 611454 196428 612528
rect 196452 611498 196518 613110
rect 197110 611498 197176 613110
rect 197208 611752 197214 613154
rect 197236 611724 197242 613154
rect 197757 613110 197788 613121
rect 197800 613110 197834 613262
rect 196452 611486 196486 611498
rect 197110 611486 197144 611498
rect 196440 611448 196490 611486
rect 197098 611448 197148 611486
rect 197692 611454 197716 612558
rect 197720 611454 197744 612530
rect 197768 611498 197834 613110
rect 197882 613200 197900 613262
rect 197914 613200 197948 613502
rect 197768 611486 197802 611498
rect 197756 611448 197806 611486
rect 194572 611414 195174 611448
rect 195230 611414 195832 611448
rect 195888 611414 196490 611448
rect 196546 611414 197148 611448
rect 197204 611414 197806 611448
rect 195124 611398 195170 611414
rect 195782 611398 195828 611414
rect 196440 611398 196486 611414
rect 197098 611398 197144 611414
rect 197756 611398 197802 611414
rect 197882 611408 197948 613200
rect 198502 612136 198622 612156
rect 198808 612138 199048 612690
rect 198808 612136 199098 612138
rect 198496 612108 198650 612128
rect 198808 612110 199048 612136
rect 198808 612108 199126 612110
rect 198808 612052 199048 612108
rect 195136 611346 195170 611398
rect 194466 611312 197814 611346
rect 195136 609566 195170 611312
rect 197104 609566 197126 609756
rect 197882 609566 197916 611408
rect 205870 610080 205872 610130
rect 205898 610080 205900 610158
rect 205318 609840 205956 610080
rect 211084 610036 211086 610114
rect 211112 610036 211114 610086
rect 211028 609796 211666 610036
rect 194364 609538 197916 609566
rect 194058 609096 194060 609144
rect 194030 609068 194060 609088
rect 194364 606528 194398 609538
rect 195136 609510 195170 609538
rect 197104 609510 197126 609538
rect 194436 609482 197854 609510
rect 194478 606624 194512 606658
rect 195136 606624 195170 609482
rect 197104 609088 197126 609482
rect 195828 606826 195834 607900
rect 195828 606658 195860 606826
rect 195794 606624 195860 606658
rect 195884 606624 195888 606854
rect 196452 606624 196486 606658
rect 197046 606624 197072 606818
rect 197104 606790 197128 607900
rect 197074 606658 197128 606790
rect 197074 606624 197144 606658
rect 197768 606624 197802 606658
rect 194446 606590 197836 606624
rect 189455 606483 190111 606517
rect 190113 606483 190769 606517
rect 190771 606483 191427 606517
rect 191429 606483 192085 606517
rect 192087 606483 192731 606517
rect 190031 606477 190035 606483
rect 190059 606449 190063 606483
rect 190065 606436 190111 606483
rect 190723 606436 190769 606483
rect 191347 606477 191351 606483
rect 191375 606449 191379 606483
rect 191381 606436 191427 606483
rect 192039 606436 192085 606483
rect 192663 606477 192667 606483
rect 192691 606449 192695 606483
rect 189407 606424 189441 606436
rect 190040 606424 190053 606435
rect 190065 606424 190099 606436
rect 190698 606424 190711 606435
rect 190723 606424 190757 606436
rect 191356 606424 191369 606435
rect 191381 606424 191415 606436
rect 192014 606424 192027 606435
rect 192039 606424 192073 606436
rect 192672 606424 192685 606435
rect 192697 606424 192731 606483
rect 189393 605120 189441 606424
rect 190051 605120 190099 606424
rect 190709 605120 190757 606424
rect 171650 603162 173160 603178
rect 172130 603144 172164 603162
rect 172888 603144 172922 603162
rect 173002 603144 173036 603162
rect 171616 603128 173126 603144
rect 172130 603082 172164 603128
rect 172888 603082 172922 603128
rect 173002 603082 173036 603128
rect 163274 603006 163596 603078
rect 171480 603048 175456 603082
rect 163076 602544 163714 603006
rect 163764 602918 164312 602952
rect 163764 602636 163798 602918
rect 163939 602838 164137 602849
rect 163828 602794 163938 602832
rect 163950 602804 164137 602838
rect 164138 602794 164248 602832
rect 163866 602760 163938 602794
rect 163939 602750 164137 602761
rect 164176 602760 164248 602794
rect 163950 602716 164137 602750
rect 164278 602636 164312 602918
rect 163764 602602 164312 602636
rect 165274 602596 165292 602796
rect 165302 602568 165320 602824
rect 159551 601606 167989 601939
rect 146208 601572 146297 601606
rect 146346 601583 172934 601606
rect 173002 601583 173036 603048
rect 146346 601572 173036 601583
rect 146208 600464 146279 601572
rect 146358 600604 146392 601572
rect 147116 601542 147150 601572
rect 147762 601542 147796 601572
rect 147874 601542 147910 601572
rect 147920 601542 147921 601572
rect 148534 601542 148579 601572
rect 148632 601542 148677 601572
rect 149192 601542 149237 601572
rect 149390 601542 149435 601572
rect 149850 601542 149895 601572
rect 150148 601542 150193 601572
rect 150508 601542 150553 601572
rect 150906 601542 150951 601572
rect 151166 601542 151211 601572
rect 151280 601542 151314 601572
rect 151664 601542 151698 601572
rect 152422 601542 152456 601572
rect 153180 601542 153214 601572
rect 153938 601542 153972 601572
rect 154696 601542 154730 601572
rect 155454 601542 155488 601572
rect 156212 601542 156246 601572
rect 156970 601542 157004 601572
rect 157728 601542 157762 601572
rect 157772 601542 157796 601568
rect 158486 601542 158520 601572
rect 159244 601542 159278 601572
rect 159551 601542 167989 601572
rect 168340 601542 168374 601572
rect 169098 601542 169132 601572
rect 169856 601542 169890 601572
rect 170614 601542 170648 601572
rect 171372 601542 171406 601572
rect 173002 601565 173036 601572
rect 146938 601504 147676 601542
rect 147762 601504 151360 601542
rect 151636 601504 151698 601542
rect 152394 601504 152456 601542
rect 153152 601504 153214 601542
rect 153910 601504 153972 601542
rect 154668 601504 154730 601542
rect 155426 601504 155488 601542
rect 156184 601504 156246 601542
rect 156942 601504 157004 601542
rect 157700 601504 167989 601542
rect 168312 601504 168374 601542
rect 169070 601504 169132 601542
rect 169828 601504 169890 601542
rect 170586 601504 170648 601542
rect 171344 601538 171406 601542
rect 171344 601510 171412 601538
rect 171338 601504 171412 601510
rect 171421 601504 173072 601565
rect 146404 601470 147150 601504
rect 147178 601470 147910 601504
rect 147116 600604 147150 601470
rect 146358 600566 146432 600604
rect 147088 600566 147150 600604
rect 147762 600566 147796 601470
rect 147874 600604 147910 601470
rect 147846 600566 147910 600604
rect 146358 600464 146392 600566
rect 146420 600532 147150 600566
rect 147162 600532 147910 600566
rect 147116 600464 147150 600532
rect 147762 600464 147796 600532
rect 147874 600464 147910 600532
rect 147920 600566 147921 601504
rect 147936 601470 148677 601504
rect 148694 601470 149435 601504
rect 149452 601470 150193 601504
rect 150210 601470 150951 601504
rect 150968 601470 151698 601504
rect 151710 601470 152456 601504
rect 152468 601470 153214 601504
rect 153226 601470 153972 601504
rect 153984 601470 154730 601504
rect 154742 601470 155488 601504
rect 155500 601470 156246 601504
rect 156258 601470 157004 601504
rect 157016 601470 157762 601504
rect 148534 600628 148579 601470
rect 148632 600628 148677 601470
rect 148534 600566 148568 600628
rect 148632 600604 148666 600628
rect 149192 600604 149237 601470
rect 149390 600604 149435 601470
rect 149850 600604 149895 601470
rect 150148 600604 150193 601470
rect 148604 600566 148666 600604
rect 149188 600566 150193 600604
rect 150508 600816 150553 601470
rect 150906 600816 150951 601470
rect 150508 600566 150542 600816
rect 150906 600604 150940 600816
rect 150966 600800 150974 600816
rect 150878 600566 150940 600604
rect 151166 600790 151211 601470
rect 151166 600566 151200 600790
rect 151280 600566 151314 601470
rect 151664 601466 151698 601470
rect 152422 601466 152456 601470
rect 153180 601466 153214 601470
rect 153938 601466 153972 601470
rect 154696 601466 154730 601470
rect 151452 601436 155130 601466
rect 151664 600604 151698 601436
rect 152422 600604 152456 601436
rect 153180 600604 153214 601436
rect 153938 600604 153972 601436
rect 154696 600604 154730 601436
rect 155454 600604 155488 601470
rect 156212 600604 156246 601470
rect 156970 600604 157004 601470
rect 157728 600604 157762 601470
rect 157772 601470 158520 601504
rect 158548 601470 159278 601504
rect 159306 601470 168374 601504
rect 168386 601470 169132 601504
rect 169144 601470 169890 601504
rect 169902 601470 170648 601504
rect 170660 601470 171412 601504
rect 171418 601470 173072 601504
rect 157772 600604 157796 601470
rect 158486 600604 158520 601470
rect 159244 600604 159278 601470
rect 159551 600604 167989 601470
rect 168340 600604 168374 601470
rect 169098 600604 169132 601470
rect 169856 600604 169890 601470
rect 170614 600604 170648 601470
rect 171338 601464 171356 601470
rect 171366 601436 171412 601470
rect 171372 600604 171406 601436
rect 151428 600566 155188 600604
rect 155426 600600 155488 600604
rect 155426 600572 155494 600600
rect 155420 600566 155494 600572
rect 155504 600566 155522 600572
rect 156184 600566 156246 600604
rect 156942 600600 157004 600604
rect 156942 600572 157010 600600
rect 156936 600566 157010 600572
rect 157020 600566 157038 600572
rect 157700 600566 167989 600604
rect 168312 600566 168374 600604
rect 169070 600566 169132 600604
rect 169828 600566 169890 600604
rect 170586 600566 170648 600604
rect 171344 600566 171406 600604
rect 171421 600566 173072 601470
rect 147920 600532 148666 600566
rect 148678 600532 149435 600566
rect 149452 600532 150193 600566
rect 150210 600532 150940 600566
rect 150952 600532 151698 600566
rect 151726 600532 152462 600566
rect 147920 600464 147921 600532
rect 148534 600464 148568 600532
rect 148632 600464 148666 600532
rect 149192 600464 149237 600532
rect 149390 600464 149435 600532
rect 149850 600464 149895 600532
rect 150148 600464 150193 600532
rect 150508 600464 150542 600532
rect 150906 600464 150940 600532
rect 151166 600464 151200 600532
rect 151280 600464 151314 600532
rect 151664 600464 151698 600532
rect 152388 600526 152406 600532
rect 152416 600498 152462 600532
rect 152472 600532 153214 600566
rect 153242 600532 153978 600566
rect 152472 600526 152490 600532
rect 152422 600464 152456 600498
rect 153180 600464 153214 600532
rect 153904 600526 153922 600532
rect 153932 600498 153978 600532
rect 153988 600532 154730 600566
rect 154758 600532 155494 600566
rect 155500 600532 156246 600566
rect 156258 600532 157010 600566
rect 157016 600532 157762 600566
rect 153988 600526 154006 600532
rect 153938 600464 153972 600498
rect 154696 600464 154730 600532
rect 155420 600526 155438 600532
rect 155448 600498 155494 600532
rect 155504 600526 155522 600532
rect 155454 600464 155488 600498
rect 156212 600464 156246 600532
rect 156936 600526 156954 600532
rect 156964 600498 157010 600532
rect 157020 600526 157038 600532
rect 156970 600464 157004 600498
rect 157728 600464 157762 600532
rect 157772 600532 158526 600566
rect 157772 600464 157796 600532
rect 158452 600526 158470 600532
rect 158480 600498 158526 600532
rect 158536 600532 159278 600566
rect 159306 600532 168374 600566
rect 168386 600532 169132 600566
rect 169144 600532 169890 600566
rect 169902 600532 170648 600566
rect 170660 600532 171406 600566
rect 171418 600532 173072 600566
rect 158536 600526 158554 600532
rect 158486 600464 158520 600498
rect 159244 600464 159278 600532
rect 159551 600464 167989 600532
rect 168340 600464 168374 600532
rect 169098 600464 169132 600532
rect 169856 600464 169890 600532
rect 170614 600464 170648 600532
rect 171372 600464 171406 600532
rect 171421 600464 173072 600532
rect 146208 600430 146297 600464
rect 146340 600430 173072 600464
rect 146208 600186 146279 600430
rect 146140 599944 146178 600130
rect 146196 599944 146279 600186
rect 142793 599617 146163 599651
rect 124842 594597 129196 594662
rect 131644 594597 133262 594692
rect 124842 593884 133262 594597
rect 134446 593934 134502 593946
rect 135690 593934 135746 593946
rect 134446 593884 134502 593890
rect 124842 593850 135136 593884
rect 135690 593878 135746 593890
rect 136288 593850 142222 595752
rect 124842 593836 133262 593850
rect 124842 593834 133428 593836
rect 100480 593498 100486 593640
rect 100474 593476 100486 593498
rect 113168 593492 113468 593511
rect 114820 593492 116320 593511
rect 117888 593505 119596 593511
rect 119606 593505 119640 593764
rect 119720 593505 119754 593764
rect 119958 593550 120014 593567
rect 121215 593533 121249 593764
rect 119765 593517 119766 593518
rect 119766 593516 119767 593517
rect 119884 593505 120014 593511
rect 121156 593505 121167 593516
rect 117888 593494 121167 593505
rect 100470 593450 100486 593476
rect 119572 593471 121167 593494
rect 100470 593420 100496 593450
rect 113412 593366 114876 593382
rect 100470 593316 100496 593344
rect 100470 593288 100492 593316
rect 100474 593280 100492 593288
rect 97364 593156 98828 593172
rect 96136 593027 96192 593044
rect 96538 593027 97420 593044
rect 98772 593027 99072 593044
rect 96136 592971 96192 592988
rect 100480 592822 100492 593280
rect 96468 592624 99291 592774
rect 96468 592590 104666 592624
rect 96468 591751 99291 592590
rect 100466 592584 100536 592586
rect 100522 592528 100536 592530
rect 100604 591976 100976 592004
rect 100566 591938 101014 591966
rect 94816 591717 99291 591751
rect 96468 591567 99291 591717
rect 94892 590844 94894 590986
rect 94882 590822 94894 590844
rect 94878 590796 94894 590822
rect 94878 590766 94904 590796
rect 95596 590696 95628 590766
rect 94878 590662 94904 590690
rect 95630 590662 95662 590800
rect 94878 590634 94900 590662
rect 94882 590626 94900 590634
rect 94892 590168 94900 590626
rect 96504 590084 96538 591567
rect 96980 591336 98382 591350
rect 112985 590485 113019 593342
rect 116510 593314 117076 593348
rect 116510 592992 116544 593314
rect 117042 593250 117076 593314
rect 117126 593250 117746 593366
rect 116694 593234 116892 593245
rect 116565 593172 116693 593219
rect 116705 593200 116892 593234
rect 116978 593219 117746 593250
rect 116893 593172 117746 593219
rect 116612 593134 116693 593172
rect 116940 593134 117746 593172
rect 116694 593106 116892 593117
rect 116950 593108 117746 593134
rect 116705 593072 116892 593106
rect 116978 593038 117746 593108
rect 117042 592992 117076 593038
rect 116510 592958 117076 592992
rect 117126 592944 117746 593038
rect 119606 592847 119640 593471
rect 119720 592847 119754 593471
rect 119766 593459 119767 593460
rect 119765 593458 119766 593459
rect 121168 593443 121249 593490
rect 119958 592934 120014 592936
rect 119958 592878 120014 592880
rect 121215 592875 121249 593443
rect 119765 592859 119766 592860
rect 119766 592858 119767 592859
rect 121156 592847 121167 592858
rect 119572 592813 121167 592847
rect 119606 592638 119640 592813
rect 119720 592799 119754 592813
rect 119766 592801 119767 592802
rect 119765 592800 119766 592801
rect 121168 592787 121296 592832
rect 121167 592786 121168 592787
rect 119742 592772 120014 592774
rect 119770 592744 120014 592746
rect 119958 592740 120014 592744
rect 121215 592740 121249 592785
rect 121317 592740 121351 593764
rect 124842 593390 133262 593834
rect 119782 592706 121351 592740
rect 121215 592638 121249 592706
rect 121317 592638 121351 592706
rect 124855 592740 124889 593390
rect 124957 593159 124991 593390
rect 125824 593143 125825 593144
rect 125823 593142 125824 593143
rect 125484 593131 125830 593137
rect 125836 593131 125870 593390
rect 128894 593230 128928 593390
rect 125881 593143 125882 593144
rect 125882 593142 125883 593143
rect 125876 593131 126166 593137
rect 128318 593131 128536 593142
rect 128860 593137 128866 593230
rect 128882 593143 128883 593144
rect 128881 593142 128882 593143
rect 128888 593137 128928 593230
rect 128894 593131 128928 593137
rect 129008 593131 129042 593390
rect 124910 593069 124991 593116
rect 125050 593097 129042 593131
rect 129886 593118 131386 593137
rect 131680 593131 131714 593390
rect 131782 593254 131816 593390
rect 133085 593239 133119 593390
rect 133038 593238 133119 593239
rect 133038 593226 133135 593238
rect 131735 593164 131816 593211
rect 131875 593192 133135 593226
rect 132738 593180 133135 593192
rect 132738 593174 133119 593180
rect 131782 593144 131816 593164
rect 133079 593159 133119 593174
rect 133079 593148 133094 593159
rect 133079 593147 133125 593148
rect 131646 593097 131714 593131
rect 131735 593143 131816 593144
rect 131735 593131 131863 593143
rect 133026 593137 133037 593142
rect 132738 593131 133038 593137
rect 131735 593120 133038 593131
rect 133187 593120 133221 593390
rect 135690 593274 135746 593288
rect 135690 593218 135746 593232
rect 134446 593174 134502 593176
rect 131735 593119 134502 593120
rect 131735 593118 133079 593119
rect 133125 593118 134502 593119
rect 131735 593097 133037 593118
rect 125823 593085 125824 593086
rect 125824 593084 125825 593085
rect 124957 592740 124991 593069
rect 125836 592799 125870 593097
rect 128894 593091 128928 593097
rect 125882 593085 125883 593086
rect 125881 593084 125882 593085
rect 128860 593008 128866 593091
rect 128881 593085 128882 593086
rect 128882 593084 128883 593085
rect 128888 593008 128928 593091
rect 128894 592992 128928 593008
rect 129008 592992 129042 593097
rect 131680 593008 131714 593097
rect 131766 593085 131863 593097
rect 131330 592992 131776 593008
rect 128460 592876 129080 592992
rect 129130 592940 129696 592974
rect 129130 592876 129164 592940
rect 128460 592845 129228 592876
rect 129501 592860 129512 592871
rect 125037 592787 125038 592788
rect 128460 592787 129266 592845
rect 129325 592826 129512 592860
rect 129513 592798 129594 592845
rect 125038 592786 125039 592787
rect 125808 592740 125855 592787
rect 128318 592760 129266 592787
rect 129560 592760 129594 592798
rect 128318 592740 129256 592760
rect 124855 592706 125855 592740
rect 125898 592734 129256 592740
rect 125898 592706 129228 592734
rect 129501 592732 129512 592743
rect 124855 592638 124889 592706
rect 124957 592638 124991 592706
rect 128460 592664 129228 592706
rect 129325 592698 129512 592732
rect 128460 592638 129080 592664
rect 119606 592604 129080 592638
rect 116986 592392 117434 592604
rect 117078 592382 117210 592392
rect 113060 592270 121276 592281
rect 113071 592258 121265 592270
rect 113060 592247 121276 592258
rect 113087 592201 113121 592247
rect 113996 592189 114452 592208
rect 121215 592201 121249 592247
rect 113180 592143 121156 592189
rect 113180 592133 121167 592143
rect 113087 591537 113121 592127
rect 114034 592118 114490 592133
rect 121215 591984 121249 592127
rect 121317 591984 121351 592604
rect 124855 591984 124889 592604
rect 128460 592570 129080 592604
rect 129130 592618 129164 592664
rect 129662 592618 129696 592940
rect 129130 592584 129696 592618
rect 126110 592504 126764 592506
rect 131680 592454 131714 592992
rect 131782 592596 131816 593085
rect 133038 593069 133119 593116
rect 133085 592581 133119 593069
rect 133038 592580 133119 592581
rect 133038 592568 133135 592580
rect 131875 592537 133135 592568
rect 131875 592534 133150 592537
rect 133038 592522 133150 592534
rect 131742 592454 133026 592488
rect 133085 592485 133119 592488
rect 133187 592454 133221 593118
rect 134446 592614 134502 592630
rect 135690 592614 135746 592630
rect 134446 592558 134502 592574
rect 135690 592558 135746 592574
rect 131680 592420 135136 592454
rect 128772 592018 129220 592230
rect 133187 592026 133221 592420
rect 128996 592008 129128 592018
rect 131680 591992 135136 592026
rect 119642 591950 129078 591984
rect 116986 591928 117434 591938
rect 116978 591726 117434 591928
rect 116978 591716 117426 591726
rect 119642 591542 119676 591950
rect 121215 591882 121249 591950
rect 121317 591882 121351 591950
rect 119818 591848 121351 591882
rect 121167 591801 121168 591802
rect 121168 591800 121169 591801
rect 119745 591789 119790 591800
rect 116120 591531 119676 591542
rect 119756 591552 119790 591789
rect 120036 591602 120092 591628
rect 119756 591531 120440 591552
rect 121156 591531 121167 591542
rect 121215 591537 121249 591848
rect 113180 591475 121167 591531
rect 113087 591447 113121 591451
rect 119642 591417 119676 591475
rect 119756 591417 119790 591475
rect 119802 591463 119803 591464
rect 119801 591462 119802 591463
rect 119806 591454 120460 591475
rect 120036 591438 120092 591454
rect 121168 591447 121249 591494
rect 121215 591430 121249 591447
rect 121168 591417 121249 591430
rect 121317 591417 121351 591848
rect 124855 591907 124889 591950
rect 124928 591907 124951 591944
rect 124997 591907 125312 591944
rect 126170 591916 128702 591944
rect 126136 591907 128942 591916
rect 129044 591907 129078 591950
rect 131680 591907 131714 591992
rect 131720 591912 132788 591922
rect 133038 591912 133150 591924
rect 131720 591909 133150 591912
rect 131720 591907 133135 591909
rect 133187 591907 133221 591992
rect 124855 591873 133221 591907
rect 124855 591849 125891 591873
rect 125934 591854 128949 591873
rect 125918 591849 128949 591854
rect 124855 591848 128949 591849
rect 113049 591383 121351 591417
rect 119642 590851 119676 591383
rect 119756 590851 119790 591383
rect 120036 591382 120092 591383
rect 120036 590886 120092 590913
rect 121215 590879 121249 591383
rect 119801 590863 119802 590864
rect 119802 590862 119803 590863
rect 120036 590851 120092 590857
rect 121156 590851 121167 590862
rect 119608 590817 121167 590851
rect 113412 590712 114876 590728
rect 119642 590485 119676 590817
rect 119756 590485 119790 590817
rect 119802 590805 119803 590806
rect 119801 590804 119802 590805
rect 121168 590789 121249 590836
rect 121215 590490 121249 590789
rect 112189 590451 120459 590485
rect 94816 590050 99260 590084
rect 96504 589970 96538 590050
rect 96606 590004 96640 590050
rect 99226 589992 99260 590050
rect 96690 589970 99260 589992
rect 96470 589958 99260 589970
rect 96470 589946 99074 589958
rect 96470 589936 99085 589946
rect 94874 589930 94948 589932
rect 94930 589874 94948 589876
rect 96504 589312 96538 589936
rect 96568 589930 96678 589936
rect 96590 589924 96678 589930
rect 96606 589362 96640 589924
rect 99086 589908 99158 589946
rect 99124 589346 99158 589908
rect 99086 589334 99174 589346
rect 99226 589334 99260 589958
rect 96690 589312 99260 589334
rect 96504 589300 99260 589312
rect 96504 589278 99074 589300
rect 96504 589220 96538 589278
rect 99124 589250 99158 589254
rect 99226 589220 99260 589300
rect 96504 589186 104756 589220
rect 99226 588851 99260 589186
rect 96463 588646 99296 588851
rect 94816 588620 99296 588646
rect 92742 587344 92754 587374
rect 92770 587344 92782 587402
rect 92742 587266 92754 587298
rect 92770 587238 92782 587298
rect 96463 586496 99296 588620
rect 96499 586161 96533 586496
rect 104688 586356 104901 588851
rect 104688 586345 105797 586356
rect 104688 586333 105786 586345
rect 104688 586322 105797 586333
rect 104688 586253 104901 586322
rect 104688 586242 105697 586253
rect 91634 586148 92308 586161
rect 91003 586127 92308 586148
rect 94816 586127 99273 586161
rect 91018 585985 91638 586127
rect 91688 586093 92222 586112
rect 91722 586078 92220 586093
rect 91009 585946 91638 585985
rect 90936 585860 91638 585946
rect 91009 585708 91638 585860
rect 91688 586053 92254 586059
rect 91688 586047 91722 586053
rect 92220 586047 92254 586053
rect 96499 586047 96533 586127
rect 96601 586081 96635 586127
rect 99239 586069 99273 586127
rect 96554 586047 96635 586054
rect 96694 586047 99273 586069
rect 91688 586044 92254 586047
rect 91688 585972 91722 586044
rect 91845 586032 92097 586036
rect 91833 586013 92109 586032
rect 92059 585998 92070 586001
rect 91867 585983 92075 585998
rect 91743 585972 91824 585983
rect 91867 585979 92152 585983
rect 91688 585930 91728 585972
rect 91736 585936 91824 585972
rect 91883 585964 92070 585979
rect 92071 585936 92152 585979
rect 91736 585930 91756 585936
rect 91688 585756 91722 585930
rect 91790 585898 91824 585936
rect 92118 585898 92152 585936
rect 92059 585870 92070 585881
rect 91883 585836 92070 585870
rect 92220 585756 92254 586044
rect 96465 586035 99273 586047
rect 96465 586023 99078 586035
rect 96465 586013 99089 586023
rect 91688 585722 92254 585756
rect 91009 585654 91043 585708
rect 91009 585417 91638 585654
rect 91018 585232 91638 585417
rect 91688 585602 92254 585636
rect 91688 585389 91722 585602
rect 92059 585522 92070 585533
rect 91736 585395 91738 585482
rect 91743 585460 91824 585507
rect 91883 585488 92070 585522
rect 92071 585460 92152 585507
rect 91790 585406 91824 585460
rect 92118 585423 92152 585460
rect 92110 585414 92162 585423
rect 92112 585410 92158 585414
rect 92118 585406 92152 585410
rect 91872 585401 92070 585405
rect 91883 585389 92059 585394
rect 92082 585389 92190 585395
rect 92220 585389 92254 585602
rect 91688 585355 92254 585389
rect 91688 585280 91722 585355
rect 92220 585280 92254 585355
rect 91688 585246 92254 585280
rect 96499 585389 96533 586013
rect 96554 586007 96682 586013
rect 96585 586001 96682 586007
rect 96601 585439 96635 586001
rect 99090 585985 99171 586032
rect 99137 585423 99171 585985
rect 99090 585411 99187 585423
rect 99239 585411 99273 586035
rect 96694 585389 99273 585411
rect 96499 585377 99273 585389
rect 96499 585355 99078 585377
rect 99090 585365 99218 585374
rect 96499 585297 96533 585355
rect 99137 585327 99171 585331
rect 99239 585297 99273 585377
rect 104688 585297 104901 586242
rect 104910 586208 105697 586242
rect 96499 585263 104901 585297
rect 91516 584628 91716 584638
rect 91488 584600 91744 584610
rect 97382 584162 98846 584178
rect 96154 584033 96210 584050
rect 96556 584033 97438 584050
rect 98790 584033 99090 584050
rect 96154 583977 96210 583994
rect 99239 583780 99273 585263
rect 104688 585227 104901 585263
rect 100498 584504 100504 584646
rect 100492 584482 100504 584504
rect 100488 584456 100504 584482
rect 100488 584426 100514 584456
rect 100488 584322 100514 584350
rect 100488 584294 100510 584322
rect 100492 584286 100510 584294
rect 100498 583828 100510 584286
rect 96486 583744 99309 583780
rect 104724 583744 104758 585227
rect 104826 583744 104860 585227
rect 105686 583838 105697 583849
rect 104910 583804 105697 583838
rect 96486 583710 104774 583744
rect 104799 583737 104870 583744
rect 104779 583724 104870 583737
rect 105736 583724 105770 586322
rect 96486 583630 99309 583710
rect 96486 583596 104684 583630
rect 104690 583602 104700 583630
rect 104724 583602 104758 583710
rect 104779 583690 105804 583724
rect 104690 583596 104758 583602
rect 96486 582757 99309 583596
rect 100484 583590 100554 583592
rect 104700 583580 104758 583596
rect 104700 583568 104774 583580
rect 100540 583534 100554 583536
rect 104724 583498 104792 583568
rect 104810 583526 104826 583626
rect 104724 583050 104806 583498
rect 100622 582982 100994 583010
rect 104724 583000 104792 583050
rect 104810 583022 104834 583526
rect 104724 582988 104774 583000
rect 100584 582944 101032 582972
rect 104690 582944 104700 582972
rect 104724 582944 104758 582988
rect 104810 582984 104826 583022
rect 104690 582938 104758 582944
rect 104700 582922 104758 582938
rect 104700 582910 104774 582922
rect 94816 582723 99309 582757
rect 96486 582573 99309 582723
rect 104724 582846 104792 582910
rect 104810 582874 104826 582968
rect 104836 582874 104870 583690
rect 104810 582846 104870 582874
rect 94910 581850 94912 581992
rect 94900 581828 94912 581850
rect 94896 581802 94912 581828
rect 94896 581772 94922 581802
rect 95614 581702 95646 581772
rect 94896 581668 94922 581696
rect 95648 581668 95680 581806
rect 94896 581640 94918 581668
rect 94900 581632 94918 581640
rect 93356 581202 93508 581226
rect 93636 581216 93782 581224
rect 93614 581202 93782 581216
rect 93384 581174 93480 581198
rect 93064 581126 93098 581137
rect 93392 581126 93426 581137
rect 92926 581090 93564 581126
rect 93614 581090 93648 581202
rect 93664 581174 93754 581196
rect 93716 581104 93750 581137
rect 94026 581104 94060 581137
rect 94128 581090 94162 581216
rect 94336 581142 94340 581316
rect 94370 581176 94374 581350
rect 94910 581174 94918 581632
rect 96522 581090 96556 582573
rect 104724 582450 104870 582846
rect 105838 582450 105872 588914
rect 103516 582380 105908 582450
rect 96998 582342 98400 582356
rect 92926 581056 99278 581090
rect 92926 580908 93564 581056
rect 93710 580988 94066 581010
rect 93614 580962 94162 580988
rect 96522 580976 96556 581056
rect 96624 581038 96664 581056
rect 96618 581014 96664 581038
rect 96624 581010 96658 581014
rect 99244 580998 99278 581056
rect 96708 580976 99278 580998
rect 96488 580964 99278 580976
rect 96488 580952 99092 580964
rect 96488 580942 99103 580952
rect 91032 580330 91066 580362
rect 90998 580296 91100 580328
rect 96522 580318 96556 580942
rect 96586 580936 96696 580942
rect 96608 580930 96696 580936
rect 96624 580368 96658 580930
rect 99104 580914 99176 580952
rect 99142 580352 99176 580914
rect 99104 580340 99192 580352
rect 99244 580340 99278 580964
rect 96708 580318 99278 580340
rect 96522 580306 99278 580318
rect 96522 580284 99092 580306
rect 91540 579862 92720 580234
rect 96522 580226 96556 580284
rect 99142 580256 99176 580260
rect 99244 580226 99278 580306
rect 103516 581036 105918 582380
rect 103516 581000 105908 581036
rect 103516 580226 104906 581000
rect 96522 580192 104906 580226
rect 91406 579688 92808 579702
rect 95218 579660 95896 579752
rect 96664 579720 97212 579754
rect 96664 579692 96698 579720
rect 97178 579692 97212 579720
rect 96630 579660 96732 579692
rect 97144 579660 97246 579692
rect 97262 579660 97900 579808
rect 95218 579626 99092 579660
rect 95218 579418 95896 579626
rect 96546 579588 96632 579606
rect 94816 579276 95896 579418
rect 96664 579438 96698 579626
rect 96728 579596 96800 579626
rect 96850 579614 97026 579626
rect 96850 579606 97037 579614
rect 97038 579596 97110 579626
rect 96766 579562 96800 579596
rect 97068 579592 97072 579596
rect 97026 579552 97037 579563
rect 97076 579562 97110 579596
rect 96850 579518 97037 579552
rect 97068 579542 97072 579562
rect 97040 579514 97072 579534
rect 97178 579438 97212 579626
rect 96664 579404 97212 579438
rect 97262 579346 97900 579626
rect 94816 579206 95252 579276
rect 96664 579244 97212 579278
rect 96664 578962 96698 579244
rect 97026 579164 97037 579175
rect 96728 579120 96800 579158
rect 96850 579130 97037 579164
rect 97038 579120 97110 579158
rect 96766 579086 96800 579120
rect 96810 579086 97066 579110
rect 97076 579086 97110 579120
rect 97026 579082 97037 579086
rect 96838 579058 97038 579082
rect 96850 579042 97037 579058
rect 97178 578996 97212 579244
rect 96704 578968 97212 578996
rect 97178 578962 97212 578968
rect 96664 578928 97212 578962
rect 97262 578870 97900 579332
rect 97738 578850 97794 578870
rect 87549 578532 87757 578562
rect 99244 578549 99278 580192
rect 103516 580156 104906 580192
rect 87515 578498 87791 578528
rect 90894 578513 93129 578549
rect 97785 578518 99314 578549
rect 89161 578479 93129 578513
rect 85948 577208 87128 577580
rect 89065 576713 89099 578417
rect 89541 578411 89575 578449
rect 89672 578411 90852 578434
rect 90894 578411 93129 578479
rect 89241 578377 93129 578411
rect 89541 576713 89575 578377
rect 89672 578329 90852 578377
rect 89644 578318 90852 578329
rect 89655 578062 90852 578318
rect 89655 577098 89700 578062
rect 89837 577502 89882 578062
rect 90313 577502 90358 578062
rect 89820 577098 89890 577502
rect 90296 577098 90366 577502
rect 89626 577046 90366 577098
rect 89626 576814 90304 577046
rect 89608 576738 90304 576814
rect 89626 576713 90304 576738
rect 90313 576713 90358 577046
rect 90495 576713 90540 578062
rect 90894 577572 93129 578377
rect 94136 578513 99314 578518
rect 102856 578513 103277 578549
rect 94136 578484 103277 578513
rect 94136 578344 94170 578484
rect 94612 578454 94646 578484
rect 97654 578454 97688 578484
rect 97785 578479 103277 578484
rect 97785 578454 99314 578479
rect 94612 578416 94650 578454
rect 94910 578416 99314 578454
rect 94312 578411 99314 578416
rect 99689 578411 99723 578449
rect 101339 578427 101350 578438
rect 101362 578427 101373 578438
rect 101339 578411 101373 578427
rect 102856 578411 103277 578479
rect 94312 578382 101749 578411
rect 94612 578356 94646 578382
rect 96804 578376 96832 578382
rect 97456 578376 97484 578382
rect 96776 578356 96804 578376
rect 96832 578356 96860 578376
rect 97428 578356 97456 578376
rect 97484 578356 97512 578376
rect 97654 578356 97688 578382
rect 97785 578377 101749 578382
rect 102378 578377 102407 578411
rect 97785 578356 99314 578377
rect 94296 578344 99314 578356
rect 94102 578310 99314 578344
rect 94136 577686 94170 578310
rect 94250 577686 94284 578310
rect 94296 578298 94297 578299
rect 94295 578297 94296 578298
rect 94295 577698 94296 577699
rect 94296 577697 94297 577698
rect 94612 577686 94646 578310
rect 94726 577686 94760 578310
rect 94908 577896 94953 578310
rect 95384 577984 95429 578310
rect 95566 577984 95611 578310
rect 96042 577984 96087 578310
rect 96224 577984 96269 578310
rect 96700 577984 96745 578310
rect 96882 577984 96927 578310
rect 97358 577984 97403 578310
rect 97540 577984 97585 578310
rect 97654 577984 97688 578310
rect 97785 577984 99314 578310
rect 95056 577952 99314 577984
rect 99689 577952 99723 578377
rect 99792 578318 99848 578329
rect 99898 578318 99954 578329
rect 100450 578318 100506 578329
rect 100556 578318 100612 578329
rect 101108 578318 101164 578329
rect 101214 578318 101270 578329
rect 99803 577952 99848 578318
rect 99909 577952 99954 578318
rect 95056 577918 100182 577952
rect 95056 577897 99314 577918
rect 99689 577897 99723 577918
rect 99803 577897 99848 577918
rect 99909 577897 99954 577918
rect 94908 577686 94942 577896
rect 95056 577850 100053 577897
rect 95056 577816 99395 577850
rect 99438 577816 100053 577850
rect 95056 577686 99314 577816
rect 99365 577757 99421 577768
rect 94102 577652 99314 577686
rect 94136 577572 94170 577652
rect 94250 577572 94284 577652
rect 94612 577572 94646 577652
rect 94726 577572 94771 577652
rect 94908 577580 94953 577652
rect 95056 577580 99314 577652
rect 94816 577578 99314 577580
rect 94876 577572 99314 577578
rect 90894 577538 99314 577572
rect 90894 577502 93129 577538
rect 90971 576713 91016 577502
rect 91036 577136 91064 577140
rect 91092 577136 91120 577140
rect 91153 577136 91198 577502
rect 91629 577486 91674 577502
rect 91608 577364 91678 577486
rect 91608 577292 91704 577364
rect 91608 577136 91678 577292
rect 91036 577030 91678 577136
rect 91706 577118 91734 577140
rect 91762 577118 91790 577140
rect 91811 577118 91856 577502
rect 91706 577084 92272 577118
rect 91706 577040 91740 577084
rect 91036 576714 91674 577030
rect 91698 576990 91740 577040
rect 91762 577046 91790 577084
rect 91762 576990 91802 577046
rect 91698 576984 91746 576990
rect 91762 576989 91774 576990
rect 91811 576989 91856 577084
rect 91890 577004 92088 577015
rect 91761 576984 91858 576989
rect 91706 576864 91746 576984
rect 91754 576976 91858 576984
rect 91754 576942 91876 576976
rect 91901 576970 92088 577004
rect 92089 576942 92217 576989
rect 91754 576864 91774 576942
rect 91808 576915 91876 576942
rect 91800 576904 91876 576915
rect 92136 576904 92217 576942
rect 91698 576808 91746 576864
rect 91036 576713 91064 576714
rect 91092 576713 91120 576714
rect 91153 576713 91198 576714
rect 87293 576679 91225 576713
rect 89065 576664 89099 576679
rect 89173 576664 89219 576679
rect 89541 576664 89575 576679
rect 89626 576664 90304 576679
rect 90313 576664 90358 576679
rect 90495 576664 90540 576679
rect 90715 576664 90749 576679
rect 88646 576658 90870 576664
rect 90971 576658 91016 576679
rect 91036 576660 91064 576679
rect 91092 576660 91120 576679
rect 91153 576660 91225 576679
rect 91629 576660 91674 576714
rect 91706 576790 91746 576808
rect 91762 576790 91774 576864
rect 91706 576762 91740 576790
rect 91762 576762 91802 576790
rect 91811 576762 91856 576904
rect 91890 576876 92088 576887
rect 91901 576842 92088 576876
rect 92238 576762 92272 577084
rect 91706 576754 92272 576762
rect 92287 576754 92332 577502
rect 92414 577026 92442 577140
rect 92414 576754 92442 576840
rect 92469 576754 92514 577502
rect 92583 576754 92617 577502
rect 91706 576728 93129 576754
rect 91706 576668 91734 576728
rect 91762 576668 91790 576728
rect 91036 576658 91674 576660
rect 88646 576649 91674 576658
rect 87197 575859 87231 576617
rect 87673 576611 87707 576649
rect 88550 576630 91674 576649
rect 91811 576642 91856 576728
rect 92232 576718 93129 576728
rect 94136 576718 94170 577538
rect 94612 576718 94646 577538
rect 94726 576718 94771 577538
rect 94876 577510 99314 577538
rect 94908 577456 94953 577510
rect 95056 577502 99314 577510
rect 95056 577456 98200 577502
rect 94876 577414 98200 577456
rect 94870 577408 98200 577414
rect 94802 576718 94830 577140
rect 94908 576718 94953 577408
rect 95056 577046 98200 577408
rect 95384 576718 95429 577046
rect 95454 576718 95482 577046
rect 95510 576718 95538 577046
rect 95566 576718 95611 577046
rect 96042 576718 96087 577046
rect 96112 576718 96140 577046
rect 96168 576718 96196 577046
rect 96224 576718 96269 577046
rect 92232 576684 96296 576718
rect 92232 576642 93129 576684
rect 88550 576611 88584 576630
rect 89065 576611 89099 576630
rect 89167 576611 91674 576630
rect 87673 576600 91674 576611
rect 91706 576616 93129 576642
rect 93586 576622 93614 576654
rect 93642 576622 93670 576654
rect 94136 576616 94170 576684
rect 94244 576654 94290 576684
rect 94612 576654 94646 576684
rect 94726 576654 94771 576684
rect 94802 576654 94830 576684
rect 94908 576654 94953 576684
rect 95384 576654 95429 576684
rect 95454 576654 95482 576684
rect 95510 576654 95538 576684
rect 95566 576654 95611 576684
rect 95786 576654 95820 576684
rect 96042 576654 96087 576684
rect 96112 576654 96140 576684
rect 94238 576616 96158 576654
rect 91706 576608 96158 576616
rect 87361 576571 87428 576584
rect 87673 576577 91663 576600
rect 83569 575825 87501 575859
rect 83473 574059 83507 575763
rect 83949 575757 83983 575795
rect 86991 575773 87002 575784
rect 87014 575773 87025 575784
rect 86991 575757 87025 575773
rect 87197 575757 87231 575825
rect 87311 575791 87358 575804
rect 87311 575788 87359 575791
rect 87299 575757 87359 575788
rect 83649 575723 87359 575757
rect 83949 574059 83983 575723
rect 84052 575664 84108 575675
rect 84234 575664 84290 575675
rect 84710 575664 84766 575675
rect 84892 575664 84948 575675
rect 85368 575664 85413 575675
rect 85550 575664 85595 575675
rect 86026 575664 86071 575675
rect 86208 575664 86253 575675
rect 86684 575664 86729 575675
rect 86866 575664 86911 575675
rect 84063 575408 84784 575664
rect 84063 574059 84108 575408
rect 84124 574059 84152 575340
rect 84245 574059 84290 575408
rect 84721 574059 84766 575408
rect 84782 574059 84810 575340
rect 84838 574059 84866 575340
rect 84903 574059 84948 575664
rect 81701 574025 85157 574059
rect 83473 567527 83507 574025
rect 83949 574004 83983 574025
rect 84063 574022 84108 574025
rect 84063 574004 84097 574022
rect 83587 573988 83634 574004
rect 83575 573957 83634 573988
rect 83665 573963 83712 574004
rect 83648 573957 83712 573963
rect 83949 573957 83996 574004
rect 84063 573957 84110 574004
rect 84124 573976 84152 574025
rect 84245 574022 84290 574025
rect 84721 574022 84766 574025
rect 84245 574004 84279 574022
rect 84721 574004 84755 574022
rect 84245 573957 84292 574004
rect 84323 573957 84370 574004
rect 84721 573957 84768 574004
rect 84782 573976 84810 574025
rect 84838 573976 84866 574025
rect 84903 574022 84948 574025
rect 84903 574004 84937 574022
rect 84903 573957 84950 574004
rect 84981 573957 85028 574004
rect 83575 573923 83712 573957
rect 83755 573923 84370 573957
rect 84413 573923 85028 573957
rect 83575 573917 83677 573923
rect 83575 573876 83633 573917
rect 83704 573889 83705 573923
rect 83587 573632 83621 573876
rect 83682 573864 83727 573875
rect 83587 572168 83627 573632
rect 83644 572224 83655 573576
rect 83587 567688 83621 572168
rect 83631 568012 83662 569414
rect 83687 567984 83690 569442
rect 83693 567676 83727 573864
rect 83949 567676 83983 573923
rect 84063 567688 84097 573923
rect 84245 567688 84279 573923
rect 84340 573864 84385 573875
rect 84351 571866 84385 573864
rect 84282 571858 84494 571866
rect 84282 571418 84694 571858
rect 84351 567676 84385 571418
rect 84482 571410 84694 571418
rect 84721 567688 84755 573923
rect 84903 567688 84937 573923
rect 84998 573864 85043 573875
rect 85009 571858 85043 573864
rect 85123 571866 85157 574025
rect 85345 574022 85360 575128
rect 85123 571858 85340 571866
rect 84958 571418 85340 571858
rect 84958 571410 85170 571418
rect 85009 567676 85043 571410
rect 83681 567629 83740 567676
rect 83949 567629 83996 567676
rect 84339 567629 84398 567676
rect 84997 567629 85055 567676
rect 83649 567595 85055 567629
rect 83581 567533 83604 567589
rect 83681 567579 83739 567595
rect 83693 567527 83727 567561
rect 83949 567527 83983 567595
rect 84286 567582 84397 567595
rect 84339 567580 84397 567582
rect 84314 567579 84397 567580
rect 84997 567579 85055 567595
rect 84314 567527 84345 567579
rect 85040 567564 85055 567579
rect 85123 567629 85157 571410
rect 85379 567688 85413 575664
rect 85444 569990 85472 575340
rect 85500 569990 85528 575340
rect 85444 567635 85472 569804
rect 85500 567635 85528 569804
rect 85561 567688 85595 575664
rect 85812 571858 85816 571866
rect 85824 571418 85828 571858
rect 86037 570724 86071 575664
rect 86037 570534 86082 570724
rect 86114 570534 86142 575340
rect 86170 570534 86198 575340
rect 86219 570724 86253 575664
rect 86695 574100 86729 575664
rect 86822 574100 86850 575340
rect 86877 574100 86911 575664
rect 86991 574100 87025 575723
rect 87197 574100 87231 575723
rect 87299 575714 87341 575723
rect 87299 575676 87345 575714
rect 87311 574100 87345 575676
rect 87353 575675 87379 575680
rect 87353 574100 87387 575675
rect 87467 574100 87501 575825
rect 87673 574100 87707 576577
rect 87876 576571 87904 576577
rect 88534 576571 88584 576577
rect 87776 576518 87821 576529
rect 87848 576528 87876 576571
rect 87958 576518 88003 576529
rect 88434 576518 88479 576529
rect 88506 576528 88534 576571
rect 88550 576528 88590 576571
rect 89065 576562 89099 576577
rect 89167 576562 89226 576577
rect 89541 576562 89575 576577
rect 89643 576562 89702 576577
rect 89837 576562 89884 576577
rect 90301 576562 90360 576577
rect 90495 576562 90542 576577
rect 90694 576562 90749 576577
rect 88710 576543 90749 576562
rect 88726 576539 90749 576543
rect 89065 576530 90749 576539
rect 87787 575874 87821 576518
rect 87969 575874 88003 576518
rect 88445 575874 88479 576518
rect 88550 575900 88584 576528
rect 88616 576518 88661 576529
rect 88726 576528 90749 576530
rect 88627 576480 88661 576518
rect 88664 576480 88695 576485
rect 89065 576481 89149 576528
rect 88627 576469 88698 576480
rect 88627 575900 88661 576469
rect 88664 575900 88698 576469
rect 89065 575900 89099 576481
rect 89103 575984 89137 576481
rect 89179 575984 89213 576528
rect 89274 576518 89319 576528
rect 89285 575984 89319 576518
rect 89103 575900 89148 575984
rect 89179 575900 89224 575984
rect 89285 575900 89330 575984
rect 89541 575900 89575 576528
rect 89655 575984 89689 576528
rect 89749 576481 89807 576528
rect 89761 575984 89795 576481
rect 89837 575984 89871 576528
rect 89932 576518 89977 576528
rect 89943 575984 89977 576518
rect 90313 575984 90347 576528
rect 90407 576481 90465 576528
rect 90419 575984 90453 576481
rect 90495 575984 90529 576528
rect 90590 576518 90635 576528
rect 90601 575984 90635 576518
rect 90715 576480 90749 576528
rect 90715 575984 90756 576480
rect 89655 575900 89700 575984
rect 89761 575900 89806 575984
rect 89837 575900 89882 575984
rect 89943 575900 89988 575984
rect 90313 575900 90358 575984
rect 90419 575900 90464 575984
rect 90495 575900 90540 575984
rect 90601 575900 90646 575984
rect 90715 575900 90767 575984
rect 90836 575900 90870 576577
rect 90894 576270 90904 576577
rect 90959 576530 91663 576577
rect 90971 576528 91663 576530
rect 90971 576270 91016 576528
rect 90971 575984 91005 576270
rect 91036 576238 91663 576528
rect 91706 576584 91740 576608
rect 91811 576600 91856 576608
rect 91706 576570 91762 576584
rect 91706 576528 91740 576570
rect 91762 576528 91790 576570
rect 91706 576514 91762 576528
rect 91706 576286 91740 576514
rect 91811 576513 91845 576600
rect 92232 576582 96158 576608
rect 92077 576528 92088 576539
rect 91761 576500 91858 576513
rect 91761 576466 91876 576500
rect 91901 576494 92088 576528
rect 92089 576466 92170 576513
rect 91808 576439 91876 576466
rect 91800 576428 91876 576439
rect 92136 576428 92170 576466
rect 91811 576286 91845 576428
rect 92077 576400 92088 576411
rect 91901 576366 92088 576400
rect 92232 576286 93129 576582
rect 93614 576576 93642 576582
rect 93505 576532 93561 576543
rect 91706 576252 93129 576286
rect 91077 575984 91111 576238
rect 91153 575984 91187 576238
rect 91191 575984 91225 576238
rect 90971 575900 91016 575984
rect 91077 575900 91122 575984
rect 91153 575900 91225 575984
rect 91629 575984 91663 576238
rect 91811 575984 91845 576252
rect 91629 575900 91674 575984
rect 91811 575900 91856 575984
rect 92232 575900 93129 576252
rect 88508 575895 93129 575900
rect 93516 575895 93561 576532
rect 93586 576528 93614 576576
rect 93642 576528 93670 576576
rect 94136 576543 94170 576582
rect 94238 576576 94300 576582
rect 94238 576544 94296 576576
rect 93687 576532 93743 576543
rect 93698 575895 93743 576532
rect 94136 576532 94219 576543
rect 94136 576276 94170 576532
rect 94174 576276 94219 576532
rect 94244 576528 94295 576544
rect 94300 576543 94346 576576
rect 94300 576532 94401 576543
rect 94300 576528 94346 576532
rect 94250 576276 94295 576528
rect 94356 576276 94401 576532
rect 94612 576276 94646 576582
rect 94714 576544 94772 576582
rect 94726 576276 94771 576544
rect 94821 576532 94877 576543
rect 94832 576276 94877 576532
rect 94908 576276 94953 576582
rect 95372 576544 95430 576582
rect 95003 576532 95059 576543
rect 95014 576276 95059 576532
rect 95384 576276 95429 576544
rect 95479 576532 95535 576543
rect 95490 576276 95535 576532
rect 95566 576276 95611 576582
rect 95661 576532 95717 576543
rect 95672 576276 95717 576532
rect 95786 576276 95820 576582
rect 96030 576544 96140 576582
rect 96168 576544 96196 576684
rect 96042 576543 96140 576544
rect 96142 576543 96196 576544
rect 96042 576532 96196 576543
rect 96042 576528 96140 576532
rect 96142 576528 96196 576532
rect 96042 576276 96087 576528
rect 96148 576276 96193 576528
rect 96224 576276 96296 576684
rect 96700 576282 96745 577046
rect 96776 576528 96804 577046
rect 96832 576528 96860 577046
rect 96882 576282 96927 577046
rect 97358 576282 97403 577046
rect 97428 576592 97456 577046
rect 97484 576528 97512 577046
rect 97540 576282 97585 577046
rect 97654 576282 97688 577046
rect 97785 576713 98200 577046
rect 98550 576713 98556 577140
rect 98604 576747 98638 577502
rect 98654 577012 98678 577140
rect 98718 576781 98763 577502
rect 98593 576716 98638 576747
rect 98654 576716 98678 576772
rect 99251 576769 99296 577502
rect 99376 576781 99421 577757
rect 99689 576769 99723 577816
rect 99803 576814 99848 577816
rect 99909 576814 99954 577816
rect 100023 577757 100079 577768
rect 99760 576769 99954 576814
rect 100034 576781 100079 577757
rect 98733 576722 100053 576769
rect 98593 576713 98678 576716
rect 98780 576713 99395 576722
rect 99438 576713 100053 576722
rect 100148 576713 100182 577918
rect 100461 577140 100506 578318
rect 100567 577140 100612 578318
rect 101119 577950 101164 578318
rect 101225 577950 101270 578318
rect 101339 577950 101373 578377
rect 102416 578339 102445 578406
rect 102497 578377 103277 578411
rect 100461 576713 100546 577140
rect 100561 576713 100612 577140
rect 100690 577916 102268 577950
rect 100690 576713 100724 577916
rect 101119 577895 101164 577916
rect 101225 577895 101270 577916
rect 101339 577895 101373 577916
rect 100819 577848 101481 577895
rect 101777 577864 101824 577895
rect 101765 577848 101824 577864
rect 102092 577848 102139 577895
rect 100866 577814 101481 577848
rect 101524 577816 102139 577848
rect 101518 577814 102139 577816
rect 100793 577755 100849 577766
rect 100804 576779 100849 577755
rect 101119 577416 101164 577814
rect 101225 577464 101270 577814
rect 101210 577416 101280 577464
rect 101028 577262 101280 577416
rect 101119 576767 101164 577262
rect 101210 577008 101280 577262
rect 101225 576767 101270 577008
rect 101339 576767 101373 577814
rect 101518 577780 101576 577782
rect 101765 577767 101823 577814
rect 101451 577755 101507 577766
rect 101462 576779 101507 577755
rect 101777 577604 101811 577767
rect 102109 577755 102154 577766
rect 102120 577604 102154 577755
rect 101777 577486 101822 577604
rect 101756 577412 101826 577486
rect 101676 577266 101926 577412
rect 101756 577030 101826 577266
rect 101777 576767 101822 577030
rect 102120 576779 102165 577604
rect 100819 576720 102139 576767
rect 100866 576713 101481 576720
rect 97785 576686 101481 576713
rect 101524 576686 102139 576720
rect 97785 576679 101373 576686
rect 97785 576658 98200 576679
rect 98550 576672 98556 576679
rect 98593 576658 98638 576679
rect 99239 576672 99297 576679
rect 99251 576664 99285 576672
rect 99372 576664 99416 576679
rect 99689 576664 99723 576679
rect 99803 576664 99848 576679
rect 99860 576678 99871 576679
rect 99909 576664 99954 576679
rect 100148 576664 100182 576679
rect 100461 576672 100546 576679
rect 100461 576664 100506 576672
rect 100561 576664 100612 576679
rect 100690 576664 100724 576679
rect 98698 576658 101018 576664
rect 97785 576630 101018 576658
rect 97785 576620 98732 576630
rect 99245 576620 99263 576630
rect 99273 576620 99291 576630
rect 99372 576626 99416 576630
rect 99689 576620 99723 576630
rect 99803 576627 99848 576630
rect 99791 576620 99849 576627
rect 99903 576620 99954 576630
rect 100086 576620 100786 576630
rect 97785 576618 100786 576620
rect 100984 576618 101018 576630
rect 101119 576627 101164 576679
rect 101182 576648 101187 576679
rect 101225 576645 101270 576679
rect 101107 576618 101165 576627
rect 101219 576618 101270 576645
rect 101339 576618 101373 576679
rect 101765 576670 101823 576686
rect 102234 576618 102268 577916
rect 97785 576611 102268 576618
rect 97785 576609 100612 576611
rect 97785 576600 100614 576609
rect 100629 576600 102268 576611
rect 97785 576586 102268 576600
rect 97785 576577 98633 576586
rect 98639 576584 102268 576586
rect 98639 576577 101270 576584
rect 97785 576282 98200 576577
rect 98500 576571 98577 576577
rect 98587 576543 98633 576577
rect 98643 576571 98732 576577
rect 94034 575895 96342 576276
rect 96612 576246 98200 576282
rect 98593 576246 98627 576543
rect 98698 576246 98732 576571
rect 99239 576562 99298 576577
rect 99689 576562 99723 576577
rect 99791 576562 99850 576577
rect 99909 576562 99956 576577
rect 100449 576562 100508 576577
rect 100567 576562 100614 576577
rect 100842 576562 100889 576577
rect 98858 576543 100889 576562
rect 98874 576528 100889 576543
rect 99239 576481 99297 576528
rect 98801 576469 98846 576480
rect 98812 576326 98846 576469
rect 98812 576246 98857 576326
rect 96612 576212 98884 576246
rect 96612 576144 98200 576212
rect 98698 576191 98732 576212
rect 98593 576160 98640 576191
rect 98581 576144 98640 576160
rect 98698 576144 98745 576191
rect 96612 576110 98745 576144
rect 96612 575900 98200 576110
rect 98581 576063 98639 576110
rect 98593 575984 98627 576063
rect 98698 576062 98732 576110
rect 98736 576062 98766 576067
rect 98698 576051 98770 576062
rect 98593 575900 98638 575984
rect 98698 575900 98732 576051
rect 98736 575984 98770 576051
rect 98736 575900 98781 575984
rect 98812 575900 98884 576212
rect 99251 575984 99285 576481
rect 99251 575900 99296 575984
rect 99689 575900 99723 576528
rect 99803 575984 99837 576528
rect 99897 576481 99955 576528
rect 99909 575984 99943 576481
rect 99803 575900 99848 575984
rect 99909 575900 99954 575984
rect 100461 575900 100495 576528
rect 100555 576481 100613 576528
rect 100567 575900 100601 576481
rect 100859 576469 100904 576480
rect 100870 575900 100904 576469
rect 100984 575900 101018 576577
rect 101107 576530 101165 576577
rect 101191 576571 101209 576577
rect 101219 576543 101270 576577
rect 101119 576338 101164 576530
rect 101225 576338 101270 576543
rect 101339 576338 101373 576584
rect 101777 576338 101811 576372
rect 102435 576338 102469 578318
rect 102856 577988 103277 578377
rect 103516 578518 105954 578554
rect 106182 578518 106216 590322
rect 106296 587764 106330 590232
rect 106284 587730 106800 587764
rect 106296 587700 106330 587730
rect 106754 587700 106788 587730
rect 106296 587662 106680 587700
rect 106726 587662 106788 587700
rect 106806 587692 106822 587730
rect 106296 580104 106330 587662
rect 106358 587628 106788 587662
rect 106754 580244 106788 587628
rect 106726 580206 106788 580244
rect 106342 580172 106788 580206
rect 106754 580104 106788 580172
rect 106810 580104 106822 580144
rect 106278 580070 106800 580104
rect 106806 580070 106822 580104
rect 106776 579982 106788 580070
rect 106810 580016 106822 580070
rect 106868 578518 106902 590322
rect 112093 585450 112127 590389
rect 112985 588934 113019 590451
rect 113040 590371 113168 590383
rect 119642 590382 119676 590451
rect 116120 590371 119676 590382
rect 119756 590371 119790 590451
rect 120264 590371 120275 590382
rect 113040 590337 120275 590371
rect 113071 590325 113168 590337
rect 113025 590296 113081 590310
rect 113068 590280 113081 590296
rect 113040 590252 113081 590254
rect 113087 590221 113121 590325
rect 119642 590310 119676 590337
rect 113127 590280 119750 590310
rect 119642 590254 119676 590280
rect 113127 590252 119750 590254
rect 119642 590204 119676 590252
rect 116120 590193 119676 590204
rect 119756 590193 119790 590337
rect 119796 590280 120092 590310
rect 120276 590309 120357 590356
rect 119796 590252 120092 590254
rect 120036 590224 120092 590252
rect 120323 590206 120357 590309
rect 120276 590193 120357 590206
rect 120425 590204 120459 590451
rect 121215 590221 121296 590490
rect 120422 590193 121167 590204
rect 113040 590131 113121 590178
rect 113180 590159 121167 590193
rect 113087 589726 113121 590131
rect 113040 589725 113121 589726
rect 113040 589713 113168 589725
rect 119642 589724 119676 590159
rect 116120 589713 119676 589724
rect 119756 589713 119790 590159
rect 120323 589741 120357 590159
rect 120264 589713 120275 589724
rect 113040 589679 120275 589713
rect 113071 589667 113168 589679
rect 113087 589563 113121 589667
rect 119642 589652 119676 589679
rect 113127 589618 119750 589652
rect 119642 589596 119676 589618
rect 113127 589562 119750 589596
rect 119642 589546 119676 589562
rect 116120 589535 119676 589546
rect 119756 589535 119790 589679
rect 119796 589618 120092 589652
rect 120276 589651 120357 589698
rect 119796 589562 120092 589596
rect 120323 589548 120357 589651
rect 120276 589535 120357 589548
rect 120425 589546 120459 590159
rect 121168 590131 121296 590178
rect 121215 589563 121296 590131
rect 120422 589535 121167 589546
rect 113040 589473 113121 589520
rect 113180 589501 121167 589535
rect 113087 589068 113121 589473
rect 113040 589067 113121 589068
rect 113040 589055 113168 589067
rect 119642 589066 119676 589501
rect 116120 589055 119676 589066
rect 119756 589055 119790 589501
rect 120323 589083 120357 589501
rect 120264 589055 120275 589066
rect 113040 589021 120275 589055
rect 113071 589009 113168 589021
rect 113068 588960 113081 588962
rect 112985 588904 113081 588934
rect 113087 588905 113121 589009
rect 119642 588962 119676 589021
rect 113127 588960 119750 588962
rect 119642 588934 119676 588960
rect 113127 588904 119750 588934
rect 112985 588763 113019 588904
rect 119642 588888 119676 588904
rect 116120 588877 119676 588888
rect 119756 588877 119790 589021
rect 120276 588993 120357 589040
rect 120036 588962 120092 588990
rect 119796 588960 120092 588962
rect 119796 588904 120092 588934
rect 120323 588890 120357 588993
rect 120276 588877 120357 588890
rect 120425 588888 120459 589501
rect 121168 589473 121296 589520
rect 121215 588905 121296 589473
rect 120422 588877 121167 588888
rect 113180 588843 121167 588877
rect 119642 588763 119676 588843
rect 119756 588763 119790 588843
rect 120323 588763 120357 588843
rect 120425 588763 120459 588843
rect 121317 588763 121351 591383
rect 122816 591076 122848 591498
rect 122854 591114 122886 591460
rect 124855 591043 124889 591848
rect 124957 591843 124991 591848
rect 125578 591842 125592 591848
rect 125792 591842 125856 591848
rect 124957 591827 124991 591836
rect 125564 591834 125578 591842
rect 125592 591834 125634 591842
rect 125094 591827 125714 591834
rect 125860 591827 126234 591848
rect 128646 591842 128914 591848
rect 125038 591821 128918 591827
rect 125038 591815 128942 591821
rect 129044 591815 129078 591873
rect 131680 591815 131714 591873
rect 131735 591850 131816 591873
rect 131863 591872 133221 591873
rect 134446 591872 134502 591876
rect 135690 591872 135746 591876
rect 133038 591866 133135 591872
rect 131782 591834 131816 591850
rect 131835 591844 132732 591866
rect 131754 591815 132210 591834
rect 133079 591831 133125 591866
rect 133085 591827 133119 591831
rect 133026 591815 133037 591826
rect 125034 591814 133037 591815
rect 124952 591800 125025 591802
rect 125038 591801 133037 591814
rect 133051 591803 133153 591820
rect 124910 591753 125038 591800
rect 125050 591759 133037 591801
rect 124957 591163 125038 591753
rect 125094 591412 125714 591759
rect 125764 591464 125798 591759
rect 125872 591691 125906 591759
rect 126135 591706 126146 591717
rect 125819 591678 125919 591691
rect 125819 591644 125934 591678
rect 125959 591672 126146 591706
rect 126147 591644 126228 591691
rect 125860 591606 125934 591644
rect 126194 591606 126228 591644
rect 125860 591590 125918 591606
rect 125872 591464 125906 591590
rect 126135 591578 126146 591589
rect 125959 591544 126146 591578
rect 126296 591464 126330 591759
rect 128930 591564 128964 591759
rect 129044 591564 129078 591759
rect 125764 591430 126330 591464
rect 128772 591554 129220 591564
rect 125094 591168 125714 591358
rect 125872 591344 125906 591430
rect 128772 591352 129228 591554
rect 125764 591310 126330 591344
rect 128780 591342 129228 591352
rect 125764 591236 125798 591310
rect 125764 591228 125866 591236
rect 125872 591228 125906 591310
rect 126135 591230 126146 591241
rect 125764 591198 125804 591228
rect 125872 591215 125912 591228
rect 125819 591208 125919 591215
rect 125812 591202 125919 591208
rect 125812 591198 125934 591202
rect 125754 591184 125762 591190
rect 125012 591157 125029 591163
rect 125039 591157 125714 591168
rect 125764 591178 125798 591198
rect 125819 591178 125934 591198
rect 125959 591196 126146 591230
rect 126147 591178 126228 591215
rect 126296 591178 126330 591310
rect 125764 591168 126420 591178
rect 125764 591157 126520 591168
rect 128930 591157 128964 591342
rect 129044 591157 129078 591342
rect 131680 591157 131714 591759
rect 131716 591744 132172 591759
rect 133038 591753 133119 591800
rect 131782 591282 131816 591744
rect 133085 591266 133119 591753
rect 133038 591254 133135 591266
rect 133187 591254 133221 591872
rect 134446 591816 134502 591820
rect 135690 591816 135746 591820
rect 134446 591314 134502 591316
rect 135690 591314 135746 591316
rect 134446 591258 134502 591260
rect 135690 591258 135746 591260
rect 131735 591232 131816 591239
rect 131735 591228 131850 591232
rect 131735 591204 131816 591228
rect 131875 591220 135136 591254
rect 133038 591219 133135 591220
rect 131863 591214 133135 591219
rect 132692 591208 133135 591214
rect 131735 591192 131822 591204
rect 132692 591202 133119 591208
rect 131776 591172 131822 591192
rect 131782 591169 131822 591172
rect 131766 591163 131863 591169
rect 131766 591158 132692 591163
rect 131766 591157 131863 591158
rect 133026 591157 133037 591168
rect 125012 591120 133037 591157
rect 133079 591163 133119 591202
rect 133079 591156 133094 591163
rect 124910 591073 125038 591120
rect 125050 591101 133037 591120
rect 124957 591056 125038 591073
rect 124910 591043 125038 591056
rect 125094 591043 125714 591101
rect 125746 591080 126400 591101
rect 128917 591089 128918 591090
rect 128918 591088 128919 591089
rect 125764 591043 125798 591080
rect 125872 591064 125906 591080
rect 125959 591077 126146 591080
rect 125943 591068 126151 591077
rect 125872 591046 125912 591064
rect 126170 591052 126226 591080
rect 126142 591046 126226 591052
rect 125872 591043 125906 591046
rect 126296 591043 126330 591080
rect 128930 591043 128964 591101
rect 129044 591043 129078 591101
rect 131680 591043 131714 591101
rect 131766 591089 131863 591101
rect 131782 591043 131816 591089
rect 133038 591073 133119 591120
rect 133085 591056 133119 591073
rect 133038 591043 133119 591056
rect 133187 591043 133221 591220
rect 124855 591009 133221 591043
rect 112985 588729 121351 588763
rect 119642 588510 119676 588729
rect 112182 588486 112189 588510
rect 112235 588486 119750 588510
rect 119642 588397 119676 588486
rect 119756 588397 119790 588729
rect 119796 588486 120092 588510
rect 120036 588430 120092 588454
rect 120323 588425 120357 588729
rect 119801 588409 119802 588410
rect 119802 588408 119803 588409
rect 120264 588397 120275 588408
rect 119608 588363 120275 588397
rect 119642 587831 119676 588363
rect 119756 587831 119790 588363
rect 119802 588351 119803 588352
rect 119801 588350 119802 588351
rect 120276 588335 120357 588382
rect 120323 587831 120357 588335
rect 120425 587831 120459 588729
rect 122816 588422 122848 588844
rect 122854 588460 122886 588806
rect 124855 588389 124889 591009
rect 124957 590588 125038 591009
rect 125094 590936 125714 591009
rect 125764 590988 125798 591009
rect 125872 590988 125906 591009
rect 125912 591008 125946 591009
rect 126142 590990 126226 591009
rect 126296 590988 126330 591009
rect 125764 590954 126330 590988
rect 124957 590570 124991 590588
rect 125872 590570 125906 590954
rect 128930 590918 128964 591009
rect 129044 590918 129078 591009
rect 128772 590706 129220 590918
rect 128804 590570 129080 590706
rect 131680 590578 131714 591009
rect 131782 590624 131816 591009
rect 133085 590609 133119 591009
rect 133038 590608 133119 590609
rect 133038 590596 133135 590608
rect 131875 590578 133135 590596
rect 131410 590576 131776 590578
rect 131822 590576 133135 590578
rect 131680 590570 131714 590576
rect 131863 590570 133135 590576
rect 133187 590570 133221 591009
rect 134446 590650 134502 590658
rect 135690 590650 135746 590658
rect 134446 590594 134502 590602
rect 135690 590594 135746 590602
rect 124952 590462 133372 590570
rect 134446 590556 134502 590564
rect 135690 590556 135856 590584
rect 134446 590500 134502 590508
rect 135690 590500 135746 590528
rect 124910 590415 133372 590462
rect 124952 589804 133372 590415
rect 124910 589757 133372 589804
rect 124952 589754 133372 589757
rect 124952 589146 133257 589754
rect 124910 589099 133257 589146
rect 124952 588389 133257 589099
rect 124855 588355 133257 588389
rect 112168 587820 120459 587831
rect 112179 587808 120459 587820
rect 112168 587797 120459 587808
rect 112195 587751 112229 587797
rect 112578 587760 113980 587776
rect 112984 587739 113638 587760
rect 119642 587739 119676 587797
rect 119756 587739 119790 587797
rect 119801 587751 119802 587752
rect 120323 587751 120357 587797
rect 119802 587750 119803 587751
rect 120264 587739 120275 587750
rect 112288 587683 120275 587739
rect 112195 587087 112229 587677
rect 113004 587662 113658 587683
rect 116018 587488 116466 587498
rect 116010 587286 116466 587488
rect 116010 587276 116458 587286
rect 119034 587096 119440 587474
rect 118954 587092 119440 587096
rect 119642 587092 119676 587683
rect 116120 587081 119676 587092
rect 119756 587081 119790 587683
rect 120276 587677 120357 587724
rect 120264 587081 120275 587092
rect 120323 587087 120357 587677
rect 112288 587025 120275 587081
rect 118992 587006 119448 587025
rect 112195 586997 112229 587001
rect 119034 586967 119440 587006
rect 119642 586967 119676 587025
rect 119756 586967 119790 587025
rect 119802 587013 119803 587014
rect 119801 587012 119802 587013
rect 120276 586997 120357 587044
rect 120323 586980 120357 586997
rect 120276 586967 120357 586980
rect 120425 586967 120459 587797
rect 112157 586933 120459 586967
rect 116234 586822 116366 586832
rect 116010 586610 116458 586822
rect 119642 586401 119676 586933
rect 119756 586401 119790 586933
rect 120323 586429 120357 586933
rect 119801 586413 119802 586414
rect 119802 586412 119803 586413
rect 120264 586401 120275 586412
rect 119608 586367 120275 586401
rect 114702 586264 115012 586270
rect 115698 586176 116318 586270
rect 116368 586222 116934 586256
rect 116368 586176 116402 586222
rect 115698 586127 116466 586176
rect 116552 586142 116750 586153
rect 115698 586042 116551 586127
rect 116563 586108 116750 586142
rect 116751 586080 116879 586127
rect 116798 586042 116879 586080
rect 115698 586016 116494 586042
rect 115698 585964 116466 586016
rect 116552 586014 116750 586025
rect 116563 585980 116750 586014
rect 115698 585848 116318 585964
rect 116368 585900 116402 585964
rect 116900 585900 116934 586222
rect 116368 585866 116934 585900
rect 119642 585848 119676 586367
rect 119756 585848 119790 586367
rect 119802 586355 119803 586356
rect 119801 586354 119802 586355
rect 120276 586339 120357 586386
rect 118568 585832 120032 585848
rect 112276 585703 115556 585720
rect 117124 585703 118624 585722
rect 119642 585652 119676 585832
rect 119750 585801 119796 585832
rect 120276 585801 120277 585802
rect 120323 585801 120357 586339
rect 120275 585800 120276 585801
rect 119722 585777 119824 585792
rect 119722 585773 120298 585777
rect 119818 585755 120298 585773
rect 120323 585755 120357 585792
rect 119802 585754 120298 585755
rect 119802 585739 120276 585754
rect 120285 585739 120395 585754
rect 119802 585722 120415 585739
rect 120425 585722 120459 586933
rect 124952 588319 133257 588355
rect 124952 587880 129114 588319
rect 124952 587869 133261 587880
rect 124952 587857 133250 587869
rect 124952 587846 133261 587857
rect 124952 587788 129114 587846
rect 131762 587800 132220 587820
rect 133200 587800 133234 587846
rect 131722 587788 132220 587800
rect 124952 587742 133150 587788
rect 124952 587732 133161 587742
rect 124952 587552 129114 587732
rect 131722 587728 132220 587732
rect 131722 587708 132180 587728
rect 131466 587684 132570 587704
rect 131438 587656 132598 587676
rect 124952 587340 129310 587552
rect 124952 587312 129292 587340
rect 124952 587130 129114 587312
rect 133150 587130 133161 587141
rect 133200 587136 133234 587726
rect 124952 587120 133161 587130
rect 124952 587074 133150 587120
rect 124952 587016 129114 587074
rect 133200 587046 133234 587050
rect 124952 586982 133268 587016
rect 124952 586880 129114 586982
rect 124952 586668 129304 586880
rect 124952 586512 129114 586668
rect 124952 586478 129154 586512
rect 124952 586450 129114 586478
rect 129120 586450 129154 586478
rect 124952 586444 129154 586450
rect 124952 586412 129114 586444
rect 129120 586412 129154 586444
rect 124952 586410 129154 586412
rect 124952 586196 129114 586410
rect 129120 586196 129154 586410
rect 124952 586162 129154 586196
rect 124952 585753 129114 586162
rect 129204 586104 129842 586566
rect 119802 585712 120459 585722
rect 121684 585712 121740 585722
rect 119802 585704 120415 585712
rect 119976 585703 120276 585704
rect 120261 585697 120276 585703
rect 120323 585693 120357 585697
rect 120317 585666 120363 585693
rect 120425 585666 120459 585712
rect 124675 585682 129114 585753
rect 120276 585656 121740 585666
rect 120425 585652 120459 585656
rect 124675 585652 129238 585682
rect 119642 585618 129238 585652
rect 120425 585450 120459 585618
rect 124675 585582 129238 585618
rect 129106 585564 129238 585582
rect 128858 585499 129306 585564
rect 133302 585499 133336 589754
rect 112080 584243 120495 585450
rect 124952 584292 133367 585499
rect 112116 581752 112150 584243
rect 115986 584178 116434 584243
rect 116234 584060 116366 584178
rect 112592 584012 113994 584026
rect 118892 583988 120312 584018
rect 120328 583996 120362 584035
rect 120430 583988 120464 584243
rect 125148 584024 128428 584039
rect 129996 584024 131496 584039
rect 132848 584024 133148 584039
rect 124929 583988 133367 584024
rect 118796 583954 133367 583988
rect 114642 583640 115036 583676
rect 114702 583580 115012 583616
rect 115734 583546 116282 583580
rect 115734 583264 115768 583546
rect 116096 583466 116107 583477
rect 115798 583422 115870 583460
rect 115920 583432 116107 583466
rect 116108 583422 116180 583460
rect 115836 583388 115870 583422
rect 115880 583410 116136 583412
rect 116096 583384 116107 583389
rect 116146 583388 116180 583422
rect 115908 583382 116108 583384
rect 116096 583378 116107 583382
rect 115920 583360 116107 583378
rect 115904 583344 116112 583360
rect 116142 583358 116232 583360
rect 115908 583338 115910 583344
rect 116104 583338 116108 583344
rect 116248 583332 116282 583546
rect 115880 583326 115910 583332
rect 116104 583330 116282 583332
rect 116104 583326 116136 583330
rect 115870 583310 116146 583326
rect 115882 583306 116134 583310
rect 116248 583298 116282 583330
rect 115774 583292 116282 583298
rect 116248 583264 116282 583292
rect 115734 583230 116282 583264
rect 116332 583176 116970 583638
rect 118796 583326 118830 583954
rect 120328 583926 120362 583938
rect 119640 583886 119678 583924
rect 120294 583892 120314 583898
rect 120322 583892 120362 583926
rect 120328 583886 120362 583892
rect 118972 583852 119678 583886
rect 119730 583852 120414 583886
rect 120289 583814 120290 583815
rect 120290 583813 120291 583814
rect 118899 583802 118944 583813
rect 119657 583802 119702 583813
rect 118910 583326 118944 583802
rect 118955 583338 118956 583339
rect 119656 583338 119657 583339
rect 118956 583337 118957 583338
rect 119655 583337 119656 583338
rect 119668 583326 119702 583802
rect 120328 583410 120362 583852
rect 120392 583410 120400 583842
rect 119713 583338 119714 583339
rect 119714 583337 119715 583338
rect 120278 583326 120289 583337
rect 118762 583292 120289 583326
rect 120294 583314 120314 583410
rect 120322 583354 120362 583410
rect 120420 583382 120428 583814
rect 120322 583342 120342 583354
rect 120294 583302 120314 583304
rect 115984 582862 116432 583074
rect 118796 582760 118830 583292
rect 118910 582760 118944 583292
rect 118956 583280 118957 583281
rect 119655 583280 119656 583281
rect 118955 583279 118956 583280
rect 119656 583279 119657 583280
rect 119668 582760 119702 583292
rect 119714 583280 119715 583281
rect 119713 583279 119714 583280
rect 120290 583264 120362 583302
rect 120294 583194 120314 583264
rect 120322 583194 120362 583264
rect 120328 582760 120362 583194
rect 120430 582760 120464 583954
rect 120472 583852 120511 583886
rect 112191 582749 120464 582760
rect 112202 582737 120464 582749
rect 112191 582726 120464 582737
rect 112218 582680 112252 582726
rect 112984 582668 113638 582686
rect 118796 582668 118830 582726
rect 118910 582668 118944 582726
rect 118955 582680 118956 582681
rect 119656 582680 119657 582681
rect 118956 582679 118957 582680
rect 119655 582679 119656 582680
rect 119668 582668 119702 582726
rect 119713 582680 119714 582681
rect 119714 582679 119715 582680
rect 120278 582668 120289 582679
rect 112302 582612 120289 582668
rect 120294 582656 120314 582726
rect 120322 582684 120362 582726
rect 120328 582680 120362 582684
rect 120294 582644 120314 582646
rect 112218 582016 112252 582606
rect 113020 582588 113674 582612
rect 115972 582402 116420 582430
rect 115972 582218 116438 582402
rect 115990 582190 116438 582218
rect 118796 582086 118830 582612
rect 118566 582066 118904 582086
rect 118796 582058 118830 582066
rect 118594 582038 118904 582058
rect 118796 582010 118830 582038
rect 118910 582034 118944 582612
rect 118950 582066 119052 582086
rect 119556 582066 119662 582086
rect 118950 582038 119052 582058
rect 119556 582038 119662 582058
rect 118850 582014 119308 582034
rect 118850 582010 119348 582014
rect 119668 582010 119702 582612
rect 120290 582606 120362 582644
rect 120294 582542 120314 582606
rect 120322 582542 120362 582606
rect 120420 582542 120422 582570
rect 120328 582066 120362 582542
rect 120392 582514 120394 582542
rect 120392 582066 120400 582514
rect 120278 582010 120289 582021
rect 112302 581954 120289 582010
rect 120294 581976 120314 582066
rect 120322 582016 120362 582066
rect 120420 582038 120428 582542
rect 120322 582004 120342 582016
rect 120294 581964 120314 581966
rect 117906 581948 118162 581954
rect 112218 581896 112252 581930
rect 117934 581920 118134 581934
rect 118796 581896 118830 581954
rect 118850 581942 119348 581954
rect 119655 581942 119656 581943
rect 118890 581922 119348 581942
rect 119656 581941 119657 581942
rect 118910 581896 118944 581922
rect 119668 581896 119702 581954
rect 119714 581942 119715 581943
rect 119713 581941 119714 581942
rect 120290 581926 120362 581964
rect 120294 581900 120314 581926
rect 120322 581900 120362 581926
rect 120290 581896 120362 581900
rect 120430 581896 120464 582726
rect 112171 581862 120464 581896
rect 112218 581752 112252 581862
rect 112116 581666 112252 581752
rect 112116 581268 112150 581666
rect 112218 581362 112252 581666
rect 112258 581390 112806 581424
rect 112258 581362 112292 581390
rect 112772 581362 112806 581390
rect 112212 581346 112292 581362
rect 112258 581334 112292 581346
rect 112184 581318 112292 581334
rect 112738 581330 112840 581362
rect 112856 581348 113494 581478
rect 112856 581330 113646 581348
rect 117906 581336 117920 581414
rect 117934 581336 117948 581414
rect 118796 581330 118830 581862
rect 118910 581330 118944 581862
rect 118955 581342 118956 581343
rect 119656 581342 119657 581343
rect 118956 581341 118957 581342
rect 119655 581341 119656 581342
rect 119668 581330 119702 581862
rect 120328 581414 120362 581862
rect 120392 581414 120404 581862
rect 119713 581342 119714 581343
rect 119714 581341 119715 581342
rect 120278 581330 120289 581341
rect 112116 581190 112252 581268
rect 112116 580223 112150 581190
rect 112218 580700 112252 581190
rect 112258 581108 112292 581318
rect 112302 581296 112806 581330
rect 112322 581266 112394 581296
rect 112444 581284 112620 581296
rect 112444 581276 112631 581284
rect 112632 581266 112704 581296
rect 112360 581232 112394 581266
rect 112620 581222 112631 581233
rect 112670 581232 112704 581266
rect 112444 581188 112631 581222
rect 112662 581212 112666 581232
rect 112634 581184 112666 581204
rect 112772 581108 112806 581296
rect 112258 581074 112806 581108
rect 112856 581296 114976 581330
rect 118762 581296 120289 581330
rect 120294 581318 120314 581414
rect 120322 581358 120362 581414
rect 120420 581386 120464 581862
rect 120322 581346 120342 581358
rect 120294 581306 120314 581308
rect 112856 581274 113646 581296
rect 112856 581016 113494 581274
rect 112258 580914 112806 580948
rect 112258 580632 112292 580914
rect 112620 580834 112631 580845
rect 112322 580790 112394 580828
rect 112444 580800 112631 580834
rect 112632 580790 112704 580828
rect 112360 580756 112394 580790
rect 112404 580756 112660 580780
rect 112670 580756 112704 580790
rect 112620 580752 112631 580756
rect 112432 580728 112632 580752
rect 112444 580712 112631 580728
rect 112772 580666 112806 580914
rect 112298 580638 112806 580666
rect 112772 580632 112806 580638
rect 112258 580598 112806 580632
rect 112856 580540 113494 581002
rect 118796 580672 118830 581296
rect 118910 580672 118944 581296
rect 118956 581284 118957 581285
rect 119655 581284 119656 581285
rect 118955 581283 118956 581284
rect 119656 581283 119657 581284
rect 118955 580684 118956 580685
rect 119656 580684 119657 580685
rect 118956 580683 118957 580684
rect 119655 580683 119656 580684
rect 119668 580672 119702 581296
rect 119714 581284 119715 581285
rect 119713 581283 119714 581284
rect 120290 581268 120362 581306
rect 120294 581204 120314 581268
rect 120322 581204 120362 581268
rect 120328 580756 120362 581204
rect 120392 580856 120400 581204
rect 120420 580856 120428 581232
rect 119713 580684 119714 580685
rect 119714 580683 119715 580684
rect 120278 580672 120289 580683
rect 118762 580638 120289 580672
rect 120294 580660 120314 580756
rect 120322 580700 120368 580756
rect 120322 580688 120342 580700
rect 120356 580688 120368 580700
rect 120384 580660 120396 580756
rect 120294 580648 120314 580650
rect 118796 580223 118830 580638
rect 118910 580223 118944 580638
rect 118956 580626 118957 580627
rect 119655 580626 119656 580627
rect 118955 580625 118956 580626
rect 119656 580625 119657 580626
rect 119668 580223 119702 580638
rect 119714 580626 119715 580627
rect 119713 580625 119714 580626
rect 120290 580622 120362 580648
rect 120290 580610 120368 580622
rect 120294 580540 120314 580610
rect 120322 580540 120368 580610
rect 120384 580540 120396 580650
rect 120328 580223 120362 580540
rect 112080 580192 120395 580223
rect 103516 578484 108216 578518
rect 103516 578416 105954 578484
rect 106182 578416 106216 578484
rect 106410 578454 106444 578484
rect 106284 578416 106542 578454
rect 106754 578447 106792 578454
rect 106868 578450 106902 578484
rect 106754 578432 106800 578447
rect 106742 578416 106800 578432
rect 103516 578382 106800 578416
rect 106804 578382 106836 578416
rect 103516 577988 105954 578382
rect 106182 578366 106216 578382
rect 106156 578343 106216 578366
rect 106284 578344 106342 578382
rect 106156 578332 106235 578343
rect 106182 577988 106250 578332
rect 106274 577988 106286 577994
rect 106296 577988 106341 578344
rect 102856 577952 106382 577988
rect 102794 577918 106382 577952
rect 102794 576338 102828 577918
rect 102856 577590 106382 577918
rect 106410 577590 106444 578382
rect 106742 578344 106800 578382
rect 106838 578366 106902 578450
rect 106838 578348 106916 578366
rect 106754 577778 106788 578344
rect 106754 577604 106794 577778
rect 106754 577602 106799 577604
rect 106780 577590 106794 577602
rect 102856 577518 106764 577590
rect 106808 577562 106822 577750
rect 102856 577450 106382 577518
rect 106410 577450 106444 577518
rect 106868 577512 106916 578348
rect 106868 577450 106902 577512
rect 102856 577416 106902 577450
rect 102856 576718 106382 577416
rect 106410 576718 106444 577416
rect 102856 576684 106444 576718
rect 102856 576338 106382 576684
rect 106410 576584 106444 576684
rect 101119 576304 106382 576338
rect 101119 576286 101194 576304
rect 101119 576256 101153 576286
rect 101119 575900 101159 576256
rect 101160 576200 101194 576286
rect 101225 576286 101270 576304
rect 101160 575900 101215 576200
rect 101225 575900 101259 576286
rect 101339 576236 101373 576304
rect 102435 576283 102469 576304
rect 102794 576296 102828 576304
rect 102856 576296 106382 576304
rect 101777 576252 101824 576283
rect 101765 576236 101824 576252
rect 101904 576236 101951 576283
rect 102435 576252 102482 576283
rect 102423 576236 102482 576252
rect 102562 576236 102609 576283
rect 102794 576246 106382 576296
rect 102794 576240 102828 576246
rect 102856 576240 106382 576246
rect 102794 576236 106382 576240
rect 101320 576202 101951 576236
rect 101994 576202 102609 576236
rect 102652 576202 106382 576236
rect 101274 576154 101293 576159
rect 101305 576154 101308 576159
rect 101263 576143 101308 576154
rect 101274 575900 101308 576143
rect 101339 575900 101373 576202
rect 101765 576155 101823 576202
rect 101777 575900 101811 576155
rect 101854 576150 101864 576196
rect 101910 576150 101920 576196
rect 102423 576155 102481 576202
rect 101898 575958 101920 576150
rect 101921 576143 101966 576154
rect 101854 575900 101864 575958
rect 101910 575900 101920 575958
rect 101932 575900 101966 576143
rect 102435 575900 102469 576155
rect 102506 575900 102526 576196
rect 102562 576154 102582 576196
rect 102794 576190 106382 576202
rect 102562 576143 102624 576154
rect 102562 575900 102582 576143
rect 102590 575900 102624 576143
rect 96612 575895 102756 575900
rect 87787 574100 87832 575874
rect 87848 574858 87876 575340
rect 87848 574658 87892 574858
rect 87848 574100 87876 574658
rect 87904 574630 87920 574886
rect 87969 574100 88014 575874
rect 88445 574100 88490 575874
rect 88508 575608 102756 575895
rect 102794 575608 102828 576190
rect 102856 575608 106382 576190
rect 106390 575716 108348 576584
rect 108450 576450 108464 576816
rect 108490 576176 108506 576362
rect 109172 576342 109206 576376
rect 109286 576342 109320 576452
rect 109938 576342 109972 576456
rect 111482 576420 111516 576456
rect 110052 576342 110086 576376
rect 110710 576342 110744 576376
rect 111124 576342 111516 576420
rect 111993 576454 112027 580091
rect 112080 580042 120400 580192
rect 112080 580002 120396 580042
rect 112080 579992 120395 580002
rect 112080 579990 120396 579992
rect 112080 579384 120400 579990
rect 120420 579412 120422 579466
rect 112080 579242 120395 579384
rect 120430 579266 120464 581386
rect 120420 579242 120466 579266
rect 120472 579242 120490 579302
rect 121178 579242 121224 579266
rect 112080 579208 120464 579242
rect 122828 579214 122840 579266
rect 124929 579221 133367 583954
rect 134178 583950 134378 583952
rect 136288 583850 142208 593850
rect 142248 593810 142249 593811
rect 142247 593809 142248 593810
rect 136234 583846 142208 583850
rect 136288 583717 142208 583846
rect 134239 583686 142208 583717
rect 142496 593798 142574 595804
rect 142677 595400 142725 599555
rect 142805 599565 142839 599617
rect 143463 599596 143497 599617
rect 143421 599565 143497 599596
rect 143520 599596 143531 599614
rect 144121 599596 144155 599617
rect 144779 599596 144813 599617
rect 145042 599596 145254 599617
rect 145437 599596 145471 599617
rect 146095 599596 146129 599617
rect 142805 599468 142851 599565
rect 143421 599549 143509 599565
rect 143520 599549 146129 599596
rect 146208 599555 146279 599944
rect 142853 599522 143509 599549
rect 143511 599522 144167 599549
rect 142853 599515 144167 599522
rect 144169 599522 144825 599549
rect 144827 599522 145483 599549
rect 144169 599515 145483 599522
rect 145485 599515 146129 599549
rect 142880 599509 142908 599515
rect 143370 599509 143433 599515
rect 143457 599481 143461 599515
rect 143463 599509 143566 599515
rect 144028 599509 144080 599515
rect 143463 599468 143509 599509
rect 142805 599456 142839 599468
rect 143438 599456 143451 599467
rect 143463 599456 143497 599468
rect 142791 598812 142839 599456
rect 143449 598812 143497 599456
rect 143520 598812 143531 599509
rect 144121 599468 144167 599515
rect 144188 599509 144228 599515
rect 144690 599509 144749 599515
rect 144773 599481 144777 599515
rect 144779 599509 144898 599515
rect 144779 599468 144825 599509
rect 144096 599456 144109 599467
rect 144121 599456 144166 599468
rect 144754 599456 144767 599467
rect 144779 599456 144824 599468
rect 142791 598140 142850 598812
rect 143449 598140 143508 598812
rect 144107 598140 144166 599456
rect 144688 598140 144690 598278
rect 144716 598140 144718 598278
rect 144765 598140 144824 599456
rect 145042 599288 145254 599515
rect 145360 599509 145400 599515
rect 145437 599468 145483 599515
rect 145508 599509 145550 599515
rect 146012 599509 146065 599515
rect 146089 599481 146093 599515
rect 145412 599456 145425 599467
rect 145437 599456 145482 599468
rect 146070 599456 146083 599467
rect 146095 599456 146129 599515
rect 145028 598964 145368 599288
rect 145423 598140 145482 599456
rect 146010 598140 146012 598278
rect 146038 598140 146040 598278
rect 146081 598140 146129 599456
rect 142791 598093 146129 598140
rect 142791 597991 142850 598093
rect 142855 598059 143508 598093
rect 143525 598059 144166 598093
rect 142855 598053 142873 598059
rect 143437 598043 143508 598059
rect 144095 598043 144166 598059
rect 144171 598059 144824 598093
rect 144841 598059 145482 598093
rect 144171 598053 144189 598059
rect 143449 597991 143508 598043
rect 144107 597991 144166 598043
rect 144688 597991 144690 598053
rect 144716 597991 144718 598053
rect 144753 598043 144824 598059
rect 145411 598043 145482 598059
rect 145487 598059 146129 598093
rect 145487 598053 145505 598059
rect 144765 597991 144824 598043
rect 145423 597991 145482 598043
rect 146010 597991 146012 598053
rect 146038 597991 146040 598053
rect 146069 598043 146129 598059
rect 146081 597991 146129 598043
rect 146162 597991 146166 598198
rect 142779 597957 146166 597991
rect 142791 596997 142850 597957
rect 143449 596997 143508 597957
rect 144107 596997 144166 597957
rect 144688 597788 144690 597957
rect 144716 597816 144718 597957
rect 144765 596997 144824 597957
rect 145423 596997 145482 597957
rect 146010 597758 146012 597957
rect 146038 597786 146040 597957
rect 146081 596997 146129 597957
rect 146162 597786 146166 597957
rect 142779 596963 146163 596997
rect 142791 596960 142850 596963
rect 143449 596960 143508 596963
rect 142791 596895 142839 596960
rect 143449 596942 143497 596960
rect 143421 596895 143497 596942
rect 143520 596942 143531 596960
rect 144107 596942 144166 596963
rect 144765 596942 144824 596963
rect 145423 596942 145482 596963
rect 146081 596942 146129 596963
rect 143520 596895 146129 596942
rect 142791 596861 142850 596895
rect 142853 596861 143508 596895
rect 143511 596861 144166 596895
rect 144169 596861 144824 596895
rect 144827 596861 145482 596895
rect 145485 596861 146129 596895
rect 142791 595498 142839 596861
rect 143449 595498 143497 596861
rect 142791 595400 142825 595498
rect 143449 595486 143483 595498
rect 143486 595486 143497 595498
rect 143520 595486 143531 596861
rect 144107 595498 144166 596861
rect 144107 595486 144141 595498
rect 144688 595486 144690 596424
rect 144716 595486 144718 596424
rect 144765 595498 144824 596861
rect 145423 595498 145482 596861
rect 144765 595486 144799 595498
rect 145423 595486 145457 595498
rect 146010 595486 146012 596424
rect 146038 595486 146040 596424
rect 146081 595498 146129 596861
rect 146195 596720 146279 599555
rect 146358 597734 146392 600430
rect 146476 599600 146502 599606
rect 146504 599600 146530 599634
rect 146884 599542 147346 600180
rect 147762 599656 147796 600430
rect 147874 599656 147910 600430
rect 147920 599656 147921 600430
rect 148534 600134 148568 600430
rect 148532 599868 148574 600134
rect 148532 599754 148579 599868
rect 148588 599810 148602 600134
rect 148632 599868 148666 600430
rect 148534 599656 148579 599754
rect 148632 599656 148677 599868
rect 149192 599656 149237 600430
rect 149262 599656 149298 600134
rect 149318 599656 149354 600134
rect 149390 599656 149435 600430
rect 149850 599656 149895 600430
rect 150148 599656 150193 600430
rect 150508 599868 150542 600430
rect 150906 599868 150940 600430
rect 151166 599868 151200 600430
rect 150508 599656 150553 599868
rect 150906 599656 150951 599868
rect 151166 599656 151211 599868
rect 151280 599656 151314 600430
rect 153938 599687 153972 600430
rect 147748 599622 151314 599656
rect 146942 599458 147292 599492
rect 146942 599006 146976 599458
rect 147062 599424 147154 599428
rect 147062 599390 147168 599424
rect 147100 599356 147168 599390
rect 147104 599318 147150 599356
rect 147045 599306 147101 599317
rect 147056 599130 147101 599306
rect 147116 599306 147150 599318
rect 147162 599306 147189 599317
rect 147116 599130 147189 599306
rect 147116 599118 147150 599130
rect 147062 599114 147154 599118
rect 147062 599080 147168 599114
rect 147100 599046 147168 599080
rect 147104 599030 147150 599046
rect 147258 599006 147292 599458
rect 147748 599006 147796 599622
rect 147874 599592 147910 599622
rect 147920 599592 147921 599622
rect 148120 599592 148332 599622
rect 148534 599592 148579 599622
rect 148632 599592 148677 599622
rect 148786 599592 148998 599622
rect 149192 599592 149237 599622
rect 149248 599592 149298 599622
rect 149318 599592 149354 599622
rect 149390 599592 149646 599622
rect 149850 599592 149895 599622
rect 150148 599592 150193 599622
rect 150508 599592 150553 599622
rect 150906 599592 150951 599622
rect 147874 599554 148530 599592
rect 147874 599514 147921 599554
rect 147924 599520 148530 599554
rect 148534 599554 149188 599592
rect 148534 599522 148579 599554
rect 148582 599522 149188 599554
rect 148534 599520 149188 599522
rect 149192 599554 149846 599592
rect 147948 599514 147970 599520
rect 147851 599470 147862 599481
rect 147874 599470 147948 599514
rect 147862 599466 147948 599470
rect 147970 599466 147976 599514
rect 147862 599006 147921 599466
rect 148120 599368 148332 599520
rect 148534 599514 148678 599520
rect 148534 599481 148579 599514
rect 148620 599482 148678 599514
rect 148509 599470 148579 599481
rect 148520 599466 148579 599470
rect 148626 599466 148630 599482
rect 148520 599458 148626 599466
rect 148098 599006 148420 599368
rect 148520 599006 148579 599458
rect 148632 599006 148677 599482
rect 148786 599368 148998 599520
rect 149192 599510 149237 599554
rect 149240 599520 149846 599554
rect 149850 599554 150504 599592
rect 149298 599514 149304 599520
rect 149248 599510 149298 599514
rect 149174 599481 149298 599510
rect 149167 599470 149298 599481
rect 149174 599466 149298 599470
rect 149304 599466 149354 599514
rect 149378 599482 149646 599520
rect 149174 599368 149248 599466
rect 149298 599458 149304 599466
rect 148786 599196 149248 599368
rect 148888 599006 149248 599196
rect 149390 599380 149646 599482
rect 149850 599481 149895 599554
rect 149898 599520 150504 599554
rect 150508 599554 151162 599592
rect 150136 599482 150194 599520
rect 150508 599502 150553 599554
rect 150556 599520 151162 599554
rect 149825 599470 149895 599481
rect 149836 599380 149895 599470
rect 149390 599200 149936 599380
rect 149390 599006 149435 599200
rect 149614 599006 149936 599200
rect 150148 599006 150193 599482
rect 150490 599481 150564 599502
rect 150894 599482 150952 599520
rect 150483 599470 150564 599481
rect 150490 599402 150564 599470
rect 150360 599006 150682 599402
rect 150906 599006 150951 599482
rect 151166 599481 151211 599622
rect 151141 599470 151211 599481
rect 151152 599006 151211 599470
rect 151266 599006 151314 599622
rect 151397 599006 155021 599687
rect 156470 599006 156498 599690
rect 157738 599656 157762 600430
rect 157772 599656 157796 600430
rect 159551 599656 167989 600430
rect 146942 598944 156498 599006
rect 146970 598936 156498 598944
rect 156504 599622 167989 599656
rect 146314 597712 146434 597734
rect 146314 597586 146726 597712
rect 146320 597182 146726 597586
rect 146358 596872 146392 597182
rect 146970 596720 156478 598936
rect 156504 597002 156538 599622
rect 157738 599592 157762 599622
rect 157772 599592 157796 599622
rect 159244 599592 159278 599622
rect 159551 599592 167989 599622
rect 156970 599570 157008 599592
rect 156958 599554 157016 599570
rect 157248 599554 157286 599592
rect 157728 599570 157766 599592
rect 157772 599570 157944 599592
rect 157716 599554 157944 599570
rect 157958 599554 158602 599592
rect 158616 599554 167989 599592
rect 156680 599520 157286 599554
rect 157338 599520 157944 599554
rect 157996 599520 158602 599554
rect 156958 599482 157016 599520
rect 157716 599482 157796 599520
rect 158474 599514 158576 599520
rect 158642 599514 158648 599522
rect 158654 599520 159284 599554
rect 159172 599514 159284 599520
rect 159300 599520 167989 599554
rect 159300 599514 159376 599520
rect 158474 599482 158532 599514
rect 156607 599470 156652 599481
rect 156618 597002 156652 599470
rect 156970 597002 157004 599482
rect 157265 599470 157310 599481
rect 157276 597002 157310 599470
rect 157728 597002 157762 599482
rect 157772 598370 157796 599482
rect 157923 599470 157979 599481
rect 157934 598370 157979 599470
rect 157828 597550 157850 597854
rect 157884 597550 157906 597854
rect 157934 597002 157968 598370
rect 158486 598346 158531 599482
rect 158620 599481 158632 599482
rect 158581 599470 158637 599481
rect 158592 598346 158637 599470
rect 158648 599466 158660 599510
rect 159232 599486 159284 599514
rect 159232 599482 159238 599486
rect 159244 599470 159278 599486
rect 158486 597002 158520 598346
rect 158592 597784 158626 598346
rect 158558 597002 158570 597784
rect 158586 597002 158632 597784
rect 158648 597489 158660 597784
rect 159244 597489 159284 599470
rect 159290 597489 159295 599481
rect 159551 598315 167989 599520
rect 159908 597786 159942 598315
rect 159874 597489 159900 597786
rect 159902 597489 159948 597786
rect 159962 597489 159976 597786
rect 160022 597489 160056 598315
rect 165192 597489 165202 597684
rect 165220 597489 165230 597656
rect 158648 597002 167097 597489
rect 156504 596968 167097 597002
rect 156504 596720 156538 596968
rect 156618 596860 156652 596968
rect 156970 596938 157004 596968
rect 157276 596938 157310 596968
rect 156970 596900 157008 596938
rect 157248 596900 157310 596938
rect 157728 596938 157762 596968
rect 157934 596938 157968 596968
rect 157728 596900 157766 596938
rect 157906 596900 157968 596938
rect 158486 596938 158520 596968
rect 158586 596938 158632 596968
rect 158486 596900 158524 596938
rect 158564 596906 158632 596938
rect 158648 596906 167097 596968
rect 158558 596900 158632 596906
rect 158642 596900 167097 596906
rect 156664 596866 157310 596900
rect 157322 596866 157968 596900
rect 157980 596866 158632 596900
rect 158638 596866 167097 596900
rect 169856 596872 169890 600430
rect 171421 598228 173072 600430
rect 171421 598208 173150 598228
rect 171421 598200 173072 598208
rect 171421 598180 173122 598200
rect 171421 598125 173072 598180
rect 171421 598091 175456 598125
rect 171421 597941 173072 598091
rect 171732 597940 172280 597941
rect 172330 597886 172968 597941
rect 172262 597774 172266 597776
rect 172904 597556 172922 597714
rect 172942 597590 172960 597676
rect 173002 597556 173036 597941
rect 172904 597552 173122 597556
rect 172922 597538 173122 597552
rect 173002 597522 173036 597538
rect 172922 597504 173156 597522
rect 173002 597502 173036 597504
rect 171590 597468 175456 597502
rect 157276 596860 157310 596866
rect 157934 596860 157968 596866
rect 158558 596860 158576 596866
rect 158586 596860 158632 596866
rect 158642 596860 167097 596866
rect 156606 596822 156664 596860
rect 156942 596822 156980 596860
rect 157264 596822 157322 596860
rect 157700 596822 157738 596860
rect 157922 596822 157980 596860
rect 158458 596822 158496 596860
rect 158580 596828 158638 596860
rect 158648 596828 167097 596860
rect 156606 596788 156980 596822
rect 157032 596788 157738 596822
rect 157790 596788 158496 596822
rect 158536 596822 158638 596828
rect 158659 596822 167097 596828
rect 158536 596788 167097 596822
rect 168278 596804 168324 596828
rect 156606 596772 156664 596788
rect 157264 596772 157322 596788
rect 157922 596772 157980 596788
rect 158536 596782 158564 596788
rect 158580 596772 158638 596788
rect 156606 596757 156652 596772
rect 156618 596720 156652 596757
rect 157276 596720 157310 596772
rect 157934 596720 157968 596772
rect 158592 596720 158626 596772
rect 158659 596720 167097 596788
rect 168286 596782 168324 596804
rect 168342 596754 168352 596856
rect 171590 596822 171624 597468
rect 172130 597388 172164 597468
rect 172292 597388 172876 597399
rect 172888 597388 172922 597468
rect 173002 597388 173036 597468
rect 179764 597394 179780 597500
rect 171654 597326 171726 597364
rect 171776 597354 173070 597388
rect 172117 597342 172118 597343
rect 172118 597341 172119 597342
rect 171692 596822 171726 597326
rect 172130 596872 172164 597354
rect 172176 597342 172177 597343
rect 172875 597342 172876 597343
rect 172888 597342 172922 597354
rect 172175 597341 172176 597342
rect 172876 597341 172877 597342
rect 172888 597078 172933 597342
rect 173002 597078 173036 597354
rect 179754 597348 179780 597394
rect 179764 597270 179780 597348
rect 179782 597320 179792 597422
rect 179782 597276 179796 597298
rect 179754 597248 179796 597270
rect 171763 596860 171764 596861
rect 171764 596859 171765 596860
rect 172102 596822 172140 596860
rect 172438 596822 175404 597078
rect 171590 596788 172140 596822
rect 172192 596796 175404 596822
rect 171590 596720 171624 596788
rect 171692 596758 171726 596788
rect 172002 596782 172114 596788
rect 172180 596782 175404 596796
rect 172438 596768 175404 596782
rect 172030 596754 172142 596768
rect 172152 596754 175404 596768
rect 171692 596742 171726 596754
rect 171776 596720 175404 596754
rect 146195 596686 146297 596720
rect 146970 596686 175404 596720
rect 146195 596650 146279 596686
rect 146970 596650 156478 596686
rect 146081 595486 146115 595498
rect 142827 595400 142831 595473
rect 142855 595439 142859 595445
rect 143435 595439 146115 595486
rect 142851 595405 142859 595439
rect 142867 595405 143483 595439
rect 143509 595405 143517 595439
rect 143525 595405 144141 595439
rect 142855 595400 142859 595405
rect 143437 595400 143483 595405
rect 144095 595400 144141 595405
rect 144143 595400 144147 595439
rect 144171 595400 144175 595439
rect 144183 595405 144799 595439
rect 144841 595405 145457 595439
rect 142641 595337 144354 595400
rect 144688 595392 144690 595399
rect 144716 595364 144718 595399
rect 144753 595389 144799 595405
rect 145411 595389 145457 595405
rect 144765 595337 144799 595389
rect 145423 595337 145457 595389
rect 145459 595371 145463 595439
rect 145487 595399 145491 595439
rect 145499 595405 146115 595439
rect 146010 595392 146012 595399
rect 146038 595364 146040 595399
rect 146069 595389 146115 595405
rect 146081 595337 146115 595389
rect 146195 595399 146243 596650
rect 147006 596126 147040 596650
rect 147002 596092 147296 596126
rect 147006 595965 147040 596092
rect 147120 596071 147154 596092
rect 146986 595931 147040 595965
rect 147008 595755 147074 595931
rect 147086 595796 147096 595982
rect 147108 595943 147154 596071
rect 147114 595931 147154 595943
rect 147166 595931 147193 595942
rect 147114 595768 147193 595931
rect 147120 595755 147193 595768
rect 147006 595594 147040 595755
rect 147120 595743 147154 595755
rect 147108 595631 147154 595743
rect 147120 595594 147154 595631
rect 147262 595594 147296 596092
rect 147002 595560 147296 595594
rect 147712 596072 151350 596650
rect 151433 596072 151467 596650
rect 151547 596636 151592 596650
rect 151547 596124 151581 596636
rect 151734 596634 152124 596650
rect 151734 596136 151768 596634
rect 151948 596566 151995 596613
rect 151910 596532 151995 596566
rect 151837 596473 151882 596484
rect 151965 596473 152010 596484
rect 151848 596297 151882 596473
rect 151976 596297 152010 596473
rect 151948 596238 151995 596285
rect 151910 596204 151995 596238
rect 152090 596136 152124 596634
rect 151547 596100 151592 596124
rect 151734 596102 152124 596136
rect 152205 596634 152600 596650
rect 152205 596572 152250 596634
rect 152205 596198 152244 596572
rect 152416 596566 152471 596613
rect 152386 596532 152471 596566
rect 152313 596473 152358 596484
rect 152441 596473 152497 596484
rect 152324 596297 152358 596473
rect 152452 596297 152497 596473
rect 152416 596238 152471 596285
rect 152386 596204 152471 596238
rect 152205 596136 152250 596198
rect 152566 596136 152600 596634
rect 152205 596102 152600 596136
rect 152748 596514 153589 596650
rect 151488 596072 151592 596100
rect 151964 596072 152036 596100
rect 147712 596052 152058 596072
rect 152205 596052 152250 596102
rect 147712 596014 152138 596052
rect 152192 596014 152614 596052
rect 147006 595510 147040 595560
rect 142641 595303 146127 595337
rect 142496 583686 142560 593798
rect 142641 591468 144354 595303
rect 144765 591468 144799 593342
rect 145423 591468 145457 593342
rect 146081 591468 146115 593342
rect 142641 591421 146115 591468
rect 142641 591387 144805 591421
rect 142641 591319 144354 591387
rect 144731 591381 144749 591387
rect 144759 591353 144805 591387
rect 144815 591387 145463 591421
rect 144815 591381 144833 591387
rect 145389 591381 145407 591387
rect 145417 591353 145463 591387
rect 145473 591387 146115 591421
rect 145473 591381 145491 591387
rect 146047 591381 146065 591387
rect 146075 591353 146115 591387
rect 144765 591319 144799 591353
rect 145423 591319 145457 591353
rect 146081 591319 146115 591353
rect 142641 591285 146149 591319
rect 142641 588950 144354 591285
rect 146195 588727 146229 595399
rect 146970 595226 147314 595510
rect 147712 595432 152614 596014
rect 147712 595226 152510 595432
rect 152748 595226 153566 596514
rect 154179 595226 154224 596650
rect 154837 596124 154871 596650
rect 154837 596062 154882 596124
rect 154951 596062 154985 596650
rect 156294 596218 156328 596650
rect 156294 596136 156384 596218
rect 155662 596092 156052 596126
rect 154396 595512 155220 596062
rect 155662 595594 155696 596092
rect 155791 596024 155923 596071
rect 155838 595990 155923 596024
rect 155765 595931 155821 595942
rect 155893 595931 155949 595942
rect 155776 595755 155821 595931
rect 155904 595755 155949 595931
rect 155791 595696 155923 595743
rect 155838 595662 155923 595696
rect 156018 595594 156052 596092
rect 155662 595560 156052 595594
rect 154430 595226 154642 595512
rect 154822 595492 154892 595512
rect 154837 595226 154882 595492
rect 154951 595226 154985 595512
rect 155086 595426 155204 595512
rect 155648 595226 156070 595510
rect 156294 595226 156328 596136
rect 146970 595192 156340 595226
rect 146970 595171 147314 595192
rect 147712 595171 152510 595192
rect 152748 595171 153566 595192
rect 154179 595171 154224 595192
rect 146970 595124 154462 595171
rect 154837 595124 154871 595192
rect 154951 595124 154985 595192
rect 155648 595124 156070 595192
rect 156294 595171 156328 595192
rect 156266 595124 156328 595171
rect 146970 595090 156328 595124
rect 146970 594890 147314 595090
rect 147006 594374 147040 594890
rect 147006 594106 147278 594374
rect 146978 593984 147278 594106
rect 147006 593930 147278 593984
rect 147006 593472 147040 593930
rect 147002 593438 147296 593472
rect 147006 593342 147040 593438
rect 147012 593311 147040 593342
rect 146986 593277 147040 593311
rect 147108 593401 147120 593417
rect 147108 593386 147123 593401
rect 147108 593342 147136 593386
rect 147108 593289 147154 593342
rect 147120 593277 147154 593289
rect 147166 593277 147193 593288
rect 147008 593101 147074 593277
rect 147120 593101 147193 593277
rect 147006 592940 147040 593101
rect 147120 593089 147154 593101
rect 147108 592977 147154 593089
rect 147120 592940 147154 592977
rect 147262 592940 147296 593438
rect 147002 592906 147296 592940
rect 147006 592856 147040 592906
rect 146970 592787 147314 592856
rect 147712 592787 152510 595090
rect 152748 595084 153566 595090
rect 152748 592787 153589 595084
rect 154179 592787 154224 595090
rect 146970 592740 154462 592787
rect 154837 592740 154871 595090
rect 154951 592740 154985 595090
rect 155648 594890 156070 595090
rect 156294 593564 156328 595090
rect 156294 593482 156376 593564
rect 155662 593438 156052 593472
rect 155662 592940 155696 593438
rect 155876 593370 155923 593417
rect 155838 593336 155923 593370
rect 155765 593277 155810 593288
rect 155893 593277 155938 593288
rect 155776 593101 155810 593277
rect 155904 593101 155938 593277
rect 155876 593042 155923 593089
rect 155838 593008 155923 593042
rect 156018 592940 156052 593438
rect 155662 592906 156052 592940
rect 155648 592740 156070 592856
rect 156294 592787 156328 593482
rect 156266 592740 156328 592787
rect 146970 592706 156328 592740
rect 146970 592638 147314 592706
rect 147712 592650 152510 592706
rect 152748 592700 153566 592706
rect 147712 592638 152586 592650
rect 152748 592638 153589 592700
rect 154179 592638 154224 592706
rect 154837 592638 154871 592706
rect 154951 592638 154985 592706
rect 155648 592638 156070 592706
rect 156294 592638 156328 592706
rect 146970 592604 156340 592638
rect 156346 592604 156362 592638
rect 146970 592236 147314 592604
rect 147712 592118 152510 592604
rect 152552 592118 152586 592604
rect 147712 592084 152586 592118
rect 147006 591984 147040 592038
rect 147712 592034 152510 592084
rect 147104 591984 147154 592018
rect 147712 591984 152600 592034
rect 152748 591984 153589 592604
rect 154179 591984 154224 592604
rect 154837 591984 154871 592604
rect 154951 591984 154985 592604
rect 155648 592236 156070 592604
rect 156294 591984 156328 592604
rect 147042 591950 147094 591984
rect 147108 591950 156340 591984
rect 147008 591888 147040 591922
rect 147042 584024 147076 591950
rect 147108 591827 147130 591950
rect 147712 591929 152600 591950
rect 152748 591929 153589 591950
rect 154179 591929 154224 591950
rect 147171 591882 154462 591929
rect 154837 591882 154871 591950
rect 154951 591882 154985 591950
rect 156294 591929 156328 591950
rect 156294 591898 156340 591929
rect 156282 591882 156340 591898
rect 147218 591848 156340 591882
rect 147108 589055 147154 591827
rect 147166 591789 147201 591800
rect 147108 589043 147130 589055
rect 147156 589043 147201 591789
rect 147712 591468 152600 591848
rect 152748 591842 153566 591848
rect 152748 591468 153589 591842
rect 154179 591468 154224 591848
rect 154837 591468 154871 591848
rect 147712 591421 154462 591468
rect 154809 591421 154871 591468
rect 147712 591387 154224 591421
rect 154241 591387 154871 591421
rect 147712 591319 152510 591387
rect 152748 591319 153589 591387
rect 154179 591319 154224 591387
rect 154837 591319 154871 591387
rect 154951 591319 154985 591848
rect 156282 591839 156318 591848
rect 156282 591801 156328 591839
rect 147712 591285 154985 591319
rect 147712 590622 152510 591285
rect 152748 590940 153589 591285
rect 147712 589382 151336 590622
rect 151433 589382 151467 590622
rect 151547 590186 151581 590622
rect 152205 590186 152239 590622
rect 151547 589964 151592 590186
rect 152205 589996 152250 590186
rect 151547 589382 151581 589964
rect 151720 589962 152110 589996
rect 151720 589464 151754 589962
rect 151934 589894 151981 589941
rect 151896 589860 151981 589894
rect 151823 589801 151868 589812
rect 151951 589801 151996 589812
rect 151834 589625 151868 589801
rect 151962 589625 151996 589801
rect 151934 589566 151981 589613
rect 151896 589532 151981 589566
rect 152076 589464 152110 589962
rect 152196 589962 152586 589996
rect 152196 589934 152239 589962
rect 152196 589537 152264 589934
rect 152410 589894 152457 589941
rect 152372 589860 152457 589894
rect 152299 589801 152344 589812
rect 152427 589801 152483 589812
rect 152310 589625 152344 589801
rect 152438 589625 152483 589801
rect 152410 589566 152457 589613
rect 152194 589526 152264 589537
rect 152372 589532 152457 589566
rect 151720 589430 152110 589464
rect 152196 589464 152239 589526
rect 152552 589464 152586 589962
rect 152196 589430 152586 589464
rect 152748 589752 153566 590940
rect 152205 589382 152239 589430
rect 147712 589380 152520 589382
rect 147712 589348 152600 589380
rect 147712 589268 151336 589348
rect 151433 589338 151490 589348
rect 151433 589320 151467 589338
rect 151484 589320 151490 589338
rect 151388 589282 151467 589320
rect 151428 589268 151467 589282
rect 151547 589268 151581 589348
rect 151702 589268 152124 589348
rect 152178 589268 152600 589348
rect 147712 589234 152600 589268
rect 147712 589043 151336 589234
rect 151428 589230 151467 589234
rect 151428 589168 151430 589230
rect 147144 588996 151336 589043
rect 151433 588996 151467 589230
rect 151484 589168 151486 589230
rect 151547 589043 151581 589234
rect 151547 588996 151594 589043
rect 151702 588996 152124 589234
rect 152178 588996 152600 589234
rect 152748 589043 153589 589752
rect 154179 589043 154224 591285
rect 154837 589043 154871 591285
rect 152630 588996 154462 589043
rect 154837 588996 154884 589043
rect 154951 588996 154985 591285
rect 155560 591336 155950 591370
rect 155560 590838 155594 591336
rect 155774 591268 155821 591315
rect 155736 591234 155821 591268
rect 155663 591175 155708 591186
rect 155791 591175 155836 591186
rect 155674 590999 155708 591175
rect 155802 590999 155836 591175
rect 155774 590940 155821 590987
rect 155736 590906 155821 590940
rect 155916 590838 155950 591336
rect 155560 590804 155950 590838
rect 155542 590134 155964 590754
rect 156294 590746 156328 591801
rect 156330 591789 156362 591805
rect 156330 590746 156364 591789
rect 156408 590806 156442 596650
rect 156468 596124 156478 596650
rect 156468 595192 156498 596124
rect 156468 592020 156478 595192
rect 156504 592020 156538 596686
rect 156468 591950 156538 592020
rect 156444 590806 156538 591950
rect 156618 591478 156652 596686
rect 156656 595526 156658 595582
rect 156656 595270 156658 595326
rect 156656 595126 156658 595182
rect 156656 594870 156658 594926
rect 156656 592872 156690 592928
rect 156684 592672 156690 592872
rect 156712 592672 156718 592872
rect 156656 592616 156690 592672
rect 156656 592472 156690 592528
rect 156684 592272 156690 592472
rect 156712 592272 156718 592472
rect 156656 592216 156690 592272
rect 157276 591482 157310 596686
rect 157934 591482 157968 596686
rect 158552 595130 158564 596234
rect 158592 591482 158626 596686
rect 158659 596650 167097 596686
rect 158659 594690 160092 596650
rect 171590 595370 171624 596686
rect 171692 596652 171726 596684
rect 172438 596140 175404 596686
rect 175950 595644 177600 597082
rect 178036 595642 179686 597080
rect 179764 596944 179780 597248
rect 179802 596758 179836 597326
rect 179842 597276 179896 597298
rect 179842 597248 179868 597270
rect 179764 596638 179780 596642
rect 171416 595364 173724 595370
rect 169466 595334 173724 595364
rect 169516 595182 169530 595284
rect 169544 595210 169586 595256
rect 171190 595216 171412 595236
rect 171228 595178 171374 595198
rect 158659 594673 165384 594690
rect 158659 594656 160092 594673
rect 158659 594622 165446 594656
rect 158659 594542 160092 594622
rect 160570 594542 165262 594553
rect 158659 594508 165262 594542
rect 158659 594049 160092 594508
rect 165263 594480 165391 594527
rect 161860 594222 162306 594328
rect 161724 594146 162306 594222
rect 161860 594086 162306 594146
rect 160666 594060 162986 594072
rect 165310 594062 165391 594480
rect 165263 594060 165391 594062
rect 160570 594049 165391 594060
rect 165412 594049 165446 594622
rect 171416 594424 173724 595334
rect 173994 594428 176302 595376
rect 176464 594848 176720 594850
rect 176492 594820 176692 594822
rect 179764 594762 179780 594866
rect 179754 594716 179780 594762
rect 173994 594424 177600 594428
rect 158659 594015 165480 594049
rect 158659 593935 160092 594015
rect 160666 593935 160700 594015
rect 162810 593970 162857 594015
rect 160842 593969 162857 593970
rect 160826 593936 162857 593969
rect 161004 593935 161060 593936
rect 162554 593935 162610 593936
rect 162952 593935 162986 594015
rect 165263 594008 165391 594015
rect 165263 594003 165375 594008
rect 165192 593935 165304 593940
rect 165350 593935 165352 593940
rect 165412 593935 165446 594015
rect 171416 593938 177600 594424
rect 158659 593901 166965 593935
rect 171416 593932 175416 593938
rect 158659 593890 160092 593901
rect 160666 593900 160700 593901
rect 160194 593896 160828 593900
rect 160194 593890 162826 593896
rect 162838 593890 162872 593893
rect 162952 593890 162986 593901
rect 165220 593890 165304 593901
rect 158659 593889 165304 593890
rect 158659 593884 161060 593889
rect 162554 593884 165304 593889
rect 158659 593878 165304 593884
rect 165350 593878 165408 593901
rect 158659 593867 165267 593878
rect 158659 593865 160092 593867
rect 159044 592454 160092 593865
rect 160666 593850 163026 593867
rect 160666 593226 160700 593850
rect 160780 593226 160814 593850
rect 162770 593844 162832 593850
rect 160826 593838 160827 593839
rect 160825 593837 160826 593838
rect 162798 593816 162832 593842
rect 162838 593800 162872 593850
rect 162878 593844 163026 593850
rect 162952 593842 162986 593844
rect 162878 593816 162998 593842
rect 162952 593800 162986 593816
rect 162836 593752 162986 593800
rect 162826 593682 162986 593752
rect 161870 593428 162316 593670
rect 162826 593450 162886 593682
rect 161990 593342 162230 593428
rect 161004 593274 161060 593288
rect 162700 593274 162756 593288
rect 160825 593238 160826 593239
rect 162826 593238 162827 593239
rect 162838 593238 162872 593450
rect 160826 593237 160827 593238
rect 161004 593226 161060 593232
rect 162300 593226 162920 593238
rect 162952 593226 162986 593682
rect 165412 593342 165446 593901
rect 171684 593748 171718 593932
rect 172438 593914 175404 593932
rect 175950 593914 177600 593938
rect 178036 593914 179686 594426
rect 179764 594290 179780 594716
rect 179782 594688 179792 594790
rect 179802 594784 179836 595352
rect 179802 594126 179836 594694
rect 180084 594290 180094 594514
rect 180084 593984 180094 593988
rect 173424 593886 173720 593914
rect 174768 593886 175064 593914
rect 175986 593800 176020 593914
rect 176342 593912 176594 593914
rect 176376 593878 176598 593882
rect 176088 593800 176118 593818
rect 171476 593714 172300 593748
rect 160666 593224 162986 593226
rect 160666 593192 163536 593224
rect 160666 592650 160700 593192
rect 160780 592840 160814 593192
rect 160826 593180 160827 593181
rect 160825 593179 160826 593180
rect 162300 592976 162920 593192
rect 161870 592958 162920 592976
rect 161614 592844 162920 592958
rect 160780 592650 160825 592840
rect 161870 592816 162920 592844
rect 162952 593190 163536 593192
rect 162952 592868 163004 593190
rect 163502 593176 163536 593190
rect 163342 593166 164382 593176
rect 163341 593110 163352 593121
rect 163025 593048 163106 593095
rect 163165 593076 163352 593110
rect 163353 593048 163434 593095
rect 163072 593010 163106 593048
rect 163400 593010 163434 593048
rect 163341 592982 163352 592993
rect 163165 592948 163352 592982
rect 163502 592868 163536 593166
rect 162952 592834 163536 592868
rect 164226 592900 165482 592936
rect 169370 592900 169404 593342
rect 164226 592866 169582 592900
rect 161870 592734 162316 592816
rect 160476 592616 160866 592650
rect 160476 592568 160510 592616
rect 160666 592582 160700 592616
rect 160618 592581 160700 592582
rect 160605 592568 160700 592581
rect 160780 592568 160814 592616
rect 160825 592580 160826 592581
rect 160826 592579 160827 592580
rect 160832 592568 160866 592616
rect 160952 592616 161342 592650
rect 160952 592568 160986 592616
rect 161094 592581 161200 592582
rect 161081 592568 161213 592581
rect 161308 592568 161342 592616
rect 162826 592580 162827 592581
rect 162825 592579 162826 592580
rect 162158 592568 162376 592579
rect 162706 592568 162756 592574
rect 162838 592568 162872 592816
rect 162952 592568 162986 592834
rect 164226 592568 165482 592866
rect 160476 592534 165482 592568
rect 160476 592462 160510 592534
rect 160621 592522 160724 592534
rect 160666 592514 160724 592522
rect 160780 592521 160814 592534
rect 160278 592454 160568 592462
rect 160590 592454 160624 592488
rect 160666 592454 160700 592514
rect 160768 592495 160818 592521
rect 160754 592494 160818 592495
rect 160746 592488 160754 592494
rect 160718 592467 160754 592488
rect 160718 592462 160758 592467
rect 160768 592462 160818 592494
rect 160832 592462 160866 592534
rect 160952 592462 160986 592534
rect 161004 592494 161060 592518
rect 161128 592514 161213 592534
rect 161066 592466 161100 592488
rect 161194 592466 161228 592488
rect 161055 592462 161100 592466
rect 160718 592454 160752 592462
rect 160754 592454 160818 592462
rect 160820 592455 161100 592462
rect 161183 592455 161228 592466
rect 160820 592454 161060 592455
rect 161066 592454 161100 592455
rect 161194 592454 161228 592455
rect 161308 592454 161342 592534
rect 162158 592468 162376 592488
rect 162838 592454 162872 592534
rect 162952 592454 162986 592534
rect 164226 592454 165482 592534
rect 159044 592420 165482 592454
rect 159044 592418 160092 592420
rect 160476 592418 160510 592420
rect 160666 592418 160700 592420
rect 160718 592418 160734 592420
rect 160742 592418 160752 592420
rect 160768 592418 160818 592420
rect 160832 592418 160866 592420
rect 160952 592418 160986 592420
rect 161066 592418 161100 592420
rect 161194 592418 161228 592420
rect 161308 592418 161342 592420
rect 162952 592418 162986 592420
rect 164226 592418 165482 592420
rect 159044 592384 165482 592418
rect 159250 592382 159284 592384
rect 159908 592382 159942 592384
rect 160022 592382 160056 592384
rect 160440 592382 163022 592384
rect 164262 592382 164296 592384
rect 164376 592382 164410 592384
rect 158718 592348 167066 592382
rect 158718 591482 158752 592348
rect 159160 592274 159172 592332
rect 159188 592274 159200 592304
rect 159250 592268 159284 592348
rect 159908 592268 159942 592348
rect 160022 592268 160056 592348
rect 158782 592206 158854 592244
rect 158904 592234 160056 592268
rect 158820 591638 158854 592206
rect 159160 592168 159172 592228
rect 159188 592196 159200 592228
rect 159237 592222 159238 592223
rect 159238 592221 159239 592222
rect 159250 592062 159284 592234
rect 159296 592222 159297 592223
rect 159895 592222 159896 592223
rect 159295 592221 159296 592222
rect 159896 592221 159897 592222
rect 159908 592062 159942 592234
rect 160022 592062 160056 592234
rect 160440 592062 163022 592348
rect 164262 592268 164296 592348
rect 164376 592268 164410 592348
rect 164422 592268 166891 592279
rect 164262 592234 166891 592268
rect 164262 592062 164296 592234
rect 164376 592222 164410 592234
rect 164422 592222 164423 592223
rect 164376 592221 164422 592222
rect 164376 592062 164421 592221
rect 166892 592206 167002 592244
rect 159044 591926 165482 592062
rect 166892 591926 166893 591927
rect 166930 591926 167002 592206
rect 159044 591888 166892 591926
rect 166930 591888 166964 591926
rect 167032 591888 167066 592348
rect 159044 591854 167066 591888
rect 159044 591786 165482 591854
rect 166930 591786 166964 591854
rect 167032 591786 167066 591854
rect 169370 591786 169404 592866
rect 169406 592764 169438 592798
rect 169456 592726 169464 592856
rect 169472 592726 169506 592752
rect 169441 592714 169506 592726
rect 169434 592220 169506 592714
rect 169434 592189 169480 592220
rect 169434 592182 169468 592189
rect 169434 592168 169438 592182
rect 169434 592130 169480 592168
rect 169434 591938 169506 592130
rect 169516 592124 169530 592226
rect 169548 592198 169582 592866
rect 171476 592716 171510 593714
rect 171594 593662 171632 593704
rect 171556 593574 171582 593596
rect 171602 593578 171622 593662
rect 171636 593652 171674 593662
rect 171636 593630 171678 593652
rect 171684 593630 171718 593714
rect 171636 593606 171718 593630
rect 171614 593574 171616 593578
rect 171636 593574 171674 593606
rect 171556 593562 171654 593574
rect 171578 592716 171650 593562
rect 171684 592716 171718 593606
rect 172630 593486 173622 593784
rect 173940 593486 174932 593792
rect 175108 593486 175404 593800
rect 175950 593534 176118 593800
rect 176268 593722 177600 593804
rect 178036 593722 179686 593804
rect 176212 593700 177726 593722
rect 177918 593700 179694 593722
rect 176212 593698 177746 593700
rect 177756 593698 179720 593700
rect 176212 593690 177726 593698
rect 177918 593690 179694 593698
rect 175806 593532 176118 593534
rect 176268 593672 177600 593690
rect 178036 593672 179686 593690
rect 176268 593670 177718 593672
rect 177784 593670 179692 593672
rect 176268 593666 177600 593670
rect 178036 593666 179686 593670
rect 176268 593662 177726 593666
rect 177918 593662 179722 593666
rect 175806 593498 176134 593532
rect 176268 593498 177600 593662
rect 175154 593480 175178 593486
rect 175270 593480 175292 593486
rect 175208 593446 175232 593480
rect 175246 593446 175756 593480
rect 175174 593384 175178 593418
rect 172734 593314 172820 593342
rect 172648 593298 172820 593314
rect 172648 593160 172802 593298
rect 175208 593164 175242 593446
rect 175246 593360 175296 593446
rect 175383 593366 175581 593377
rect 175246 593322 175382 593360
rect 175394 593332 175581 593366
rect 175582 593322 175692 593360
rect 175246 593272 175304 593322
rect 175310 593288 175382 593322
rect 175383 593278 175581 593289
rect 175620 593288 175692 593322
rect 175246 593164 175296 593272
rect 175394 593244 175581 593278
rect 175722 593164 175756 593446
rect 175208 593130 175232 593164
rect 175246 593130 175756 593164
rect 175806 593464 177600 593498
rect 175806 593384 176134 593464
rect 176213 593384 176224 593395
rect 175806 593350 176224 593384
rect 176268 593369 177600 593464
rect 175806 593256 176134 593350
rect 176146 593338 176147 593339
rect 176145 593337 176146 593338
rect 176225 593322 177600 593369
rect 176145 593268 176146 593269
rect 176146 593267 176147 593268
rect 176213 593256 176224 593267
rect 175806 593222 176224 593256
rect 175806 593221 176134 593222
rect 175806 593210 176100 593221
rect 175806 593209 176118 593210
rect 175806 593114 176100 593209
rect 176268 593176 177600 593322
rect 176162 593162 177600 593176
rect 176268 593142 177600 593162
rect 176135 593131 177600 593142
rect 176146 593114 177600 593131
rect 175806 593108 177600 593114
rect 175806 593072 176100 593108
rect 175950 592990 176100 593072
rect 176268 592990 177600 593108
rect 173976 592722 174010 592740
rect 171416 592431 172432 592716
rect 172630 592431 173622 592716
rect 173976 592686 174932 592722
rect 173654 592431 173688 592584
rect 173994 592467 174932 592686
rect 173940 592431 174932 592467
rect 175108 592498 176100 592722
rect 176112 592498 176116 592503
rect 175108 592431 176116 592498
rect 176118 592431 176152 592465
rect 176232 592431 176266 592590
rect 176268 592467 176302 592722
rect 176304 592467 176320 592740
rect 176418 592467 176452 592990
rect 178036 592988 179686 593662
rect 178400 592974 179196 592988
rect 180176 592721 180210 596950
rect 180984 596858 180988 596863
rect 180984 596672 181012 596858
rect 180984 594392 180988 596672
rect 182916 594392 182920 596863
rect 183440 595534 183688 595554
rect 183460 595343 183461 595534
rect 183668 595343 183688 595534
rect 183460 595342 183688 595343
rect 180278 594358 183626 594392
rect 180290 594324 180324 594358
rect 180948 594352 180982 594358
rect 180984 594352 180988 594358
rect 180942 594337 180988 594352
rect 181606 594337 181640 594358
rect 182264 594337 182298 594358
rect 182916 594352 182920 594358
rect 182922 594352 182956 594358
rect 182916 594337 182962 594352
rect 183580 594337 183614 594358
rect 180290 594222 180330 594324
rect 180920 594296 180988 594337
rect 180340 594290 180358 594296
rect 180914 594290 180988 594296
rect 180998 594290 181016 594296
rect 181578 594290 181640 594337
rect 182236 594290 182298 594337
rect 182894 594296 182962 594337
rect 183552 594296 183614 594337
rect 182888 594290 182962 594296
rect 182972 594290 182990 594296
rect 183546 594290 183614 594296
rect 180336 594256 180988 594290
rect 180994 594256 181640 594290
rect 181652 594256 182298 594290
rect 182310 594256 182962 594290
rect 182968 594256 183614 594290
rect 180340 594250 180358 594256
rect 180914 594250 180932 594256
rect 180290 592850 180324 594222
rect 180942 594204 180988 594256
rect 180998 594250 181016 594256
rect 180948 594194 181012 594204
rect 180948 592878 180982 594194
rect 180984 594018 181012 594194
rect 180984 593836 180988 594018
rect 180984 592878 180988 593698
rect 180942 592863 180988 592878
rect 181606 592863 181640 594256
rect 182264 592863 182298 594256
rect 182888 594250 182906 594256
rect 182916 594194 182962 594256
rect 182972 594250 182990 594256
rect 183546 594250 183564 594256
rect 183574 594222 183614 594256
rect 182916 593076 182920 594194
rect 180290 592748 180330 592850
rect 180920 592822 180988 592863
rect 180340 592816 180358 592822
rect 180914 592816 180988 592822
rect 180998 592816 181016 592822
rect 181578 592816 181640 592863
rect 182236 592816 182298 592863
rect 182730 592816 182806 592986
rect 182810 592816 182866 593046
rect 182894 592878 182920 593076
rect 182922 592878 182956 594194
rect 183580 592900 183614 594222
rect 183440 592880 183688 592900
rect 182894 592868 182956 592878
rect 182916 592863 182962 592868
rect 182894 592822 182962 592863
rect 182888 592816 182962 592822
rect 182972 592816 182990 592822
rect 183460 592816 183461 592880
rect 183580 592863 183614 592880
rect 183552 592822 183614 592863
rect 183546 592816 183614 592822
rect 180336 592782 180988 592816
rect 180994 592782 181640 592816
rect 181652 592782 182298 592816
rect 182310 592782 182962 592816
rect 182968 592782 183614 592816
rect 180340 592776 180358 592782
rect 180914 592776 180932 592782
rect 176268 592431 179892 592467
rect 171416 592397 179892 592431
rect 171416 592364 172432 592397
rect 172630 592364 173622 592397
rect 171416 592328 171754 592364
rect 171416 592317 172212 592328
rect 172224 592317 172258 592364
rect 172270 592317 172870 592328
rect 172882 592317 172916 592364
rect 172928 592317 173528 592328
rect 173540 592317 173574 592364
rect 173654 592317 173688 592397
rect 169544 592152 169586 592198
rect 171098 592158 171224 592230
rect 169441 591926 169506 591938
rect 169406 591854 169438 591888
rect 169456 591838 169464 591926
rect 169472 591900 169506 591926
rect 169548 591786 169582 592152
rect 171042 592126 171224 592158
rect 171416 592204 171754 592317
rect 171762 592283 173688 592317
rect 171820 592204 172072 592283
rect 172211 592271 172212 592272
rect 172224 592271 172258 592283
rect 172838 592277 172876 592283
rect 172270 592271 172271 592272
rect 172869 592271 172870 592272
rect 172882 592271 172916 592283
rect 172922 592277 172980 592283
rect 172928 592271 172929 592272
rect 173527 592271 173528 592272
rect 173540 592271 173574 592283
rect 172212 592270 172213 592271
rect 172224 592270 172270 592271
rect 172870 592270 172871 592271
rect 172882 592270 172928 592271
rect 173528 592270 173529 592271
rect 172224 592228 172269 592270
rect 172882 592264 172927 592270
rect 172866 592249 172876 592264
rect 172882 592249 172980 592264
rect 172194 592208 172218 592228
rect 172224 592208 172288 592228
rect 171042 591988 171210 592126
rect 171222 591974 171226 591996
rect 171222 591918 171282 591940
rect 171416 591932 172104 592204
rect 172224 592200 172269 592208
rect 172166 592180 172218 592200
rect 172224 592180 172316 592200
rect 159044 591752 169582 591786
rect 159044 591654 165482 591752
rect 159044 591632 166316 591654
rect 159044 591610 165482 591632
rect 158782 591548 158854 591586
rect 158904 591576 165482 591610
rect 156618 591376 156658 591478
rect 156668 591444 156686 591450
rect 157248 591444 157310 591482
rect 157656 591444 158756 591482
rect 158820 591444 158854 591548
rect 159044 591444 165482 591576
rect 156664 591410 157310 591444
rect 157322 591410 158632 591444
rect 156668 591404 156686 591410
rect 156618 591342 156652 591376
rect 157276 591342 157310 591410
rect 157908 591372 157968 591410
rect 158558 591404 158576 591410
rect 158586 591376 158632 591410
rect 158642 591442 165482 591444
rect 167032 591442 167066 591752
rect 169370 591442 169404 591752
rect 171416 591670 171754 591932
rect 172224 591672 172269 592180
rect 172882 591772 172927 592249
rect 172930 592128 173312 592200
rect 172930 592022 173398 592128
rect 172930 591962 173312 592022
rect 172860 591678 172940 591772
rect 172212 591671 172213 591672
rect 172224 591671 172270 591672
rect 172211 591670 172212 591671
rect 171416 591659 172212 591670
rect 172224 591659 172258 591671
rect 172270 591670 172271 591671
rect 172458 591670 173112 591678
rect 173528 591671 173529 591672
rect 173540 591671 173585 592271
rect 173527 591670 173528 591671
rect 172270 591659 173528 591670
rect 173540 591659 173574 591671
rect 173654 591659 173688 592283
rect 173940 592328 174932 592397
rect 175108 592328 176116 592397
rect 173940 592323 176116 592328
rect 173940 592317 176100 592323
rect 176118 592317 176152 592397
rect 176232 592317 176266 592397
rect 176268 592317 179892 592397
rect 173940 592306 179892 592317
rect 173940 592283 176266 592306
rect 173734 592128 173740 592280
rect 173762 592150 173796 592280
rect 173940 591864 174932 592283
rect 175108 591864 176100 592283
rect 176105 592271 176106 592272
rect 176106 592270 176107 592271
rect 176112 592200 176116 592277
rect 173940 591854 174988 591864
rect 175052 591860 176100 591864
rect 175108 591856 176100 591860
rect 173940 591772 174932 591854
rect 175108 591780 176110 591856
rect 171416 591620 171754 591659
rect 171762 591625 173688 591659
rect 169445 591609 171754 591620
rect 172211 591613 172212 591614
rect 172224 591613 172258 591625
rect 172270 591613 172271 591614
rect 172212 591612 172213 591613
rect 172224 591612 172270 591613
rect 169456 591597 171754 591609
rect 169445 591586 171754 591597
rect 169472 591442 169506 591586
rect 171416 591517 171754 591586
rect 169545 591506 171012 591517
rect 171122 591506 171754 591517
rect 172224 591509 172269 591612
rect 172458 591604 173112 591625
rect 173527 591613 173528 591614
rect 173540 591613 173574 591625
rect 173528 591612 173529 591613
rect 172860 591520 172940 591604
rect 172882 591509 172927 591520
rect 173540 591509 173585 591613
rect 169556 591497 171754 591506
rect 169556 591472 173559 591497
rect 171416 591450 173559 591472
rect 158642 591410 170990 591442
rect 158642 591404 158660 591410
rect 157934 591342 157968 591372
rect 158592 591342 158626 591376
rect 158718 591342 158752 591410
rect 158820 591346 158854 591410
rect 159044 591408 170990 591410
rect 159044 591362 165482 591408
rect 167032 591362 167066 591408
rect 159044 591354 166930 591362
rect 166964 591354 169248 591362
rect 158820 591342 158892 591346
rect 159044 591342 165482 591354
rect 156600 591328 165482 591342
rect 166892 591328 166995 591340
rect 167032 591328 167066 591354
rect 169370 591328 169404 591408
rect 170302 591354 170854 591362
rect 169441 591339 169544 591340
rect 169441 591332 170302 591339
rect 169434 591328 170302 591332
rect 170804 591328 170815 591339
rect 156600 591320 169248 591328
rect 169336 591320 170820 591328
rect 156600 591308 166980 591320
rect 156400 590746 156540 590806
rect 156204 590660 156540 590746
rect 156204 590358 156538 590660
rect 156294 589055 156328 590358
rect 156296 589043 156328 589055
rect 156266 589039 156328 589043
rect 156266 588996 156313 589039
rect 156330 589017 156364 590358
rect 156330 589005 156362 589017
rect 147166 588962 156313 588996
rect 147166 588946 147202 588962
rect 147712 588894 151336 588962
rect 151433 588894 151467 588962
rect 151547 588894 151581 588962
rect 151702 588894 152124 588962
rect 152178 588894 152600 588962
rect 152748 588894 153566 588962
rect 154179 588894 154224 588962
rect 154837 588894 154871 588962
rect 154951 588894 154985 588962
rect 156408 588894 156442 590358
rect 147102 588860 147110 588894
rect 147144 588860 156376 588894
rect 156410 588860 156442 588894
rect 147712 588618 151336 588860
rect 151433 588836 151467 588860
rect 151547 588836 151581 588860
rect 151702 588836 152124 588860
rect 152178 588836 152600 588860
rect 151354 588826 152600 588836
rect 151433 588665 151467 588826
rect 151702 588814 152124 588826
rect 152178 588814 152600 588826
rect 152748 588826 153566 588860
rect 154179 588826 154224 588860
rect 154837 588826 154871 588860
rect 152748 588814 153561 588826
rect 151562 588767 152600 588814
rect 152630 588767 154462 588814
rect 154809 588767 154856 588814
rect 151609 588760 153540 588767
rect 151609 588733 152224 588760
rect 152267 588733 153540 588760
rect 153583 588733 154198 588767
rect 154241 588733 154856 588767
rect 152384 588665 152465 588733
rect 152486 588665 152520 588733
rect 152748 588665 153540 588733
rect 154951 588665 154985 588860
rect 151433 588631 154985 588665
rect 156444 588750 156538 590358
rect 157276 588840 157310 591308
rect 157934 588840 157968 591308
rect 158718 588864 158752 591308
rect 158820 590980 158892 591308
rect 159044 591294 166980 591308
rect 166998 591294 167066 591320
rect 169336 591294 170815 591320
rect 159044 590963 165482 591294
rect 166892 591282 166980 591294
rect 166930 590980 166964 591282
rect 158893 590952 165482 590963
rect 166880 590952 166891 590963
rect 158782 590890 158892 590928
rect 158904 590918 166891 590952
rect 158820 590434 158892 590890
rect 159044 590870 165482 590918
rect 166892 590890 166964 590928
rect 166930 590882 166964 590890
rect 166892 590870 166980 590882
rect 167032 590870 167066 591294
rect 169370 590870 169404 591294
rect 169456 591282 169544 591294
rect 169472 590882 169544 591282
rect 170816 591266 170888 591304
rect 170854 590898 170888 591266
rect 169456 590881 169544 590882
rect 169456 590874 170302 590881
rect 169434 590870 170302 590874
rect 170804 590870 170815 590881
rect 159044 590854 166980 590870
rect 166998 590854 167066 590870
rect 159044 590836 167066 590854
rect 169336 590836 170815 590870
rect 159044 590830 167030 590836
rect 159044 590826 165482 590830
rect 166892 590826 166995 590830
rect 159044 590824 167002 590826
rect 159044 590802 166924 590824
rect 166970 590802 167002 590824
rect 159044 590756 165482 590802
rect 167032 590756 167066 590836
rect 169370 590756 169404 590836
rect 169441 590824 169544 590836
rect 170956 590756 170990 591408
rect 171416 591416 172243 591450
rect 172286 591416 172901 591450
rect 172944 591416 173559 591450
rect 171416 591348 171754 591416
rect 173654 591348 173688 591625
rect 171416 591314 173688 591348
rect 174030 591659 174064 591772
rect 174144 591672 174189 591772
rect 174802 591672 174847 591772
rect 175460 591766 175505 591780
rect 174144 591671 174190 591672
rect 174790 591671 174791 591672
rect 174802 591671 174848 591672
rect 174144 591659 174178 591671
rect 174190 591670 174191 591671
rect 174789 591670 174790 591671
rect 174190 591659 174790 591670
rect 174802 591659 174836 591671
rect 174848 591670 174849 591671
rect 175368 591670 175398 591752
rect 175424 591670 175426 591752
rect 175448 591671 175449 591672
rect 175447 591670 175448 591671
rect 174848 591659 175448 591670
rect 175456 591670 175776 591766
rect 176084 591670 176110 591780
rect 175456 591659 176110 591670
rect 176112 591665 176116 591752
rect 176118 591659 176152 592283
rect 176232 591659 176266 592283
rect 176268 591659 179892 592306
rect 174030 591625 179892 591659
rect 174030 591354 174064 591625
rect 174144 591613 174178 591625
rect 174190 591613 174191 591614
rect 174789 591613 174790 591614
rect 174802 591613 174836 591625
rect 174848 591613 174849 591614
rect 174144 591612 174190 591613
rect 174790 591612 174791 591613
rect 174802 591612 174848 591613
rect 174144 591515 174189 591612
rect 174802 591515 174847 591612
rect 175368 591548 175398 591619
rect 175424 591562 175426 591619
rect 175447 591613 175448 591614
rect 175448 591612 175449 591613
rect 175456 591588 175776 591625
rect 175368 591506 175426 591548
rect 175460 591515 175505 591588
rect 175532 591562 175564 591576
rect 175532 591506 175564 591548
rect 176084 591503 176110 591625
rect 176112 591562 176116 591619
rect 176118 591515 176152 591625
rect 176118 591503 176144 591515
rect 174159 591499 176144 591503
rect 174159 591456 176137 591499
rect 174206 591422 174821 591456
rect 174864 591422 175479 591456
rect 175522 591422 176137 591456
rect 176232 591354 176266 591625
rect 174030 591320 176266 591354
rect 171416 591278 171754 591314
rect 171531 591130 171754 591278
rect 171531 591094 172432 591130
rect 159044 590722 170990 590756
rect 171476 591060 172432 591094
rect 158820 590322 158854 590434
rect 159044 590294 165482 590722
rect 166896 590352 166914 590378
rect 166924 590324 166942 590378
rect 158904 590280 165482 590294
rect 158782 590232 158854 590270
rect 158904 590260 166880 590280
rect 158820 589664 158854 590232
rect 159044 590246 165482 590260
rect 167032 590246 167066 590722
rect 169370 590246 169404 590722
rect 159044 590212 169582 590246
rect 159044 590198 166298 590212
rect 159044 590182 165482 590198
rect 159044 590144 166892 590182
rect 166930 590144 166964 590212
rect 167032 590144 167066 590212
rect 159044 590110 167066 590144
rect 159044 589636 165482 590110
rect 166891 590072 166892 590073
rect 166930 590072 166964 590110
rect 166892 590071 166893 590072
rect 166930 589764 167002 590072
rect 166930 589664 166964 589764
rect 166880 589636 166891 589647
rect 158782 589574 158854 589612
rect 158904 589602 166891 589636
rect 158820 589006 158854 589574
rect 159044 589234 165482 589602
rect 166892 589574 166964 589612
rect 166892 589272 166893 589273
rect 166891 589271 166892 589272
rect 166930 589234 166964 589574
rect 167032 589234 167066 590110
rect 159044 589200 167066 589234
rect 159044 589132 165482 589200
rect 166930 589132 166964 589200
rect 167032 589132 167066 589200
rect 169370 589132 169404 590212
rect 169406 590110 169438 590144
rect 169456 590072 169464 590202
rect 169472 590072 169506 590212
rect 169441 590060 169506 590072
rect 169434 589284 169506 590060
rect 169441 589272 169506 589284
rect 169406 589200 169438 589234
rect 169456 589184 169464 589272
rect 169472 589132 169506 589272
rect 169548 589145 169582 590212
rect 171476 589780 171510 591060
rect 171531 589780 172432 591060
rect 171476 589746 172432 589780
rect 171531 589710 172432 589746
rect 172630 589710 173622 591130
rect 171531 589697 171754 589710
rect 171531 589639 171772 589697
rect 171531 589145 171754 589639
rect 173734 589468 173740 591150
rect 173762 589496 173796 591150
rect 169545 589134 170912 589145
rect 171434 589134 171754 589145
rect 169548 589132 171754 589134
rect 159044 589100 171754 589132
rect 173940 589118 174932 591138
rect 175108 589126 176100 591146
rect 159044 589098 169582 589100
rect 159044 589026 165482 589098
rect 159044 589006 166300 589026
rect 159044 588978 165482 589006
rect 158904 588944 165482 588978
rect 159044 588864 165482 588944
rect 167032 588926 167066 589098
rect 158718 588842 165482 588864
rect 158718 588830 167066 588842
rect 157818 588816 158756 588824
rect 157818 588802 157926 588816
rect 159044 588794 165482 588830
rect 157784 588768 157922 588790
rect 157980 588782 158580 588790
rect 158638 588782 158790 588790
rect 158704 588756 158866 588758
rect 156444 588654 156532 588750
rect 158742 588718 158828 588720
rect 159044 588700 160092 588794
rect 160128 588790 160290 588794
rect 160458 588788 165482 588794
rect 169370 588788 169404 589098
rect 171531 589039 171754 589100
rect 171531 589027 171772 589039
rect 176268 589027 179892 591625
rect 171531 589020 179892 589027
rect 169425 588993 179892 589020
rect 169425 588986 171772 588993
rect 171531 588981 171772 588986
rect 171531 588843 171754 588981
rect 176268 588843 179892 588993
rect 179899 588913 179910 592397
rect 180140 589990 180223 592721
rect 180290 592714 180324 592748
rect 180942 592720 180988 592782
rect 180998 592776 181016 592782
rect 180948 592714 180982 592720
rect 180984 592714 180988 592720
rect 181606 592714 181640 592782
rect 182264 592714 182298 592782
rect 182730 592734 182806 592782
rect 182730 592714 182808 592734
rect 182810 592714 182868 592782
rect 182888 592776 182906 592782
rect 182916 592720 182962 592782
rect 182972 592776 182990 592782
rect 182916 592714 182920 592720
rect 182922 592714 182956 592720
rect 183460 592714 183461 592782
rect 183546 592776 183564 592782
rect 183574 592748 183614 592782
rect 183580 592714 183614 592748
rect 180272 592689 183626 592714
rect 183632 592689 183648 592714
rect 183668 592689 183688 592880
rect 180272 592688 183688 592689
rect 180272 592680 183626 592688
rect 183632 592680 183648 592688
rect 180984 590209 180988 592680
rect 181606 590221 181640 592680
rect 182730 592650 182808 592680
rect 182810 592650 182868 592680
rect 182809 592174 182814 592438
rect 182809 592078 182820 592174
rect 182916 592014 182920 592680
rect 182850 591446 182960 592014
rect 182916 590422 182920 591446
rect 182894 590214 182920 590422
rect 182916 590209 182920 590214
rect 183694 590122 183728 596950
rect 183934 591794 184232 591810
rect 183950 591554 184232 591794
rect 160166 588752 160252 588764
rect 160458 588760 170990 588788
rect 160606 588754 170990 588760
rect 160128 588700 160152 588742
rect 160166 588700 160190 588752
rect 152384 588618 152465 588631
rect 150154 588240 150188 588618
rect 150214 588240 150337 588618
rect 152384 588253 152418 588618
rect 152337 588240 152418 588253
rect 152486 588240 152520 588631
rect 152748 588240 153540 588631
rect 156444 588618 156514 588654
rect 159044 588640 160350 588700
rect 160606 588640 165482 588754
rect 169370 588674 169404 588754
rect 169441 588685 169544 588686
rect 169441 588678 170302 588685
rect 169434 588674 170302 588678
rect 170804 588674 170815 588685
rect 169336 588640 170815 588674
rect 170820 588650 170922 588652
rect 170816 588644 170922 588650
rect 160788 588618 160792 588640
rect 160816 588634 160820 588640
rect 147144 588206 156376 588240
rect 147156 588185 147190 588206
rect 150154 588185 150188 588206
rect 147156 588138 150188 588185
rect 147156 585801 147190 588138
rect 147218 588104 150188 588138
rect 150154 587096 150188 588104
rect 150214 588185 150337 588206
rect 150214 588138 151314 588185
rect 152384 588138 152418 588206
rect 152486 588138 152520 588206
rect 152748 588185 153540 588206
rect 156330 588185 156364 588206
rect 152630 588138 154462 588185
rect 156302 588138 156364 588185
rect 150214 588104 156364 588138
rect 150214 587780 150337 588104
rect 150214 587238 150290 587780
rect 152384 587238 152418 588104
rect 150214 587222 150282 587238
rect 150214 587096 150248 587222
rect 152325 587210 152336 587221
rect 150349 587176 152336 587210
rect 152486 587096 152520 588104
rect 150154 587062 152520 587096
rect 150214 585801 150248 587062
rect 152748 587002 153540 588104
rect 153272 585801 153306 587002
rect 156330 585801 156364 588104
rect 147156 585754 148474 585801
rect 150186 585788 150248 585801
rect 153244 585788 153306 585801
rect 150186 585760 150254 585788
rect 153244 585760 153312 585788
rect 150180 585754 150254 585760
rect 150264 585754 150282 585760
rect 153238 585754 153312 585760
rect 153322 585754 153340 585760
rect 153556 585754 154470 585801
rect 156302 585760 156364 585801
rect 156296 585754 156364 585760
rect 147156 585686 147196 585754
rect 147206 585720 150254 585754
rect 150260 585720 153312 585754
rect 153318 585720 156364 585754
rect 147206 585714 147224 585720
rect 150180 585714 150198 585720
rect 150208 585686 150254 585720
rect 150264 585714 150282 585720
rect 153238 585714 153256 585720
rect 153266 585686 153312 585720
rect 153322 585714 153340 585720
rect 156296 585714 156314 585720
rect 156324 585686 156364 585720
rect 147156 585652 147190 585686
rect 150214 585652 150248 585686
rect 153272 585652 153306 585686
rect 156330 585652 156364 585686
rect 147138 585618 156398 585652
rect 156444 584024 156478 588618
rect 156502 587780 156512 588618
rect 159044 588282 159444 588318
rect 159494 588282 159528 588314
rect 159689 588282 159865 588316
rect 160026 588282 160060 588314
rect 160606 588282 165482 588318
rect 159044 588248 165482 588282
rect 159044 588006 159444 588248
rect 159494 588168 159528 588248
rect 159596 588196 159630 588206
rect 159924 588196 159958 588206
rect 159565 588168 159677 588180
rect 159877 588168 159989 588180
rect 160026 588168 160060 588248
rect 160070 588180 160152 588206
rect 159494 588142 160190 588168
rect 159494 588134 160060 588142
rect 159494 588054 159528 588134
rect 160026 588132 160060 588134
rect 159872 588128 160060 588132
rect 160026 588054 160060 588128
rect 159494 588020 160060 588054
rect 160606 588102 165482 588248
rect 169370 588216 169404 588640
rect 169456 588628 169544 588640
rect 169472 588476 169544 588628
rect 170816 588624 170888 588644
rect 170816 588612 170894 588624
rect 170848 588588 170894 588612
rect 170848 588578 170888 588588
rect 170854 588460 170888 588578
rect 169545 588448 170302 588459
rect 170816 588448 170904 588460
rect 169434 588386 169544 588424
rect 169556 588414 170904 588448
rect 169472 588228 169544 588386
rect 170302 588380 170306 588410
rect 170816 588402 170904 588414
rect 170854 588278 170888 588402
rect 170848 588252 170888 588278
rect 170848 588232 170894 588252
rect 169456 588227 169544 588228
rect 169456 588220 170306 588227
rect 169434 588216 170306 588220
rect 170804 588216 170815 588227
rect 169336 588182 170815 588216
rect 169370 588102 169404 588182
rect 169441 588170 169544 588182
rect 170956 588102 170990 588754
rect 184343 588727 184377 599555
rect 184507 599509 184574 599522
rect 185022 599509 185099 599522
rect 185165 599509 185232 599522
rect 185680 599509 185757 599522
rect 185823 599509 185894 599522
rect 186342 599509 186415 599522
rect 186481 599509 186564 599522
rect 187012 599509 187073 599522
rect 187139 599509 187216 599522
rect 187664 599509 187731 599522
rect 187089 596997 187123 599456
rect 184445 596963 187793 596997
rect 184457 596929 184491 596963
rect 185115 596942 185149 596963
rect 185773 596942 185807 596963
rect 186431 596942 186465 596963
rect 187089 596942 187123 596963
rect 187747 596942 187781 596963
rect 185087 596929 185149 596942
rect 185745 596929 185807 596942
rect 186403 596929 186465 596942
rect 187061 596929 187123 596942
rect 184457 596827 184497 596929
rect 185087 596901 185155 596929
rect 185745 596901 185813 596929
rect 186403 596901 186471 596929
rect 187061 596901 187129 596929
rect 187719 596901 187781 596942
rect 184507 596895 184525 596901
rect 185081 596895 185155 596901
rect 185165 596895 185183 596901
rect 185739 596895 185813 596901
rect 185823 596895 185841 596901
rect 186397 596895 186471 596901
rect 186481 596895 186499 596901
rect 187055 596895 187129 596901
rect 187139 596895 187157 596901
rect 187713 596895 187781 596901
rect 184503 596861 185155 596895
rect 185161 596861 185813 596895
rect 185819 596861 186471 596895
rect 186477 596861 187129 596895
rect 187135 596861 187781 596895
rect 184507 596855 184525 596861
rect 185081 596855 185099 596861
rect 185109 596827 185155 596861
rect 185165 596855 185183 596861
rect 185739 596855 185757 596861
rect 185767 596827 185813 596861
rect 185823 596855 185841 596861
rect 186397 596855 186415 596861
rect 186425 596827 186471 596861
rect 186481 596855 186499 596861
rect 187055 596855 187073 596861
rect 187083 596827 187129 596861
rect 187139 596855 187157 596861
rect 187713 596855 187731 596861
rect 187741 596827 187781 596861
rect 184457 591455 184491 596827
rect 185115 591468 185149 596827
rect 185773 591468 185807 596827
rect 186431 591468 186465 596827
rect 187089 591468 187123 596827
rect 187747 591468 187781 596827
rect 185087 591455 185149 591468
rect 185745 591455 185807 591468
rect 186403 591455 186465 591468
rect 187061 591455 187123 591468
rect 184457 591353 184497 591455
rect 185087 591427 185155 591455
rect 185745 591427 185813 591455
rect 186403 591427 186471 591455
rect 187061 591427 187129 591455
rect 187719 591427 187781 591468
rect 184507 591421 184525 591427
rect 185081 591421 185155 591427
rect 185165 591421 185183 591427
rect 185739 591421 185813 591427
rect 185823 591421 185841 591427
rect 186397 591421 186471 591427
rect 186481 591421 186499 591427
rect 187055 591421 187129 591427
rect 187139 591421 187157 591427
rect 187713 591421 187781 591427
rect 184503 591387 185155 591421
rect 185161 591387 185813 591421
rect 185819 591387 186471 591421
rect 186477 591387 187129 591421
rect 187135 591387 187781 591421
rect 184507 591381 184525 591387
rect 185081 591381 185099 591387
rect 185109 591353 185155 591387
rect 185165 591381 185183 591387
rect 185739 591381 185757 591387
rect 185767 591353 185813 591387
rect 185823 591381 185841 591387
rect 186397 591381 186415 591387
rect 186425 591353 186471 591387
rect 186481 591381 186499 591387
rect 187055 591381 187073 591387
rect 187083 591353 187129 591387
rect 187139 591381 187157 591387
rect 187713 591381 187731 591387
rect 187741 591353 187781 591387
rect 184457 591319 184491 591353
rect 185115 591319 185149 591353
rect 185773 591319 185807 591353
rect 186431 591319 186465 591353
rect 187089 591319 187123 591353
rect 187747 591319 187781 591353
rect 184439 591285 187793 591319
rect 187799 591285 187815 591319
rect 187861 588727 187895 599555
rect 189279 598349 189313 605021
rect 189393 604959 189427 605120
rect 190051 605108 190085 605120
rect 190709 605108 190743 605120
rect 189429 604993 189433 605095
rect 189457 605061 189461 605067
rect 190037 605061 190085 605108
rect 190695 605061 190743 605108
rect 189453 605027 189461 605061
rect 189469 605027 190085 605061
rect 190111 605027 190119 605061
rect 190127 605027 190743 605061
rect 189457 605021 189461 605027
rect 190039 605011 190085 605027
rect 190697 605011 190743 605027
rect 190051 604959 190085 605011
rect 190709 604959 190743 605011
rect 190745 604993 190749 605095
rect 191290 605067 191292 606164
rect 191318 605067 191320 606136
rect 191367 605120 191415 606424
rect 192025 605120 192073 606424
rect 191367 605108 191401 605120
rect 192025 605108 192059 605120
rect 190773 605061 190777 605067
rect 191353 605061 191401 605108
rect 192011 605061 192059 605108
rect 190769 605027 190777 605061
rect 190785 605027 191401 605061
rect 191427 605027 191435 605061
rect 191443 605027 192059 605061
rect 190773 605021 190777 605027
rect 191290 605014 191292 605021
rect 191318 604986 191320 605021
rect 191355 605011 191401 605027
rect 192013 605011 192059 605027
rect 191367 604959 191401 605011
rect 192025 604959 192059 605011
rect 192061 604993 192065 605095
rect 192612 605067 192614 606134
rect 192640 605067 192642 606106
rect 192683 605120 192731 606424
rect 192683 605108 192717 605120
rect 192089 605061 192093 605067
rect 192669 605061 192717 605108
rect 192085 605027 192093 605061
rect 192101 605027 192717 605061
rect 192089 605021 192093 605027
rect 192612 605014 192614 605021
rect 192640 604986 192642 605021
rect 192671 605011 192717 605027
rect 192683 604959 192717 605011
rect 192797 605021 192845 606523
rect 194350 605044 194398 606528
rect 194478 606538 194512 606590
rect 195094 606556 195132 606560
rect 194478 606450 194524 606538
rect 195094 606522 195134 606556
rect 194526 606488 195134 606522
rect 195102 606482 195106 606488
rect 195130 606454 195134 606488
rect 195136 606538 195170 606590
rect 195136 606450 195182 606538
rect 195752 606522 195790 606560
rect 195184 606488 195790 606522
rect 195794 606528 195860 606590
rect 195884 606528 195888 606590
rect 195794 606482 195840 606528
rect 196410 606522 196448 606560
rect 195842 606488 196448 606522
rect 196452 606538 196486 606590
rect 197046 606560 197072 606590
rect 197074 606560 197144 606590
rect 197046 606538 197144 606560
rect 197726 606556 197764 606560
rect 194478 606438 194512 606450
rect 195111 606438 195124 606449
rect 195136 606438 195170 606450
rect 195769 606438 195782 606449
rect 195794 606438 195860 606482
rect 194464 605134 194512 606438
rect 189381 604925 192729 604959
rect 192797 599941 192831 605021
rect 192797 599692 192867 599941
rect 189378 598217 192867 599692
rect 194350 599687 194384 605044
rect 194464 604982 194498 605134
rect 194500 605016 194504 605118
rect 195050 605090 195058 605902
rect 195078 605090 195086 605874
rect 195122 605134 195170 606438
rect 195780 605424 195860 606438
rect 195122 605122 195156 605134
rect 195780 605122 195834 605424
rect 195884 605396 195888 606482
rect 196452 606450 196498 606538
rect 197046 606528 197156 606538
rect 197068 606522 197106 606528
rect 196500 606488 197106 606522
rect 197110 606482 197156 606528
rect 197726 606522 197766 606556
rect 197158 606488 197766 606522
rect 197734 606482 197738 606488
rect 196427 606438 196440 606449
rect 196452 606438 196486 606450
rect 196438 605134 196486 606438
rect 197046 605360 197072 606482
rect 197074 606450 197156 606482
rect 197762 606454 197766 606488
rect 197074 605388 197144 606450
rect 197743 606438 197756 606449
rect 197768 606438 197802 606590
rect 197882 606528 197916 609538
rect 205852 609534 205872 609654
rect 205880 609528 205900 609682
rect 211084 609484 211104 609638
rect 211112 609490 211132 609610
rect 198534 608174 206510 608208
rect 199116 607592 200220 607612
rect 197062 605314 197072 605360
rect 197090 605314 197144 605388
rect 197678 605314 197684 605886
rect 197706 605314 197712 605858
rect 197096 605176 197144 605314
rect 196438 605122 196472 605134
rect 194528 605084 194532 605090
rect 195108 605084 195156 605122
rect 195766 605090 195820 605122
rect 195766 605084 195814 605090
rect 194524 605050 194532 605084
rect 194540 605050 195156 605084
rect 195182 605050 195190 605084
rect 195198 605050 195814 605084
rect 194528 605044 194532 605050
rect 195050 605038 195058 605044
rect 195078 605010 195086 605044
rect 195110 605034 195156 605050
rect 195768 605044 195814 605050
rect 195816 605044 195820 605090
rect 195844 605084 195848 605090
rect 196424 605084 196472 605122
rect 197062 605090 197072 605176
rect 197090 605134 197144 605176
rect 197090 605122 197130 605134
rect 197082 605084 197130 605122
rect 195840 605050 195848 605084
rect 195856 605050 196472 605084
rect 196498 605050 196506 605084
rect 196514 605050 197130 605084
rect 195844 605044 195848 605050
rect 195768 605034 195820 605044
rect 196426 605034 196472 605050
rect 195122 604982 195156 605034
rect 195780 604988 195820 605034
rect 195780 604982 195814 604988
rect 196438 604982 196472 605034
rect 197062 604982 197072 605044
rect 197084 605034 197130 605050
rect 197090 604982 197130 605034
rect 197132 605016 197136 605118
rect 197678 605090 197684 605176
rect 197706 605090 197712 605176
rect 197754 605134 197802 606438
rect 197754 605122 197788 605134
rect 197160 605084 197164 605090
rect 197740 605084 197788 605122
rect 197156 605050 197164 605084
rect 197172 605050 197788 605084
rect 197160 605044 197164 605050
rect 197678 605032 197684 605044
rect 197706 605010 197712 605044
rect 197742 605034 197788 605050
rect 197754 604982 197788 605034
rect 197868 605044 197916 606528
rect 198312 606514 201623 606655
rect 206594 606624 206596 606658
rect 198195 606483 201623 606514
rect 198312 606480 201623 606483
rect 198115 606102 198138 606464
rect 198161 606449 201623 606480
rect 198143 606102 198166 606436
rect 198312 605462 201623 606449
rect 203106 606590 206641 606624
rect 203106 606234 203140 606590
rect 203850 606522 203888 606560
rect 204508 606522 204546 606560
rect 205166 606522 205204 606560
rect 205824 606522 205862 606560
rect 206482 606522 206520 606560
rect 203282 606488 203888 606522
rect 203940 606488 204546 606522
rect 204598 606488 205204 606522
rect 205256 606488 205862 606522
rect 205914 606488 206520 606522
rect 206560 606478 206578 606488
rect 203209 606438 203254 606449
rect 203867 606438 203912 606449
rect 204525 606438 204570 606449
rect 205183 606438 205228 606449
rect 205841 606438 205886 606449
rect 203220 606234 203254 606438
rect 203265 606246 203266 606247
rect 203866 606246 203867 606247
rect 203266 606245 203267 606246
rect 203865 606245 203866 606246
rect 203878 606234 203912 606438
rect 203923 606246 203924 606247
rect 204524 606246 204525 606247
rect 203924 606245 203925 606246
rect 204523 606245 204524 606246
rect 204536 606234 204570 606438
rect 204581 606246 204582 606247
rect 205182 606246 205183 606247
rect 204582 606245 204583 606246
rect 205181 606245 205182 606246
rect 205194 606234 205228 606438
rect 205239 606246 205240 606247
rect 205840 606246 205841 606247
rect 205240 606245 205241 606246
rect 205839 606245 205840 606246
rect 205852 606234 205886 606438
rect 206476 606326 206494 606478
rect 206554 606476 206578 606478
rect 206526 606450 206544 606454
rect 206554 606450 206582 606476
rect 206504 606449 206582 606450
rect 206499 606438 206582 606449
rect 206504 606298 206582 606438
rect 206510 606262 206582 606298
rect 206510 606250 206578 606262
rect 205897 606246 205898 606247
rect 206498 606246 206499 606247
rect 205898 606245 205899 606246
rect 206497 606245 206498 606246
rect 206510 606234 206556 606250
rect 206560 606246 206578 606250
rect 206590 606246 206594 606590
rect 206624 606262 206641 606590
rect 203072 606231 206556 606234
rect 203072 606222 206550 606231
rect 203072 606212 206544 606222
rect 206624 606219 206628 606262
rect 203072 606210 206550 606212
rect 203072 606200 206556 606210
rect 203106 605576 203140 606200
rect 203220 605576 203254 606200
rect 203266 606188 203267 606189
rect 203865 606188 203866 606189
rect 203265 606187 203266 606188
rect 203866 606187 203867 606188
rect 203265 605588 203266 605589
rect 203866 605588 203867 605589
rect 203266 605587 203267 605588
rect 203865 605587 203866 605588
rect 203878 605576 203912 606200
rect 203924 606188 203925 606189
rect 204523 606188 204524 606189
rect 203923 606187 203924 606188
rect 204524 606187 204525 606188
rect 203923 605588 203924 605589
rect 204524 605588 204525 605589
rect 203924 605587 203925 605588
rect 204523 605587 204524 605588
rect 204536 605576 204570 606200
rect 204582 606188 204583 606189
rect 205181 606188 205182 606189
rect 204581 606187 204582 606188
rect 205182 606187 205183 606188
rect 204581 605588 204582 605589
rect 205182 605588 205183 605589
rect 204582 605587 204583 605588
rect 205181 605587 205182 605588
rect 205194 605576 205228 606200
rect 205240 606188 205241 606189
rect 205839 606188 205840 606189
rect 205239 606187 205240 606188
rect 205840 606187 205841 606188
rect 205239 605588 205240 605589
rect 205840 605588 205841 605589
rect 205240 605587 205241 605588
rect 205839 605587 205840 605588
rect 205852 605576 205886 606200
rect 205898 606188 205899 606189
rect 206497 606188 206498 606189
rect 205897 606187 205898 606188
rect 206498 606187 206499 606188
rect 206510 606184 206556 606200
rect 206560 606184 206578 606188
rect 206510 606172 206578 606184
rect 206510 606122 206582 606172
rect 205897 605588 205898 605589
rect 206498 605588 206499 605589
rect 205898 605587 205899 605588
rect 206497 605587 206498 605588
rect 206510 605576 206556 606122
rect 206560 605604 206582 606122
rect 206560 605588 206578 605604
rect 206590 605588 206594 606188
rect 206624 605604 206641 606219
rect 203072 605573 206556 605576
rect 203072 605542 206544 605573
rect 206624 605554 206628 605604
rect 203106 605462 203140 605542
rect 203220 605462 203254 605542
rect 203878 605462 203912 605542
rect 204536 605462 204570 605542
rect 205194 605462 205228 605542
rect 205852 605462 205886 605542
rect 206510 605462 206544 605542
rect 198312 605428 206556 605462
rect 206624 605428 206634 605496
rect 206662 605462 206696 606678
rect 228091 606227 228125 612591
rect 230837 609144 230871 612492
rect 230837 608792 230877 609144
rect 228205 606323 228239 606357
rect 228863 606323 228897 606357
rect 229521 606323 229555 606357
rect 230179 606323 230213 606357
rect 230837 606323 230871 608792
rect 231495 606619 231529 606653
rect 231609 606619 231643 612591
rect 233934 606655 233968 612506
rect 233126 606619 234533 606655
rect 236566 606624 236600 606658
rect 236680 606624 236714 612596
rect 230945 606585 234533 606619
rect 230945 606323 230979 606585
rect 231074 606517 231541 606564
rect 231121 606483 231541 606517
rect 231483 606436 231541 606483
rect 231048 606424 231104 606435
rect 231059 606323 231104 606424
rect 231495 606357 231540 606436
rect 231495 606323 231549 606357
rect 231609 606323 231643 606585
rect 233126 606364 234533 606585
rect 228155 606289 228159 606323
rect 228171 606289 231643 606323
rect 198312 605392 201623 605428
rect 194452 604948 197800 604982
rect 195122 599687 195156 604948
rect 195780 599687 195814 604948
rect 197062 604580 197072 604948
rect 197090 604580 197128 604948
rect 196504 604074 197096 604088
rect 197130 604074 197284 604088
rect 196538 604040 197096 604054
rect 197130 604040 197284 604054
rect 197062 602120 197072 603392
rect 197090 602120 197128 603392
rect 197062 600620 197072 600932
rect 197090 600620 197128 600932
rect 195822 599694 195846 600154
rect 195828 599687 195846 599694
rect 189414 588750 189448 598217
rect 189516 596968 192864 597002
rect 189528 591478 189562 596968
rect 190186 596938 190220 596968
rect 190844 596938 190878 596968
rect 191502 596938 191536 596968
rect 192160 596938 192194 596968
rect 192818 596938 192852 596968
rect 190158 596900 190220 596938
rect 190816 596900 190878 596938
rect 191474 596900 191536 596938
rect 192132 596900 192194 596938
rect 192790 596900 192852 596938
rect 189574 596866 190220 596900
rect 190232 596866 190878 596900
rect 190890 596866 191536 596900
rect 191548 596866 192194 596900
rect 192206 596866 192852 596900
rect 189594 592644 189600 592900
rect 189622 592672 189628 592872
rect 189594 592244 189600 592500
rect 189622 592272 189628 592472
rect 190186 591482 190220 596866
rect 190844 591482 190878 596866
rect 191502 591482 191536 596866
rect 192160 591482 192194 596866
rect 192818 591482 192852 596866
rect 190158 591478 190220 591482
rect 190816 591478 190878 591482
rect 191474 591478 191536 591482
rect 192132 591478 192194 591482
rect 189528 591376 189568 591478
rect 190158 591450 190226 591478
rect 190816 591450 190884 591478
rect 191474 591450 191542 591478
rect 192132 591450 192200 591478
rect 192790 591450 192852 591482
rect 189578 591444 189596 591450
rect 190152 591444 190226 591450
rect 190236 591444 190254 591450
rect 190810 591444 190884 591450
rect 190894 591444 190912 591450
rect 191468 591444 191542 591450
rect 191552 591444 191570 591450
rect 192126 591444 192200 591450
rect 192210 591444 192228 591450
rect 192784 591444 192852 591450
rect 189574 591410 190226 591444
rect 190232 591410 190884 591444
rect 190890 591410 191542 591444
rect 191548 591410 192200 591444
rect 192206 591410 192852 591444
rect 189578 591404 189596 591410
rect 190152 591404 190170 591410
rect 190180 591376 190226 591410
rect 190236 591404 190254 591410
rect 190810 591404 190828 591410
rect 190838 591376 190884 591410
rect 190894 591404 190912 591410
rect 191468 591404 191486 591410
rect 191496 591376 191542 591410
rect 191552 591404 191570 591410
rect 192126 591404 192144 591410
rect 192154 591376 192200 591410
rect 192210 591404 192228 591410
rect 192784 591404 192802 591410
rect 192812 591376 192852 591410
rect 189528 591342 189562 591376
rect 190186 591342 190220 591376
rect 190844 591342 190878 591376
rect 191502 591342 191536 591376
rect 192160 591342 192194 591376
rect 192818 591342 192852 591376
rect 189510 591308 192886 591342
rect 190186 589044 190220 591308
rect 191516 590434 192304 590452
rect 191516 590322 191536 590434
rect 192160 590418 192208 590434
rect 191550 590384 192270 590418
rect 190154 589010 190220 589044
rect 190844 589010 190878 589044
rect 190092 588976 191240 589010
rect 190092 588688 190126 588976
rect 190186 588872 190220 588976
rect 190844 588896 190878 588976
rect 191054 588896 191065 588907
rect 190156 588850 190228 588872
rect 190278 588862 191065 588896
rect 190831 588850 190832 588851
rect 190156 588834 190232 588850
rect 190832 588849 190833 588850
rect 190844 588840 190878 588862
rect 190890 588850 190891 588851
rect 190889 588849 190890 588850
rect 191066 588834 191138 588872
rect 190174 588828 190232 588834
rect 190265 588828 190266 588829
rect 191066 588828 191067 588829
rect 190178 588824 190228 588828
rect 190266 588827 190267 588828
rect 190160 588790 190170 588796
rect 190178 588790 190234 588824
rect 190236 588790 190262 588796
rect 190816 588790 190854 588828
rect 191065 588827 191066 588828
rect 191104 588790 191138 588834
rect 191206 588790 191240 588976
rect 191550 588824 191584 590384
rect 192094 590316 192132 590354
rect 191726 590282 192132 590316
rect 192172 590282 192194 590346
rect 192126 590243 192156 590248
rect 191653 590232 191698 590243
rect 192111 590232 192156 590243
rect 191664 588828 191698 590232
rect 192122 588828 192156 590232
rect 192160 588828 192194 590282
rect 191530 588790 191584 588824
rect 190156 588756 190174 588790
rect 190178 588756 190854 588790
rect 190906 588756 191240 588790
rect 190160 588750 190170 588756
rect 190178 588740 190234 588756
rect 190236 588750 190262 588756
rect 190188 588722 190234 588740
rect 190194 588688 190228 588722
rect 191104 588688 191138 588756
rect 191206 588688 191240 588756
rect 191550 588688 191584 588790
rect 191652 588790 191710 588828
rect 192110 588824 192194 588828
rect 192110 588790 192166 588824
rect 192206 588790 192228 590346
rect 191652 588756 192166 588790
rect 191652 588740 191710 588756
rect 192110 588740 192148 588756
rect 191652 588725 191667 588740
rect 192236 588688 192270 590384
rect 192932 588750 192966 599560
rect 193099 588727 193133 599555
rect 193263 599509 193330 599522
rect 193778 599509 193855 599522
rect 193921 599509 193988 599522
rect 194314 598240 196687 599687
rect 197222 599466 197224 600174
rect 197868 598372 197902 605044
rect 198111 604972 198112 605058
rect 198149 604934 198150 605096
rect 198318 605054 198740 605392
rect 198794 605054 199216 605392
rect 201553 603909 201587 605392
rect 201588 605012 201623 605266
rect 201842 604550 201877 605012
rect 202298 604840 202400 604852
rect 203106 603945 203140 605428
rect 203182 605200 203196 605286
rect 203220 605162 203234 605324
rect 228059 604417 228125 606227
rect 228201 606237 228205 606255
rect 228201 606221 228251 606237
rect 228262 606227 228280 606242
rect 228290 606227 228308 606240
rect 228803 606221 228850 606268
rect 228859 606237 228863 606255
rect 228859 606221 228909 606237
rect 229461 606227 229508 606268
rect 229452 606221 229508 606227
rect 229517 606237 229521 606255
rect 229517 606221 229567 606237
rect 229582 606227 229588 606230
rect 229610 606227 229616 606240
rect 230119 606221 230166 606268
rect 230175 606237 230179 606255
rect 230175 606221 230225 606237
rect 230777 606227 230824 606268
rect 230837 606255 230871 606289
rect 230772 606221 230824 606227
rect 230833 606237 230871 606255
rect 230876 606237 230877 606289
rect 230945 606268 230979 606289
rect 231059 606286 231104 606289
rect 231495 606286 231540 606289
rect 231059 606268 231093 606286
rect 230833 606221 230883 606237
rect 230945 606221 230992 606268
rect 231059 606237 231106 606268
rect 231047 606221 231106 606237
rect 231435 606221 231482 606268
rect 228205 606187 228850 606221
rect 228863 606187 229508 606221
rect 229521 606187 230166 606221
rect 230179 606187 230824 606221
rect 230837 606187 231482 606221
rect 228205 606140 228251 606187
rect 228161 606128 228179 606140
rect 228205 606128 228239 606140
rect 228161 604504 228239 606128
rect 228262 604840 228280 606181
rect 228290 604812 228308 606181
rect 228863 606140 228909 606187
rect 229452 606181 229473 606187
rect 229480 606153 229501 606187
rect 229521 606140 229567 606187
rect 228820 606128 228851 606139
rect 228863 606128 228897 606140
rect 229478 606128 229509 606139
rect 229521 606128 229555 606140
rect 228760 604504 228770 605862
rect 228788 604504 228798 605834
rect 228831 604504 228897 606128
rect 229489 604504 229555 606128
rect 229582 604828 229588 606181
rect 229610 604800 229616 606181
rect 230179 606140 230225 606187
rect 230772 606181 230789 606187
rect 230800 606153 230817 606187
rect 230837 606181 230883 606187
rect 230837 606140 230908 606181
rect 230136 606128 230167 606139
rect 230179 606128 230213 606140
rect 230794 606128 230825 606139
rect 230837 606128 230871 606140
rect 230070 604504 230090 605868
rect 230098 604504 230118 605840
rect 230147 604504 230213 606128
rect 230805 604519 230871 606128
rect 230876 604806 230908 606140
rect 230876 604519 230877 604806
rect 230932 604778 230936 606181
rect 230805 604504 230877 604519
rect 230945 604504 230979 606187
rect 231047 606140 231105 606187
rect 231059 604504 231093 606140
rect 231495 606139 231529 606286
rect 231452 606128 231529 606139
rect 231463 604516 231529 606128
rect 231463 604504 231508 604516
rect 228161 604500 230526 604504
rect 228161 604490 228207 604500
rect 228220 604490 230526 604500
rect 228161 604466 230526 604490
rect 228059 604014 228093 604417
rect 228161 604355 228207 604466
rect 228220 604457 230526 604466
rect 230793 604457 230852 604504
rect 230945 604457 230992 604504
rect 231059 604457 231106 604504
rect 231463 604457 231510 604504
rect 228267 604423 228878 604457
rect 228913 604454 229536 604457
rect 228925 604423 229536 604454
rect 229583 604423 230194 604457
rect 230241 604423 230852 604457
rect 230899 604423 231510 604457
rect 228819 604407 228865 604423
rect 229477 604407 229523 604423
rect 230135 604407 230181 604423
rect 230793 604417 230839 604423
rect 230793 604407 230845 604417
rect 230805 604361 230845 604407
rect 230805 604355 230839 604361
rect 230945 604355 230979 604423
rect 231059 604355 231093 604423
rect 231463 604355 231497 604423
rect 231577 604355 231643 606289
rect 233094 606328 234533 606364
rect 236016 606590 239472 606624
rect 234592 606328 234626 606362
rect 235250 606328 235284 606362
rect 235908 606328 235942 606362
rect 236016 606328 236050 606590
rect 236566 606553 236604 606560
rect 236566 606538 236612 606553
rect 236554 606522 236612 606538
rect 236192 606488 236612 606522
rect 236554 606450 236612 606488
rect 236119 606438 236164 606449
rect 236130 606328 236164 606438
rect 236566 606362 236600 606450
rect 236566 606328 236620 606362
rect 236680 606328 236714 606590
rect 233094 606294 236714 606328
rect 233094 606264 234533 606294
rect 233094 606222 234570 606264
rect 234586 606242 234600 606288
rect 234586 606232 234638 606242
rect 234588 606226 234638 606232
rect 235190 606226 235228 606264
rect 235246 606242 235250 606260
rect 235246 606226 235296 606242
rect 235848 606226 235886 606264
rect 235904 606242 235908 606260
rect 235946 606242 235948 606294
rect 236016 606264 236050 606294
rect 236130 606264 236164 606294
rect 235904 606226 235954 606242
rect 236016 606226 236054 606264
rect 236130 606242 236168 606264
rect 236118 606226 236176 606242
rect 236506 606226 236544 606264
rect 233094 606192 234572 606222
rect 233094 606186 234544 606192
rect 231674 604778 231680 606130
rect 232440 605122 232478 605322
rect 232496 605094 232506 605350
rect 228161 604321 231643 604355
rect 233094 604480 234533 606186
rect 234550 606158 234572 606192
rect 234592 606192 235228 606226
rect 235250 606192 235886 606226
rect 235908 606192 236544 606226
rect 234550 606153 234564 606158
rect 234592 606154 234638 606192
rect 235250 606154 235296 606192
rect 235908 606186 235954 606192
rect 236016 606186 236050 606192
rect 235908 606154 235980 606186
rect 234549 606142 234580 606153
rect 234592 606142 234626 606154
rect 235207 606142 235238 606153
rect 235250 606142 235284 606154
rect 235865 606142 235896 606153
rect 235908 606142 235942 606154
rect 234550 604820 234626 606142
rect 234554 604530 234626 604820
rect 234554 604518 234594 604530
rect 234548 604480 234598 604518
rect 235150 604486 235166 605418
rect 235178 604486 235194 605418
rect 235218 604530 235284 606142
rect 235294 604728 235314 605418
rect 235876 604542 235942 606142
rect 235946 604784 235980 606154
rect 235946 604542 235948 604784
rect 236002 604728 236050 606186
rect 236118 606154 236176 606192
rect 235218 604518 235252 604530
rect 235876 604518 235948 604542
rect 236016 604518 236050 604728
rect 236130 604518 236164 606154
rect 236566 606153 236600 606294
rect 236523 606142 236600 606153
rect 236534 604530 236600 606142
rect 235206 604480 235256 604518
rect 235864 604486 235916 604518
rect 235864 604480 235914 604486
rect 236016 604480 236054 604518
rect 236130 604480 236168 604518
rect 236534 604514 236579 604530
rect 236534 604480 236572 604514
rect 233094 604446 234598 604480
rect 234654 604446 235256 604480
rect 235312 604446 235914 604480
rect 235970 604446 236572 604480
rect 233094 604378 234533 604446
rect 234548 604430 234594 604446
rect 235206 604430 235252 604446
rect 235864 604440 235910 604446
rect 235864 604430 235916 604440
rect 235876 604384 235916 604430
rect 235876 604378 235910 604384
rect 236016 604378 236050 604446
rect 236130 604382 236164 604446
rect 236534 604382 236568 604446
rect 236130 604378 236175 604382
rect 236534 604378 236579 604382
rect 236648 604378 236714 606294
rect 236750 605874 236766 605876
rect 236744 604770 236766 605874
rect 236788 605778 236822 606438
rect 236788 605696 236888 605778
rect 236750 604486 236766 604686
rect 233094 604344 236714 604378
rect 228173 604014 228207 604048
rect 228831 604014 228865 604048
rect 229489 604014 229523 604048
rect 230147 604014 230181 604048
rect 226874 603980 230330 604014
rect 203070 603909 206694 603945
rect 198353 603875 206694 603909
rect 198353 600391 198387 603875
rect 198807 603874 198841 603875
rect 198807 603801 198847 603874
rect 198866 603801 198875 603846
rect 198807 603795 198841 603801
rect 199465 603795 199499 603875
rect 200123 603795 200157 603875
rect 200781 603795 200815 603875
rect 201439 603795 201473 603875
rect 201553 603795 201587 603875
rect 198408 603733 198489 603780
rect 198548 603761 201587 603795
rect 198807 603755 198841 603761
rect 198794 603749 198795 603750
rect 198795 603748 198796 603749
rect 198455 603165 198489 603733
rect 198807 603690 198847 603755
rect 198853 603749 198854 603750
rect 198852 603748 198853 603749
rect 198866 603718 198875 603755
rect 199452 603749 199453 603750
rect 199453 603748 199454 603749
rect 198795 603149 198796 603150
rect 198794 603148 198795 603149
rect 198807 603137 198841 603690
rect 198852 603149 198853 603150
rect 199453 603149 199454 603150
rect 198853 603148 198854 603149
rect 199452 603148 199453 603149
rect 199465 603137 199499 603761
rect 199511 603749 199512 603750
rect 200110 603749 200111 603750
rect 199510 603748 199511 603749
rect 200111 603748 200112 603749
rect 199510 603149 199511 603150
rect 200111 603149 200112 603150
rect 199511 603148 199512 603149
rect 200110 603148 200111 603149
rect 200123 603137 200157 603761
rect 200169 603749 200170 603750
rect 200768 603749 200769 603750
rect 200168 603748 200169 603749
rect 200769 603748 200770 603749
rect 200168 603149 200169 603150
rect 200769 603149 200770 603150
rect 200169 603148 200170 603149
rect 200768 603148 200769 603149
rect 200781 603137 200815 603761
rect 200827 603749 200828 603750
rect 201426 603749 201427 603750
rect 200826 603748 200827 603749
rect 201427 603748 201428 603749
rect 200826 603149 200827 603150
rect 201427 603149 201428 603150
rect 200827 603148 200828 603149
rect 201426 603148 201427 603149
rect 201439 603137 201473 603761
rect 201553 603137 201587 603761
rect 203070 603137 206712 603875
rect 219912 603850 219916 603855
rect 219842 603822 219888 603827
rect 219842 603815 219910 603822
rect 219848 603812 219910 603815
rect 198408 603075 198489 603122
rect 198548 603103 206712 603137
rect 198794 603091 198795 603092
rect 198795 603090 198796 603091
rect 198455 602507 198489 603075
rect 198795 602491 198796 602492
rect 198794 602490 198795 602491
rect 198807 602479 198841 603103
rect 198853 603091 198854 603092
rect 199452 603091 199453 603092
rect 198852 603090 198853 603091
rect 199453 603090 199454 603091
rect 199465 602494 199499 603103
rect 199511 603091 199512 603092
rect 200110 603091 200111 603092
rect 199510 603090 199511 603091
rect 200111 603090 200112 603091
rect 199690 602494 199902 602626
rect 198852 602491 198853 602492
rect 198853 602490 198854 602491
rect 199380 602479 199902 602494
rect 200111 602491 200112 602492
rect 200110 602490 200111 602491
rect 200123 602479 200157 603103
rect 200169 603091 200170 603092
rect 200768 603091 200769 603092
rect 200168 603090 200169 603091
rect 200769 603090 200770 603091
rect 200168 602491 200169 602492
rect 200769 602491 200770 602492
rect 200169 602490 200170 602491
rect 200768 602490 200769 602491
rect 200781 602479 200815 603103
rect 200827 603091 200828 603092
rect 201426 603091 201427 603092
rect 200826 603090 200827 603091
rect 201427 603090 201428 603091
rect 200826 602491 200827 602492
rect 201427 602491 201428 602492
rect 200827 602490 200828 602491
rect 201426 602490 201427 602491
rect 201439 602479 201473 603103
rect 201553 602479 201587 603103
rect 202264 603060 202654 603094
rect 201618 602578 201874 602584
rect 202264 602562 202298 603060
rect 202478 602992 202525 603039
rect 202440 602958 202525 602992
rect 202367 602899 202412 602910
rect 202495 602899 202540 602910
rect 202378 602723 202412 602899
rect 202506 602723 202540 602899
rect 202478 602664 202525 602711
rect 202440 602630 202525 602664
rect 202620 602562 202654 603060
rect 202774 602578 203030 602596
rect 201646 602550 201846 602556
rect 202264 602528 202654 602562
rect 202802 602550 203002 602568
rect 198408 602417 198489 602464
rect 198548 602445 201587 602479
rect 198794 602433 198795 602434
rect 198795 602432 198796 602433
rect 198455 601849 198489 602417
rect 198795 601833 198796 601834
rect 198794 601832 198795 601833
rect 198807 601821 198841 602445
rect 198853 602433 198854 602434
rect 198852 602432 198853 602433
rect 199380 602424 199902 602445
rect 200110 602433 200111 602434
rect 200111 602432 200112 602433
rect 198847 602396 198924 602412
rect 199372 602396 199459 602412
rect 198852 601833 198853 601834
rect 199453 601833 199454 601834
rect 198853 601832 198854 601833
rect 199452 601832 199453 601833
rect 199465 601821 199499 602424
rect 199505 602396 199586 602412
rect 199690 602178 199902 602424
rect 200034 602396 200117 602412
rect 199510 601833 199511 601834
rect 200111 601833 200112 601834
rect 199511 601832 199512 601833
rect 200110 601832 200111 601833
rect 200123 601821 200157 602445
rect 200169 602433 200170 602434
rect 200768 602433 200769 602434
rect 200168 602432 200169 602433
rect 200769 602432 200770 602433
rect 200163 602396 200188 602412
rect 200168 601833 200169 601834
rect 200769 601833 200770 601834
rect 200169 601832 200170 601833
rect 200768 601832 200769 601833
rect 200781 601821 200815 602445
rect 200827 602433 200828 602434
rect 201426 602433 201427 602434
rect 200826 602432 200827 602433
rect 201427 602432 201428 602433
rect 200826 601833 200827 601834
rect 201427 601833 201428 601834
rect 200827 601832 200828 601833
rect 201426 601832 201427 601833
rect 201439 601821 201473 602445
rect 201553 601821 201587 602445
rect 201846 602364 202106 602384
rect 201846 602336 202106 602356
rect 202250 601858 202672 602478
rect 202802 602368 203002 602384
rect 202774 602340 203030 602356
rect 203070 601821 206712 603103
rect 217690 602401 218126 602424
rect 217724 602367 218092 602390
rect 218597 602302 218631 603769
rect 219856 603630 219910 603812
rect 219856 603342 219888 603630
rect 219848 603339 219888 603342
rect 219842 603327 219888 603339
rect 219912 603602 219938 603850
rect 221158 603824 221204 603827
rect 221140 603815 221204 603824
rect 227586 603826 227590 603831
rect 221140 603812 221198 603815
rect 221140 603638 221156 603812
rect 227586 603640 227614 603826
rect 219912 603299 219916 603602
rect 221158 603339 221198 603342
rect 221158 603327 221204 603339
rect 219910 603246 220478 603280
rect 222682 602980 222906 603000
rect 224874 602984 225094 603004
rect 222702 602828 222703 602980
rect 222886 602828 222906 602980
rect 224894 602828 224895 602984
rect 225074 602828 225094 602984
rect 227586 602788 227590 603640
rect 218054 602268 220194 602302
rect 211864 601864 211920 601866
rect 198408 601759 198489 601806
rect 198548 601787 206712 601821
rect 198794 601775 198795 601776
rect 198795 601774 198796 601775
rect 198455 601191 198489 601759
rect 198795 601175 198796 601176
rect 198794 601174 198795 601175
rect 198807 601163 198841 601787
rect 198853 601775 198854 601776
rect 199452 601775 199453 601776
rect 198852 601774 198853 601775
rect 199453 601774 199454 601775
rect 198852 601175 198853 601176
rect 199453 601175 199454 601176
rect 198853 601174 198854 601175
rect 199452 601174 199453 601175
rect 199465 601163 199499 601787
rect 199511 601775 199512 601776
rect 200110 601775 200111 601776
rect 199510 601774 199511 601775
rect 200111 601774 200112 601775
rect 199510 601175 199511 601176
rect 200111 601175 200112 601176
rect 199511 601174 199512 601175
rect 200110 601174 200111 601175
rect 200123 601163 200157 601787
rect 200169 601775 200170 601776
rect 200768 601775 200769 601776
rect 200168 601774 200169 601775
rect 200769 601774 200770 601775
rect 200168 601175 200169 601176
rect 200769 601175 200770 601176
rect 200169 601174 200170 601175
rect 200768 601174 200769 601175
rect 200781 601163 200815 601787
rect 200827 601775 200828 601776
rect 201426 601775 201427 601776
rect 200826 601774 200827 601775
rect 201427 601774 201428 601775
rect 200826 601175 200827 601176
rect 201427 601175 201428 601176
rect 200827 601174 200828 601175
rect 201426 601174 201427 601175
rect 201439 601163 201473 601787
rect 201553 601163 201587 601787
rect 202814 601716 202856 601722
rect 202994 601716 203022 601722
rect 202786 601688 202856 601694
rect 202994 601688 203050 601694
rect 203070 601163 206712 601787
rect 218054 601777 218088 602268
rect 218495 602200 218529 602268
rect 218597 602200 218631 602268
rect 218230 602166 218631 602200
rect 218447 602119 218448 602120
rect 218448 602118 218449 602119
rect 218157 602107 218202 602118
rect 218168 601777 218202 602107
rect 218495 601805 218529 602166
rect 218213 601789 218214 601790
rect 218214 601788 218215 601789
rect 218436 601777 218447 601788
rect 218020 601743 218447 601777
rect 211864 601702 211920 601706
rect 211864 601646 211920 601650
rect 198408 601101 198489 601148
rect 198548 601129 206712 601163
rect 198794 601117 198795 601118
rect 198795 601116 198796 601117
rect 198455 600533 198489 601101
rect 198795 600517 198796 600518
rect 198794 600516 198795 600517
rect 198807 600505 198841 601129
rect 198853 601117 198854 601118
rect 199452 601117 199453 601118
rect 198852 601116 198853 601117
rect 199453 601116 199454 601117
rect 198852 600517 198853 600518
rect 199453 600517 199454 600518
rect 198853 600516 198854 600517
rect 199452 600516 199453 600517
rect 199465 600505 199499 601129
rect 199511 601117 199512 601118
rect 200110 601117 200111 601118
rect 199510 601116 199511 601117
rect 200111 601116 200112 601117
rect 199510 600517 199511 600518
rect 200111 600517 200112 600518
rect 199511 600516 199512 600517
rect 200110 600516 200111 600517
rect 200123 600505 200157 601129
rect 200169 601117 200170 601118
rect 200768 601117 200769 601118
rect 200168 601116 200169 601117
rect 200769 601116 200770 601117
rect 200168 600517 200169 600518
rect 200769 600517 200770 600518
rect 200169 600516 200170 600517
rect 200768 600516 200769 600517
rect 200781 600505 200815 601129
rect 200827 601117 200828 601118
rect 201426 601117 201427 601118
rect 200826 601116 200827 601117
rect 201427 601116 201428 601117
rect 200826 600517 200827 600518
rect 201427 600517 201428 600518
rect 200827 600516 200828 600517
rect 201426 600516 201427 600517
rect 201439 600505 201473 601129
rect 201553 600505 201587 601129
rect 202252 601123 202508 601129
rect 202280 601095 202480 601114
rect 198548 600471 201587 600505
rect 198807 600391 198841 600471
rect 199465 600391 199499 600471
rect 200123 600391 200157 600471
rect 200781 600391 200815 600471
rect 201439 600391 201473 600471
rect 201553 600391 201587 600471
rect 203070 600391 206712 601129
rect 218054 601119 218088 601743
rect 218168 601131 218202 601743
rect 218214 601731 218215 601732
rect 218213 601730 218214 601731
rect 218448 601715 218529 601762
rect 218213 601131 218214 601132
rect 218214 601130 218215 601131
rect 218232 601130 218234 601153
rect 218495 601147 218529 601715
rect 218232 601119 218262 601125
rect 218436 601119 218447 601130
rect 218020 601085 218122 601119
rect 218130 601106 218448 601119
rect 218130 601093 218452 601106
rect 218180 601085 218452 601093
rect 218054 600970 218088 601085
rect 218190 601079 218448 601085
rect 218214 601073 218448 601079
rect 218218 601072 218270 601073
rect 218597 601072 218631 602166
rect 221372 601910 221396 602120
rect 219526 601394 219550 601402
rect 219526 601142 219552 601394
rect 219526 601130 219550 601142
rect 218214 601051 218631 601072
rect 218230 601038 218631 601051
rect 218495 600970 218529 601038
rect 218597 600970 218631 601038
rect 198353 600357 206694 600391
rect 201553 600042 201587 600357
rect 203070 600321 206694 600357
rect 198312 600006 201623 600042
rect 203106 600006 203140 600321
rect 205224 600056 205228 600218
rect 205262 600094 205266 600180
rect 198312 599972 206556 600006
rect 206624 599972 206634 600040
rect 198210 599692 198224 599830
rect 198312 599692 201623 599972
rect 203106 599892 203140 599972
rect 203220 599892 203254 599972
rect 203266 599892 203866 599903
rect 203878 599892 203912 599972
rect 203924 599892 204524 599903
rect 204536 599892 204570 599972
rect 204582 599892 205182 599903
rect 205194 599892 205228 599972
rect 205240 599892 205840 599903
rect 205852 599892 205886 599972
rect 205898 599892 206498 599903
rect 206510 599892 206544 599972
rect 206628 599910 206658 599944
rect 203072 599870 206544 599892
rect 203072 599868 206550 599870
rect 203072 599858 206556 599868
rect 198134 599656 201623 599692
rect 198134 599622 201722 599656
rect 198134 599234 201623 599622
rect 201688 599234 201722 599622
rect 202392 599488 202840 599650
rect 202316 599438 202840 599488
rect 202316 599334 202470 599438
rect 203106 599234 203140 599858
rect 203220 599846 203254 599858
rect 203266 599846 203267 599847
rect 203865 599846 203866 599847
rect 203878 599846 203912 599858
rect 203924 599846 203925 599847
rect 204523 599846 204524 599847
rect 204536 599846 204570 599858
rect 204582 599846 204583 599847
rect 205181 599846 205182 599847
rect 205194 599846 205228 599858
rect 205240 599846 205241 599847
rect 205839 599846 205840 599847
rect 205852 599846 205886 599858
rect 205898 599846 205899 599847
rect 206497 599846 206498 599847
rect 203220 599845 203266 599846
rect 203866 599845 203867 599846
rect 203878 599845 203924 599846
rect 204524 599845 204525 599846
rect 204536 599845 204582 599846
rect 205182 599845 205183 599846
rect 205194 599845 205240 599846
rect 205840 599845 205841 599846
rect 205852 599845 205898 599846
rect 206498 599845 206499 599846
rect 203220 599687 203265 599845
rect 203878 599687 203923 599845
rect 204536 599687 204581 599845
rect 205194 599687 205239 599845
rect 205852 599687 205897 599845
rect 206510 599842 206556 599858
rect 206510 599830 206578 599842
rect 206510 599774 206582 599830
rect 206510 599687 206556 599774
rect 206560 599687 206582 599774
rect 206624 599687 206641 599877
rect 206662 599687 206696 599972
rect 203211 599234 206732 599687
rect 206788 599654 206835 599687
rect 198134 599200 201722 599234
rect 203072 599200 206732 599234
rect 198134 598576 201623 599200
rect 201688 598576 201722 599200
rect 203106 598576 203140 599200
rect 203211 598576 206732 599200
rect 198134 598542 201722 598576
rect 203072 598542 206732 598576
rect 195187 596997 195221 598240
rect 195845 596997 195879 598240
rect 193201 596963 196549 596997
rect 193213 591468 193247 596963
rect 193871 596942 193905 596963
rect 194529 596942 194563 596963
rect 195187 596942 195221 596963
rect 195845 596942 195879 596963
rect 196503 596942 196537 596963
rect 193843 596895 193905 596942
rect 194501 596895 194563 596942
rect 195159 596895 195221 596942
rect 195817 596895 195879 596942
rect 196475 596895 196537 596942
rect 193259 596861 193905 596895
rect 193917 596861 194563 596895
rect 194575 596861 195221 596895
rect 195233 596861 195879 596895
rect 195891 596861 196537 596895
rect 193871 592650 193905 596861
rect 193386 592616 193776 592650
rect 193386 592118 193420 592616
rect 193600 592548 193647 592595
rect 193562 592514 193647 592548
rect 193489 592455 193534 592466
rect 193617 592455 193662 592466
rect 193500 592279 193534 592455
rect 193628 592279 193662 592455
rect 193600 592220 193647 592267
rect 193562 592186 193647 592220
rect 193742 592118 193776 592616
rect 193386 592084 193776 592118
rect 193862 592616 194252 592650
rect 193862 592118 193905 592616
rect 194076 592548 194123 592595
rect 194038 592514 194123 592548
rect 193965 592455 194010 592466
rect 194093 592455 194138 592466
rect 193976 592279 194010 592455
rect 194104 592279 194138 592455
rect 194076 592220 194123 592267
rect 194038 592186 194123 592220
rect 194218 592118 194252 592616
rect 193862 592084 194252 592118
rect 193871 592034 193905 592084
rect 193368 591468 193790 592034
rect 193844 591468 194266 592034
rect 194529 591468 194563 596861
rect 195187 591468 195221 596861
rect 195752 591714 195768 593228
rect 195845 591468 195879 596861
rect 196503 591468 196537 596861
rect 193213 591421 194266 591468
rect 194501 591455 194563 591468
rect 195159 591455 195221 591468
rect 194501 591427 194569 591455
rect 195159 591427 195227 591455
rect 195817 591427 195879 591468
rect 194495 591421 194569 591427
rect 194579 591421 194597 591427
rect 195153 591421 195227 591427
rect 195237 591421 195255 591427
rect 195783 591421 195879 591427
rect 196475 591421 196537 591468
rect 193213 591353 193253 591421
rect 193263 591414 194569 591421
rect 193263 591387 193911 591414
rect 193263 591381 193281 591387
rect 193837 591381 193855 591387
rect 193865 591353 193911 591387
rect 193921 591387 194569 591414
rect 194575 591387 195227 591421
rect 195233 591387 195879 591421
rect 195891 591387 196537 591421
rect 196538 591402 196571 595080
rect 193921 591381 193939 591387
rect 194495 591381 194513 591387
rect 194523 591353 194569 591387
rect 194579 591381 194597 591387
rect 195153 591381 195171 591387
rect 195181 591353 195227 591387
rect 195237 591381 195255 591387
rect 195783 591381 195829 591387
rect 195839 591353 195879 591387
rect 193213 591319 193247 591353
rect 193871 591319 193905 591353
rect 194529 591319 194563 591353
rect 195187 591319 195221 591353
rect 195845 591319 195879 591353
rect 196503 591319 196537 591387
rect 193195 591285 196549 591319
rect 196555 591285 196571 591319
rect 193386 589962 193776 589996
rect 193386 589464 193420 589962
rect 193600 589894 193647 589941
rect 193562 589860 193647 589894
rect 193489 589801 193534 589812
rect 193617 589801 193662 589812
rect 193500 589625 193534 589801
rect 193628 589625 193662 589801
rect 193600 589566 193647 589613
rect 193562 589532 193647 589566
rect 193742 589464 193776 589962
rect 193386 589430 193776 589464
rect 193862 589962 194252 589996
rect 193862 589934 193896 589962
rect 193862 589526 193930 589934
rect 194076 589894 194123 589941
rect 194038 589860 194123 589894
rect 193965 589801 194010 589812
rect 194093 589801 194138 589812
rect 193976 589625 194010 589801
rect 194104 589625 194138 589801
rect 194076 589566 194123 589613
rect 194038 589532 194123 589566
rect 193862 589464 193896 589526
rect 194218 589464 194252 589962
rect 194488 589612 194492 589752
rect 193862 589430 194252 589464
rect 193368 588767 193790 589380
rect 193275 588733 193843 588767
rect 193844 588760 194266 589380
rect 195872 589116 195916 589752
rect 195872 588829 195885 589116
rect 195928 589088 195944 589752
rect 195845 588826 195885 588829
rect 195839 588814 195885 588826
rect 196617 588727 196651 598240
rect 198134 598217 201623 598542
rect 198170 591380 198204 598217
rect 198314 597002 198318 598217
rect 198348 597002 198382 598217
rect 198450 597946 198484 598217
rect 198930 597930 198931 597931
rect 198929 597929 198930 597930
rect 198942 597918 198976 598217
rect 198987 597930 198988 597931
rect 199588 597930 199589 597931
rect 198988 597929 198989 597930
rect 199587 597929 199588 597930
rect 199600 597918 199634 598217
rect 199645 597930 199646 597931
rect 200246 597930 200247 597931
rect 199646 597929 199647 597930
rect 200245 597929 200246 597930
rect 200258 597918 200292 598217
rect 200303 597930 200304 597931
rect 200904 597930 200905 597931
rect 200304 597929 200305 597930
rect 200903 597929 200904 597930
rect 200916 597918 200950 598217
rect 200961 597930 200962 597931
rect 201562 597930 201563 597931
rect 200962 597929 200963 597930
rect 201561 597929 201562 597930
rect 201574 597918 201608 598217
rect 201688 597918 201722 598542
rect 203106 598310 203140 598542
rect 203211 598310 206732 598542
rect 203106 598276 206732 598310
rect 198412 597856 198484 597894
rect 198534 597884 201722 597918
rect 198929 597872 198930 597873
rect 198930 597871 198931 597872
rect 198450 597288 198484 597856
rect 198930 597272 198931 597273
rect 198929 597271 198930 597272
rect 198942 597260 198976 597884
rect 198988 597872 198989 597873
rect 199587 597872 199588 597873
rect 198987 597871 198988 597872
rect 199588 597871 199589 597872
rect 198987 597272 198988 597273
rect 199588 597272 199589 597273
rect 198988 597271 198989 597272
rect 199587 597271 199588 597272
rect 199600 597260 199634 597884
rect 199646 597872 199647 597873
rect 200245 597872 200246 597873
rect 199645 597871 199646 597872
rect 200246 597871 200247 597872
rect 199645 597272 199646 597273
rect 200246 597272 200247 597273
rect 199646 597271 199647 597272
rect 200245 597271 200246 597272
rect 200258 597260 200292 597884
rect 200304 597872 200305 597873
rect 200903 597872 200904 597873
rect 200303 597871 200304 597872
rect 200904 597871 200905 597872
rect 200303 597272 200304 597273
rect 200904 597272 200905 597273
rect 200304 597271 200305 597272
rect 200903 597271 200904 597272
rect 200916 597260 200950 597884
rect 200962 597872 200963 597873
rect 201561 597872 201562 597873
rect 200961 597871 200962 597872
rect 201562 597871 201563 597872
rect 200961 597272 200962 597273
rect 201562 597272 201563 597273
rect 200962 597271 200963 597272
rect 201561 597271 201562 597272
rect 201574 597260 201608 597884
rect 201688 597260 201722 597884
rect 198412 597198 198484 597236
rect 198534 597226 201722 597260
rect 198929 597214 198930 597215
rect 198930 597213 198931 597214
rect 198450 597002 198484 597198
rect 198942 597002 198976 597226
rect 198988 597214 198989 597215
rect 199587 597214 199588 597215
rect 198987 597213 198988 597214
rect 199588 597213 199589 597214
rect 199600 597002 199634 597226
rect 199646 597214 199647 597215
rect 200245 597214 200246 597215
rect 199645 597213 199646 597214
rect 200246 597213 200247 597214
rect 200258 597002 200292 597226
rect 200304 597214 200305 597215
rect 200903 597214 200904 597215
rect 200303 597213 200304 597214
rect 200904 597213 200905 597214
rect 200916 597002 200950 597226
rect 200962 597214 200963 597215
rect 201561 597214 201562 597215
rect 200961 597213 200962 597214
rect 201562 597213 201563 597214
rect 201574 597002 201608 597226
rect 201688 597002 201722 597226
rect 198272 596968 201722 597002
rect 198284 594971 198318 596968
rect 198348 596938 198382 596968
rect 198348 596900 198386 596938
rect 198450 596900 198484 596968
rect 198942 596938 198976 596968
rect 199600 596938 199634 596968
rect 200258 596938 200292 596968
rect 200916 596938 200950 596968
rect 201574 596938 201608 596968
rect 198914 596900 198976 596938
rect 199572 596900 199634 596938
rect 200230 596900 200292 596938
rect 200888 596900 200950 596938
rect 201546 596900 201608 596938
rect 198330 596866 198976 596900
rect 198988 596866 199634 596900
rect 199646 596866 200292 596900
rect 200304 596866 200950 596900
rect 200962 596866 201608 596900
rect 198348 596488 198382 596866
rect 198450 596630 198484 596866
rect 198930 596614 198931 596615
rect 198929 596613 198930 596614
rect 198942 596602 198976 596866
rect 198987 596614 198988 596615
rect 199588 596614 199589 596615
rect 198988 596613 198989 596614
rect 199587 596613 199588 596614
rect 199600 596602 199634 596866
rect 199645 596614 199646 596615
rect 200246 596614 200247 596615
rect 199646 596613 199647 596614
rect 200245 596613 200246 596614
rect 200258 596602 200292 596866
rect 200303 596614 200304 596615
rect 200904 596614 200905 596615
rect 200304 596613 200305 596614
rect 200903 596613 200904 596614
rect 200916 596602 200950 596866
rect 200961 596614 200962 596615
rect 201562 596614 201563 596615
rect 200962 596613 200963 596614
rect 201561 596613 201562 596614
rect 201574 596602 201608 596866
rect 201688 596602 201722 596968
rect 198534 596568 201722 596602
rect 198942 596488 198976 596568
rect 199600 596488 199634 596568
rect 200258 596488 200292 596568
rect 200916 596488 200950 596568
rect 201574 596488 201608 596568
rect 201688 596488 201722 596568
rect 203211 596488 206732 598276
rect 198348 596454 206732 596488
rect 201660 596172 201662 596202
rect 201688 594971 201722 596454
rect 203211 596418 206732 596454
rect 198284 594935 201758 594971
rect 203247 594935 203281 596418
rect 204002 595802 204053 595986
rect 203898 595684 204053 595802
rect 204002 595530 204053 595684
rect 206651 594935 206657 594969
rect 198284 594901 206697 594935
rect 198284 591524 201758 594901
rect 203247 594821 203281 594901
rect 203361 594821 203395 594901
rect 204019 594821 204053 594901
rect 204677 594821 204711 594901
rect 205335 594821 205369 594901
rect 205993 594821 206027 594901
rect 206685 594873 206697 594901
rect 206651 594839 206697 594873
rect 206524 594821 206535 594832
rect 203247 594787 206535 594821
rect 203247 594163 203281 594787
rect 203361 594163 203395 594787
rect 203407 594775 203408 594776
rect 204006 594775 204007 594776
rect 203406 594774 203407 594775
rect 204007 594774 204008 594775
rect 203406 594175 203407 594176
rect 204007 594175 204008 594176
rect 203407 594174 203408 594175
rect 204006 594174 204007 594175
rect 204019 594163 204053 594787
rect 204065 594775 204066 594776
rect 204664 594775 204665 594776
rect 204064 594774 204065 594775
rect 204665 594774 204666 594775
rect 204064 594175 204065 594176
rect 204665 594175 204666 594176
rect 204065 594174 204066 594175
rect 204664 594174 204665 594175
rect 204677 594163 204711 594787
rect 204723 594775 204724 594776
rect 205322 594775 205323 594776
rect 204722 594774 204723 594775
rect 205323 594774 205324 594775
rect 204722 594175 204723 594176
rect 205323 594175 205324 594176
rect 204723 594174 204724 594175
rect 205322 594174 205323 594175
rect 205335 594163 205369 594787
rect 205381 594775 205382 594776
rect 205980 594775 205981 594776
rect 205380 594774 205381 594775
rect 205981 594774 205982 594775
rect 205380 594175 205381 594176
rect 205981 594175 205982 594176
rect 205381 594174 205382 594175
rect 205980 594174 205981 594175
rect 205993 594163 206027 594787
rect 206039 594775 206040 594776
rect 206038 594774 206039 594775
rect 206536 594771 206617 594806
rect 206645 594797 206651 594799
rect 206536 594759 206623 594771
rect 206549 594704 206568 594759
rect 206577 594704 206623 594759
rect 206645 594732 206655 594797
rect 206583 594256 206630 594704
rect 206038 594175 206039 594176
rect 206039 594174 206040 594175
rect 206524 594163 206535 594174
rect 203247 594129 206535 594163
rect 206549 594151 206568 594256
rect 206577 594191 206623 594256
rect 206577 594179 206596 594191
rect 206617 594179 206623 594191
rect 206645 594228 206658 594732
rect 206645 594153 206655 594228
rect 206645 594151 206651 594153
rect 203247 593505 203281 594129
rect 203361 593505 203395 594129
rect 203407 594117 203408 594118
rect 204006 594117 204007 594118
rect 203406 594116 203407 594117
rect 204007 594116 204008 594117
rect 203406 593517 203407 593518
rect 204007 593517 204008 593518
rect 203407 593516 203408 593517
rect 204006 593516 204007 593517
rect 204019 593505 204053 594129
rect 204065 594117 204066 594118
rect 204664 594117 204665 594118
rect 204064 594116 204065 594117
rect 204665 594116 204666 594117
rect 204064 593517 204065 593518
rect 204665 593517 204666 593518
rect 204065 593516 204066 593517
rect 204664 593516 204665 593517
rect 204677 593505 204711 594129
rect 204723 594117 204724 594118
rect 205322 594117 205323 594118
rect 204722 594116 204723 594117
rect 205323 594116 205324 594117
rect 204722 593517 204723 593518
rect 205323 593517 205324 593518
rect 204723 593516 204724 593517
rect 205322 593516 205323 593517
rect 205335 593505 205369 594129
rect 205381 594117 205382 594118
rect 205980 594117 205981 594118
rect 205380 594116 205381 594117
rect 205981 594116 205982 594117
rect 205380 593517 205381 593518
rect 205981 593517 205982 593518
rect 205381 593516 205382 593517
rect 205980 593516 205981 593517
rect 205993 593505 206027 594129
rect 206039 594117 206040 594118
rect 206038 594116 206039 594117
rect 206536 594113 206617 594148
rect 206645 594139 206651 594141
rect 206536 594101 206623 594113
rect 206549 594052 206568 594101
rect 206577 594052 206623 594101
rect 206645 594080 206655 594139
rect 206583 593604 206630 594052
rect 206038 593517 206039 593518
rect 206039 593516 206040 593517
rect 206524 593505 206535 593516
rect 203247 593471 206535 593505
rect 206549 593493 206568 593604
rect 206577 593533 206623 593604
rect 206577 593521 206596 593533
rect 206617 593521 206623 593533
rect 206645 593576 206658 594080
rect 206645 593495 206655 593576
rect 206645 593493 206651 593495
rect 203247 592847 203281 593471
rect 203361 592847 203395 593471
rect 203407 593459 203408 593460
rect 204006 593459 204007 593460
rect 203406 593458 203407 593459
rect 204007 593458 204008 593459
rect 203406 592859 203407 592860
rect 204007 592859 204008 592860
rect 203407 592858 203408 592859
rect 204006 592858 204007 592859
rect 204019 592847 204053 593471
rect 204065 593459 204066 593460
rect 204664 593459 204665 593460
rect 204064 593458 204065 593459
rect 204665 593458 204666 593459
rect 204064 592859 204065 592860
rect 204665 592859 204666 592860
rect 204065 592858 204066 592859
rect 204664 592858 204665 592859
rect 204677 592847 204711 593471
rect 204723 593459 204724 593460
rect 205322 593459 205323 593460
rect 204722 593458 204723 593459
rect 205323 593458 205324 593459
rect 205335 592866 205369 593471
rect 205381 593459 205382 593460
rect 205980 593459 205981 593460
rect 205380 593458 205381 593459
rect 205981 593458 205982 593459
rect 205598 592866 205810 592996
rect 204722 592859 204723 592860
rect 204723 592858 204724 592859
rect 205154 592847 205810 592866
rect 205981 592859 205982 592860
rect 205980 592858 205981 592859
rect 205993 592847 206027 593471
rect 206039 593459 206040 593460
rect 206038 593458 206039 593459
rect 206536 593455 206617 593490
rect 206645 593481 206651 593483
rect 206536 593443 206623 593455
rect 206549 593382 206568 593443
rect 206577 593382 206623 593443
rect 206645 593410 206655 593481
rect 206583 592934 206630 593382
rect 206645 593342 206658 593410
rect 206685 593342 206697 594839
rect 206038 592859 206039 592860
rect 206039 592858 206040 592859
rect 206524 592847 206535 592858
rect 203247 592813 206535 592847
rect 206549 592835 206568 592934
rect 206577 592875 206623 592934
rect 206577 592863 206596 592875
rect 206617 592863 206623 592875
rect 206645 592835 206697 593342
rect 202142 592616 202532 592650
rect 201766 592149 202022 592152
rect 201794 592121 201994 592124
rect 202142 592118 202176 592616
rect 202356 592548 202403 592595
rect 202318 592514 202403 592548
rect 202245 592455 202290 592466
rect 202373 592455 202418 592466
rect 202256 592279 202290 592455
rect 202384 592279 202418 592455
rect 202356 592223 202403 592267
rect 202318 592201 202403 592223
rect 202302 592189 202403 592201
rect 202302 592170 202372 592189
rect 202498 592152 202532 592616
rect 202242 592149 202532 592152
rect 202276 592132 202396 592149
rect 202270 592121 202470 592124
rect 202270 592118 202424 592121
rect 202498 592118 202532 592149
rect 202142 592084 202532 592118
rect 202618 592616 203008 592650
rect 202618 592118 202652 592616
rect 202832 592548 202879 592595
rect 202794 592514 202879 592548
rect 202721 592455 202766 592466
rect 202849 592455 202894 592466
rect 202732 592279 202766 592455
rect 202860 592279 202894 592455
rect 202832 592223 202879 592267
rect 202794 592201 202879 592223
rect 202778 592189 202879 592201
rect 202778 592170 202848 592189
rect 202752 592132 202872 592134
rect 202974 592118 203008 592616
rect 202618 592084 203008 592118
rect 203247 592189 203281 592813
rect 203361 592189 203395 592813
rect 203407 592801 203408 592802
rect 204006 592801 204007 592802
rect 203406 592800 203407 592801
rect 204007 592800 204008 592801
rect 203406 592201 203407 592202
rect 204007 592201 204008 592202
rect 203407 592200 203408 592201
rect 204006 592200 204007 592201
rect 204019 592189 204053 592813
rect 204065 592801 204066 592802
rect 204664 592801 204665 592802
rect 204064 592800 204065 592801
rect 204665 592800 204666 592801
rect 204064 592201 204065 592202
rect 204665 592201 204666 592202
rect 204065 592200 204066 592201
rect 204664 592200 204665 592201
rect 204677 592189 204711 592813
rect 204723 592801 204724 592802
rect 204722 592800 204723 592801
rect 205154 592792 205810 592813
rect 205980 592801 205981 592802
rect 205981 592800 205982 592801
rect 204722 592201 204723 592202
rect 205323 592201 205324 592202
rect 204723 592200 204724 592201
rect 205322 592200 205323 592201
rect 205335 592189 205369 592792
rect 205598 592548 205810 592792
rect 205380 592201 205381 592202
rect 205981 592201 205982 592202
rect 205381 592200 205382 592201
rect 205980 592200 205981 592201
rect 205993 592189 206027 592813
rect 206039 592801 206040 592802
rect 206038 592800 206039 592801
rect 206536 592797 206617 592832
rect 206651 592825 206697 592835
rect 206536 592785 206623 592797
rect 206549 592720 206568 592785
rect 206577 592720 206623 592785
rect 206645 592720 206697 592825
rect 206583 592272 206617 592720
rect 206651 592272 206697 592720
rect 206038 592201 206039 592202
rect 206039 592200 206040 592201
rect 206524 592189 206535 592200
rect 203247 592155 206535 592189
rect 206549 592177 206568 592272
rect 206577 592217 206623 592272
rect 206577 592205 206596 592217
rect 206617 592205 206623 592217
rect 206645 592177 206697 592272
rect 202124 591928 202546 592034
rect 202600 591928 203022 592034
rect 202124 591716 203022 591928
rect 202124 591524 202546 591716
rect 202600 591524 203022 591716
rect 203247 591531 203281 592155
rect 203361 591531 203395 592155
rect 203407 592143 203408 592144
rect 204006 592143 204007 592144
rect 203406 592142 203407 592143
rect 204007 592142 204008 592143
rect 203406 591543 203407 591544
rect 204007 591543 204008 591544
rect 203407 591542 203408 591543
rect 204006 591542 204007 591543
rect 204019 591531 204053 592155
rect 204065 592143 204066 592144
rect 204664 592143 204665 592144
rect 204064 592142 204065 592143
rect 204665 592142 204666 592143
rect 204064 591543 204065 591544
rect 204665 591543 204666 591544
rect 204065 591542 204066 591543
rect 204664 591542 204665 591543
rect 204677 591531 204711 592155
rect 204723 592143 204724 592144
rect 205322 592143 205323 592144
rect 204722 592142 204723 592143
rect 205323 592142 205324 592143
rect 204722 591543 204723 591544
rect 205323 591543 205324 591544
rect 204723 591542 204724 591543
rect 205322 591542 205323 591543
rect 205335 591531 205369 592155
rect 205381 592143 205382 592144
rect 205980 592143 205981 592144
rect 205380 592142 205381 592143
rect 205981 592142 205982 592143
rect 205380 591543 205381 591544
rect 205981 591543 205982 591544
rect 205381 591542 205382 591543
rect 205980 591542 205981 591543
rect 205993 591531 206027 592155
rect 206039 592143 206040 592144
rect 206038 592142 206039 592143
rect 206536 592139 206617 592174
rect 206651 592167 206697 592177
rect 206536 592127 206623 592139
rect 206549 592062 206568 592127
rect 206577 592062 206623 592127
rect 206583 591614 206630 592062
rect 206038 591543 206039 591544
rect 206039 591542 206040 591543
rect 206524 591531 206535 591542
rect 198284 591497 203024 591524
rect 203247 591497 206535 591531
rect 206549 591519 206568 591614
rect 206577 591559 206623 591614
rect 206577 591547 206596 591559
rect 206617 591547 206623 591559
rect 206645 591519 206697 592167
rect 198284 591417 201758 591497
rect 202124 591490 202546 591497
rect 202600 591490 203022 591497
rect 201776 591463 203022 591490
rect 202124 591420 202546 591463
rect 202600 591420 203022 591463
rect 201852 591417 203022 591420
rect 203247 591417 203281 591497
rect 203361 591455 203395 591497
rect 204019 591468 204053 591497
rect 204677 591468 204711 591497
rect 205335 591468 205369 591497
rect 205993 591468 206027 591497
rect 206651 591468 206697 591519
rect 203991 591455 204053 591468
rect 204649 591455 204711 591468
rect 205307 591455 205369 591468
rect 205965 591455 206027 591468
rect 203361 591417 203401 591455
rect 203991 591427 204059 591455
rect 204649 591427 204717 591455
rect 205307 591427 205375 591455
rect 205965 591427 206033 591455
rect 206623 591427 206697 591468
rect 203411 591421 203429 591427
rect 203985 591421 204059 591427
rect 204069 591421 204087 591427
rect 204643 591421 204717 591427
rect 204727 591421 204745 591427
rect 205301 591421 205375 591427
rect 205385 591421 205403 591427
rect 205959 591421 206033 591427
rect 206043 591421 206061 591427
rect 206617 591421 206697 591427
rect 203407 591417 204059 591421
rect 204065 591417 204717 591421
rect 204723 591417 205375 591421
rect 205381 591417 206033 591421
rect 206039 591417 206697 591421
rect 198284 591383 206697 591417
rect 198284 591380 201758 591383
rect 198134 591378 201758 591380
rect 198170 591346 198204 591378
rect 198284 591347 201758 591378
rect 201852 591347 202822 591383
rect 198284 591346 198318 591347
rect 198168 591344 198424 591346
rect 198170 590521 198204 591344
rect 198284 591342 198318 591344
rect 198942 591342 198976 591347
rect 199600 591342 199634 591347
rect 200258 591342 200292 591347
rect 200916 591342 200950 591347
rect 201574 591342 201608 591347
rect 198266 591308 201642 591342
rect 198942 590521 198976 591308
rect 201724 591064 201736 591346
rect 201758 591098 201770 591320
rect 202106 590528 202568 590775
rect 198134 590485 201758 590521
rect 202124 590485 202546 590514
rect 203247 590485 203281 591383
rect 203383 591353 203401 591383
rect 203411 591381 203429 591383
rect 203985 591381 204003 591383
rect 204013 591353 204031 591383
rect 204041 591353 204059 591383
rect 204069 591381 204087 591383
rect 204643 591381 204661 591383
rect 204671 591353 204689 591383
rect 204699 591353 204717 591383
rect 204727 591381 204745 591383
rect 205301 591381 205319 591383
rect 205329 591353 205347 591383
rect 205357 591353 205375 591383
rect 205385 591381 205403 591383
rect 205959 591381 205977 591383
rect 205987 591353 206005 591383
rect 206015 591353 206033 591383
rect 206043 591381 206061 591383
rect 206617 591381 206635 591383
rect 206645 591353 206685 591383
rect 203361 591319 203395 591353
rect 204019 591319 204053 591353
rect 204677 591319 204711 591353
rect 205335 591319 205369 591353
rect 205993 591319 206027 591353
rect 206651 591319 206685 591353
rect 203343 591285 206697 591319
rect 206703 591285 206719 591319
rect 203361 590485 203395 590519
rect 204019 590485 204053 590519
rect 204677 590485 204711 590519
rect 205335 590485 205369 590519
rect 198134 590478 205827 590485
rect 197529 589701 197554 589752
rect 197557 589729 197582 589752
rect 198134 589719 201758 590478
rect 202124 590451 205827 590478
rect 201794 590404 201994 590405
rect 201766 590376 202022 590377
rect 202124 589894 202546 590451
rect 203094 590405 203150 590433
rect 202690 590400 203150 590405
rect 202950 590392 203150 590400
rect 202690 590372 203150 590377
rect 202922 590364 203150 590372
rect 203094 590336 203150 590364
rect 203247 590371 203281 590451
rect 203361 590371 203395 590451
rect 204019 590371 204053 590451
rect 204677 590371 204711 590451
rect 205335 590371 205369 590451
rect 205632 590371 205643 590382
rect 203247 590337 205643 590371
rect 202618 589962 203008 589996
rect 197644 589696 197920 589719
rect 198058 589696 201758 589719
rect 198134 589652 201758 589696
rect 202142 589713 202176 589894
rect 202318 589860 202403 589894
rect 202245 589801 202301 589812
rect 202373 589801 202429 589812
rect 202256 589752 202301 589801
rect 202384 589752 202429 589801
rect 202256 589713 202290 589752
rect 202301 589725 202302 589726
rect 202372 589725 202373 589726
rect 202302 589724 202303 589725
rect 202371 589724 202372 589725
rect 202384 589713 202418 589752
rect 202498 589713 202532 589894
rect 202142 589679 202532 589713
rect 202142 589652 202176 589679
rect 202256 589652 202290 589679
rect 202302 589667 202303 589668
rect 202371 589667 202372 589668
rect 202301 589666 202302 589667
rect 202372 589666 202373 589667
rect 202384 589652 202418 589679
rect 202498 589652 202532 589679
rect 202618 589713 202652 589962
rect 202832 589894 202879 589941
rect 202794 589860 202879 589894
rect 202974 589830 203008 589962
rect 202721 589801 202766 589812
rect 202849 589801 202894 589812
rect 202900 589806 203150 589830
rect 202974 589802 203008 589806
rect 202732 589713 202766 589801
rect 202777 589725 202778 589726
rect 202848 589725 202849 589726
rect 202778 589724 202779 589725
rect 202847 589724 202848 589725
rect 202860 589713 202894 589801
rect 202900 589778 203150 589802
rect 202974 589713 203008 589778
rect 203094 589750 203150 589778
rect 203247 589719 203281 590337
rect 202618 589679 203008 589713
rect 203166 589713 203328 589719
rect 203361 589713 203395 590337
rect 203407 590325 203408 590326
rect 204006 590325 204007 590326
rect 203406 590324 203407 590325
rect 204007 590324 204008 590325
rect 203406 589725 203407 589726
rect 204007 589725 204008 589726
rect 203407 589724 203408 589725
rect 204006 589724 204007 589725
rect 203436 589713 203478 589719
rect 203926 589713 203986 589719
rect 204019 589713 204053 590337
rect 204065 590325 204066 590326
rect 204664 590325 204665 590326
rect 204064 590324 204065 590325
rect 204665 590324 204666 590325
rect 204677 590196 204711 590337
rect 204723 590325 204724 590326
rect 205322 590325 205323 590326
rect 204722 590324 204723 590325
rect 205323 590324 205324 590325
rect 204656 589730 204730 590196
rect 204064 589725 204065 589726
rect 204065 589724 204066 589725
rect 204360 589713 204816 589730
rect 205323 589725 205324 589726
rect 205322 589724 205323 589725
rect 205335 589713 205369 590337
rect 205381 590325 205382 590326
rect 205380 590324 205381 590325
rect 205644 590309 205725 590356
rect 205691 589741 205725 590309
rect 205380 589725 205381 589726
rect 205381 589724 205382 589725
rect 205375 589713 205468 589719
rect 205632 589713 205643 589724
rect 203166 589696 205643 589713
rect 198134 589612 202592 589652
rect 198134 589596 201758 589612
rect 202142 589596 202176 589612
rect 202356 589596 202403 589612
rect 202498 589596 202532 589612
rect 198134 589556 202592 589596
rect 198134 589024 201758 589556
rect 202142 589464 202176 589556
rect 202318 589532 202403 589556
rect 202498 589464 202532 589556
rect 202142 589430 202532 589464
rect 202618 589464 202652 589679
rect 202732 589652 202766 589679
rect 202778 589667 202779 589668
rect 202847 589667 202848 589668
rect 202777 589666 202778 589667
rect 202848 589666 202849 589667
rect 202690 589613 202772 589652
rect 202860 589625 202894 589679
rect 202974 589624 203008 589679
rect 203247 589679 205643 589696
rect 202854 589622 203068 589624
rect 202854 589613 202900 589622
rect 202690 589612 202766 589613
rect 202832 589596 202879 589613
rect 202974 589596 203008 589622
rect 202690 589594 203068 589596
rect 202690 589585 202928 589594
rect 202690 589566 202828 589585
rect 202832 589566 202879 589585
rect 202690 589556 202879 589566
rect 202794 589532 202879 589556
rect 202974 589464 203008 589594
rect 202618 589430 203008 589464
rect 198134 589015 201774 589024
rect 198134 588996 201758 589015
rect 198134 588987 201774 588996
rect 189510 588654 192870 588688
rect 198134 588666 201758 588987
rect 202124 588934 202546 589380
rect 202600 588934 203022 589380
rect 201982 588916 203022 588934
rect 202124 588760 202546 588916
rect 202600 588760 203022 588916
rect 203247 589055 203281 589679
rect 203361 589055 203395 589679
rect 203407 589667 203408 589668
rect 204006 589667 204007 589668
rect 203406 589666 203407 589667
rect 204007 589666 204008 589667
rect 203930 589572 204013 589596
rect 203406 589067 203407 589068
rect 204007 589067 204008 589068
rect 203407 589066 203408 589067
rect 204006 589066 204007 589067
rect 204019 589055 204053 589679
rect 204065 589667 204066 589668
rect 204064 589666 204065 589667
rect 204360 589660 204816 589679
rect 205322 589667 205323 589668
rect 205323 589666 205324 589667
rect 204059 589572 204136 589596
rect 204584 589572 204636 589596
rect 204656 589542 204730 589660
rect 204744 589572 204798 589596
rect 205246 589572 205329 589596
rect 204064 589067 204065 589068
rect 204665 589067 204666 589068
rect 204065 589066 204066 589067
rect 204664 589066 204665 589067
rect 204677 589055 204711 589542
rect 204722 589067 204723 589068
rect 205323 589067 205324 589068
rect 204723 589066 204724 589067
rect 205322 589066 205323 589067
rect 205335 589055 205369 589679
rect 205381 589667 205382 589668
rect 205380 589666 205381 589667
rect 205644 589651 205725 589698
rect 205691 589083 205725 589651
rect 205380 589067 205381 589068
rect 205381 589066 205382 589067
rect 205632 589055 205643 589066
rect 203247 589021 205643 589055
rect 160606 588068 170990 588102
rect 160606 588032 165482 588068
rect 158928 587780 159030 587808
rect 158962 587746 158996 587774
rect 159044 587530 159444 587952
rect 159494 587900 160060 587934
rect 159494 587578 159528 587900
rect 159678 587820 159876 587831
rect 159562 587805 159664 587808
rect 159549 587780 159664 587805
rect 159689 587786 159876 587820
rect 159549 587758 159630 587780
rect 159877 587758 160005 587805
rect 159596 587720 159630 587758
rect 159924 587754 160005 587758
rect 159924 587720 159958 587754
rect 159865 587692 159876 587703
rect 159538 587656 159610 587662
rect 159689 587658 159876 587692
rect 159554 587600 159610 587606
rect 160026 587578 160060 587900
rect 159494 587544 160060 587578
rect 159080 587155 159114 587530
rect 159182 587522 159216 587530
rect 160092 587458 160726 587468
rect 165412 587155 165446 588032
rect 158691 587121 166865 587155
rect 159080 587102 159114 587121
rect 159120 587102 159176 587121
rect 159080 587098 159176 587102
rect 159080 587074 159114 587098
rect 159080 587053 159176 587074
rect 159080 587047 159263 587053
rect 158778 587042 159263 587047
rect 159080 587041 159114 587042
rect 159046 587007 159114 587041
rect 159135 587041 159263 587042
rect 165263 587041 165375 587053
rect 165412 587041 165446 587121
rect 159135 587038 165375 587041
rect 159135 587007 165360 587038
rect 165378 587007 165446 587041
rect 159080 586383 159114 587007
rect 159166 586995 159263 587007
rect 165263 586995 165360 587007
rect 159120 586966 159176 586980
rect 159120 586910 159176 586924
rect 159182 586880 159216 586995
rect 165310 586880 165344 586995
rect 165251 586852 165262 586863
rect 159135 586790 159216 586837
rect 159275 586818 165262 586852
rect 165263 586790 165344 586837
rect 159182 586396 159216 586790
rect 165310 586396 165344 586790
rect 165352 586476 165408 586482
rect 165352 586420 165406 586426
rect 159046 586349 159114 586383
rect 159135 586395 159216 586396
rect 165263 586395 165344 586396
rect 159135 586383 159263 586395
rect 165263 586383 165360 586395
rect 165412 586383 165446 587007
rect 159135 586349 165360 586383
rect 165378 586349 165446 586383
rect 159080 586080 159114 586349
rect 159166 586337 159263 586349
rect 165263 586337 165360 586349
rect 159182 586222 159216 586337
rect 165310 586222 165344 586337
rect 165412 586322 165446 586349
rect 165352 586298 166472 586322
rect 165352 586242 165408 586266
rect 165251 586194 165262 586205
rect 159275 586160 165262 586194
rect 165412 586080 165446 586298
rect 159080 586046 165446 586080
rect 159120 585762 160208 585766
rect 158790 585691 166766 585725
rect 160208 585626 160844 585632
rect 160152 585570 160900 585604
rect 169370 585338 169404 588068
rect 169410 586150 169430 587182
rect 169466 586150 169486 587238
rect 177970 585402 178004 586204
rect 178628 585402 178662 586204
rect 177520 585030 178700 585402
rect 164814 584906 166819 584934
rect 166865 584906 166878 584934
rect 147006 583954 156514 584024
rect 146946 583892 146956 583898
rect 147002 583892 156514 583954
rect 147006 583846 156514 583892
rect 134239 583652 142898 583686
rect 146324 583672 146344 583802
rect 146362 583730 146538 583782
rect 146358 583706 146840 583730
rect 146434 583668 146840 583706
rect 146946 583668 146956 583846
rect 147002 583668 156514 583846
rect 134239 583622 142208 583652
rect 142496 583622 142560 583652
rect 134239 583550 142760 583622
rect 134239 582460 142208 583550
rect 142396 583512 142454 583550
rect 142408 582460 142442 583512
rect 142496 582460 142560 583550
rect 142739 583500 142784 583511
rect 142750 582460 142784 583500
rect 142864 582460 142898 583652
rect 145264 583530 145624 583668
rect 146160 583556 156514 583668
rect 158559 583988 166997 584024
rect 171054 583988 171088 584114
rect 171168 583988 171202 584022
rect 171826 583988 171860 584022
rect 171940 583988 171974 584114
rect 172244 583988 172278 584114
rect 172358 583988 172392 584022
rect 158559 583954 172988 583988
rect 158559 583717 166997 583954
rect 158559 583567 168485 583717
rect 146160 583530 158154 583556
rect 145264 583496 158154 583530
rect 134239 582426 144068 582460
rect 134239 582358 142208 582426
rect 142408 582396 142442 582426
rect 142408 582374 142446 582396
rect 142396 582358 142454 582374
rect 142496 582358 142560 582426
rect 142750 582396 142784 582426
rect 142750 582358 142788 582396
rect 142864 582358 142898 582426
rect 143924 582396 143958 582426
rect 143166 582374 143204 582396
rect 143154 582358 143212 582374
rect 143520 582358 143958 582396
rect 134239 582324 143958 582358
rect 134239 581448 142208 582324
rect 142396 582286 142454 582324
rect 142408 581486 142442 582286
rect 142396 581448 142454 581486
rect 142496 581448 142560 582324
rect 142750 581486 142784 582324
rect 142750 581448 142788 581486
rect 142864 581448 142898 582324
rect 143154 582286 143212 582324
rect 143886 582290 143918 582314
rect 143166 581486 143200 582286
rect 143909 582274 143912 582285
rect 143914 582262 143918 582286
rect 143924 582274 143958 582324
rect 143920 581498 143958 582274
rect 143924 581486 143958 581498
rect 143154 581448 143212 581486
rect 143520 581448 143958 581486
rect 134239 581414 143958 581448
rect 134239 581346 142208 581414
rect 142396 581398 142454 581414
rect 142408 581370 142442 581398
rect 142408 581346 142453 581370
rect 142496 581346 142560 581414
rect 142750 581370 142784 581414
rect 142750 581346 142795 581370
rect 142864 581346 142898 581414
rect 143154 581398 143212 581414
rect 143890 581408 143904 581414
rect 143918 581380 143958 581414
rect 143924 581346 143958 581380
rect 144034 581346 144068 582426
rect 144892 581740 145214 581792
rect 144812 581370 145214 581740
rect 134239 581312 144068 581346
rect 134239 581002 142208 581312
rect 142408 581002 142453 581312
rect 142496 581002 142560 581312
rect 142750 581002 142795 581312
rect 142864 581002 142898 581312
rect 144892 581284 145214 581370
rect 145264 581230 145624 583496
rect 146160 582118 158154 583496
rect 146160 581850 156514 582118
rect 146160 581838 156856 581850
rect 146160 581230 147656 581838
rect 148896 581346 148930 581838
rect 149010 581498 149055 581838
rect 149342 581486 149387 581838
rect 150100 581486 150145 581838
rect 150858 581486 150903 581838
rect 151616 581486 151661 581838
rect 151970 581830 154278 581838
rect 151970 581672 154450 581830
rect 151782 581486 154450 581672
rect 149034 581448 154450 581486
rect 149072 581414 154450 581448
rect 149330 581398 149388 581414
rect 150088 581398 150146 581414
rect 150846 581398 150904 581414
rect 151604 581398 151662 581414
rect 151970 581346 154450 581414
rect 148896 581322 154450 581346
rect 148896 581312 154278 581322
rect 145554 581002 145588 581230
rect 145618 581140 145628 581148
rect 145646 581084 145684 581148
rect 146196 581002 146230 581230
rect 151970 581002 154278 581312
rect 154548 581002 156856 581838
rect 134239 580968 156856 581002
rect 134239 580908 142208 580968
rect 142408 580954 142453 580968
rect 134239 580888 137894 580908
rect 137906 580888 138282 580899
rect 138618 580888 138652 580908
rect 139346 580888 139410 580908
rect 139460 580894 139500 580908
rect 139518 580894 139528 580908
rect 139460 580888 139494 580894
rect 140118 580888 140168 580908
rect 140776 580888 140810 580908
rect 140892 580888 140926 580908
rect 141434 580888 141468 580908
rect 141510 580894 141538 580908
rect 141566 580894 141594 580908
rect 141650 580888 141684 580908
rect 142092 580888 142126 580908
rect 142408 580888 142442 580954
rect 142496 580888 142560 580968
rect 142750 580954 142795 580968
rect 142750 580948 142784 580954
rect 142864 580948 142898 580968
rect 143166 580948 143200 580968
rect 142692 580908 143328 580948
rect 142750 580892 142784 580908
rect 142864 580892 142898 580908
rect 143166 580892 143200 580908
rect 142636 580888 143328 580892
rect 143924 580888 143958 580968
rect 144682 580948 144716 580968
rect 144024 580908 145192 580948
rect 144682 580892 144716 580908
rect 144024 580888 145248 580892
rect 145276 580888 145310 580968
rect 134239 580866 145310 580888
rect 145442 580876 145476 580968
rect 145554 580888 145588 580968
rect 146196 580888 146230 580968
rect 146310 580888 146344 580968
rect 146356 580888 147056 580899
rect 147068 580888 147102 580968
rect 147114 580888 147814 580899
rect 147826 580888 147860 580968
rect 147872 580888 148474 580899
rect 148584 580888 148618 580968
rect 149342 580888 149376 580968
rect 150100 580888 150134 580968
rect 150858 580888 150892 580968
rect 151616 580888 151650 580968
rect 151676 580899 151684 580954
rect 151970 580899 154278 580968
rect 151676 580888 154470 580899
rect 154548 580888 156856 580968
rect 145440 580866 145476 580876
rect 134239 580864 145318 580866
rect 134239 580854 145412 580864
rect 134239 580842 137894 580854
rect 138550 580848 138612 580854
rect 137906 580842 137907 580843
rect 134239 580841 137906 580842
rect 134122 580694 134150 580750
rect 134239 580443 137905 580841
rect 138578 580820 138612 580846
rect 134239 580442 137906 580443
rect 138606 580442 138607 580443
rect 134239 580430 137894 580442
rect 137906 580441 137907 580442
rect 138605 580441 138606 580442
rect 137906 580430 138282 580441
rect 138618 580430 138652 580854
rect 138658 580848 138730 580854
rect 138658 580820 138702 580846
rect 138663 580442 138664 580443
rect 138664 580441 138665 580442
rect 139346 580430 139410 580854
rect 139460 580848 139494 580854
rect 140058 580848 140112 580854
rect 139422 580842 139423 580843
rect 139421 580841 139422 580842
rect 139460 580758 139500 580848
rect 139518 580758 139528 580848
rect 140086 580820 140112 580834
rect 139460 580514 139494 580758
rect 139421 580442 139422 580443
rect 139422 580441 139423 580442
rect 139460 580436 139500 580514
rect 139518 580436 139528 580514
rect 139460 580430 139494 580436
rect 140118 580430 140168 580854
rect 140174 580848 140238 580854
rect 140174 580820 140210 580834
rect 140776 580430 140810 580854
rect 140892 580430 140926 580854
rect 141434 580430 141468 580854
rect 141510 580758 141538 580848
rect 141566 580758 141594 580848
rect 141510 580436 141538 580514
rect 141566 580436 141594 580514
rect 141650 580430 141684 580854
rect 142092 580430 142126 580854
rect 142408 580430 142442 580854
rect 142636 580852 143328 580854
rect 142750 580430 142784 580852
rect 142864 580430 142898 580852
rect 143096 580848 143160 580852
rect 143124 580820 143160 580846
rect 143154 580442 143155 580443
rect 143153 580441 143154 580442
rect 143166 580430 143200 580852
rect 143206 580848 143276 580852
rect 143206 580820 143248 580846
rect 143911 580842 143912 580843
rect 143912 580841 143913 580842
rect 143211 580442 143212 580443
rect 143912 580442 143913 580443
rect 143212 580441 143213 580442
rect 143911 580441 143912 580442
rect 143924 580430 143958 580854
rect 144024 580852 145248 580854
rect 143970 580842 143971 580843
rect 144669 580842 144670 580843
rect 143969 580841 143970 580842
rect 144670 580841 144671 580842
rect 143969 580442 143970 580443
rect 144670 580442 144671 580443
rect 143970 580441 143971 580442
rect 144669 580441 144670 580442
rect 144682 580430 144716 580852
rect 144728 580842 144729 580843
rect 144727 580841 144728 580842
rect 145276 580838 145412 580854
rect 145434 580842 145476 580866
rect 145520 580854 145588 580888
rect 146162 580854 156856 580888
rect 145276 580826 145418 580838
rect 145276 580758 145318 580826
rect 145334 580758 145374 580826
rect 145276 580514 145310 580758
rect 145340 580514 145374 580758
rect 144727 580442 144728 580443
rect 144728 580441 144729 580442
rect 145276 580430 145318 580514
rect 145334 580446 145374 580514
rect 145340 580442 145374 580446
rect 145378 580758 145418 580826
rect 145378 580514 145412 580758
rect 145378 580446 145418 580514
rect 145378 580442 145412 580446
rect 145428 580442 145476 580842
rect 134239 580418 145318 580430
rect 145434 580418 145476 580442
rect 145554 580430 145588 580854
rect 146196 580430 146230 580854
rect 146244 580848 146304 580854
rect 146310 580842 146344 580854
rect 146350 580848 146424 580854
rect 146356 580842 146357 580843
rect 147055 580842 147056 580843
rect 147068 580842 147102 580854
rect 147114 580842 147115 580843
rect 147813 580842 147814 580843
rect 147826 580842 147860 580854
rect 147872 580842 147873 580843
rect 148571 580842 148572 580843
rect 146310 580841 146356 580842
rect 147056 580841 147057 580842
rect 147068 580841 147114 580842
rect 147814 580841 147815 580842
rect 147826 580841 147872 580842
rect 148572 580841 148573 580842
rect 146310 580838 146355 580841
rect 146272 580820 146304 580838
rect 146310 580820 146396 580838
rect 146310 580443 146355 580820
rect 147068 580443 147113 580841
rect 147826 580443 147871 580841
rect 146310 580442 146356 580443
rect 147056 580442 147057 580443
rect 147068 580442 147114 580443
rect 147814 580442 147815 580443
rect 147826 580442 147872 580443
rect 148572 580442 148573 580443
rect 146310 580430 146344 580442
rect 146356 580441 146357 580442
rect 147055 580441 147056 580442
rect 146356 580430 147056 580441
rect 147068 580430 147102 580442
rect 147114 580441 147115 580442
rect 147813 580441 147814 580442
rect 147114 580430 147814 580441
rect 147826 580430 147860 580442
rect 147872 580441 147873 580442
rect 148571 580441 148572 580442
rect 147872 580430 148474 580441
rect 148584 580430 148618 580854
rect 148630 580842 148631 580843
rect 149329 580842 149330 580843
rect 148629 580841 148630 580842
rect 149330 580841 149331 580842
rect 148629 580442 148630 580443
rect 149330 580442 149331 580443
rect 148630 580441 148631 580442
rect 149329 580441 149330 580442
rect 149342 580430 149376 580854
rect 149388 580842 149389 580843
rect 150087 580842 150088 580843
rect 149387 580841 149388 580842
rect 150088 580841 150089 580842
rect 149387 580442 149388 580443
rect 150088 580442 150089 580443
rect 149388 580441 149389 580442
rect 150087 580441 150088 580442
rect 150100 580430 150134 580854
rect 150786 580848 150852 580854
rect 150146 580842 150147 580843
rect 150845 580842 150846 580843
rect 150145 580841 150146 580842
rect 150846 580841 150847 580842
rect 150814 580820 150852 580830
rect 150145 580442 150146 580443
rect 150846 580442 150847 580443
rect 150146 580441 150147 580442
rect 150845 580441 150846 580442
rect 150858 580430 150892 580854
rect 150898 580848 150966 580854
rect 150904 580842 150905 580843
rect 151603 580842 151604 580843
rect 150903 580841 150904 580842
rect 151604 580841 151605 580842
rect 150898 580820 150938 580830
rect 150903 580442 150904 580443
rect 151604 580442 151605 580443
rect 150904 580441 150905 580442
rect 151603 580441 151604 580442
rect 151616 580430 151650 580854
rect 151662 580842 151663 580843
rect 151661 580841 151662 580842
rect 151661 580442 151662 580443
rect 151662 580441 151663 580442
rect 151676 580441 151684 580854
rect 151970 580441 154278 580854
rect 151676 580430 154470 580441
rect 154548 580430 156856 580854
rect 134239 580396 145310 580418
rect 145440 580408 145476 580418
rect 134239 580316 137894 580396
rect 138618 580316 138652 580396
rect 139346 580316 139410 580396
rect 139460 580390 139494 580396
rect 139460 580346 139500 580390
rect 139460 580316 139505 580346
rect 139518 580316 139528 580390
rect 140118 580346 140168 580396
rect 140776 580346 140810 580396
rect 140892 580346 140926 580396
rect 141434 580346 141468 580396
rect 140118 580316 140179 580346
rect 140776 580316 140821 580346
rect 140892 580316 140937 580346
rect 141434 580316 141479 580346
rect 141510 580316 141538 580390
rect 141566 580316 141594 580390
rect 141650 580346 141684 580396
rect 142092 580346 142126 580396
rect 142408 580346 142442 580396
rect 142750 580346 142784 580396
rect 141650 580316 141695 580346
rect 142092 580316 142137 580346
rect 142408 580316 142453 580346
rect 142750 580316 142795 580346
rect 142864 580316 142898 580396
rect 143166 580316 143200 580396
rect 143924 580316 143958 580396
rect 144682 580316 144716 580396
rect 145276 580374 145310 580396
rect 145222 580362 145310 580374
rect 145276 580316 145310 580362
rect 145442 580316 145476 580408
rect 145520 580396 145588 580430
rect 146162 580412 156856 580430
rect 146162 580396 155440 580412
rect 145554 580316 145588 580396
rect 146196 580316 146230 580396
rect 146310 580316 146344 580396
rect 147068 580316 147102 580396
rect 147826 580316 147860 580396
rect 148584 580316 148618 580396
rect 149342 580316 149376 580396
rect 150100 580316 150134 580396
rect 150858 580316 150892 580396
rect 151616 580316 151650 580396
rect 151676 580388 151684 580396
rect 152374 580316 152408 580396
rect 153132 580316 153166 580396
rect 153890 580316 153924 580396
rect 154648 580316 154682 580396
rect 155406 580316 155440 580396
rect 155590 580316 155624 580412
rect 134239 580282 155624 580316
rect 134064 579242 134110 579266
rect 122812 579210 122828 579214
rect 122840 579210 122884 579214
rect 112080 579172 120395 579208
rect 120414 579184 120430 579208
rect 112102 578974 112129 579136
rect 118760 579102 120395 579172
rect 122828 579158 122840 579210
rect 129280 579102 129314 579221
rect 129382 579204 129440 579221
rect 129494 579204 129532 579221
rect 130040 579204 130098 579221
rect 130252 579204 130290 579221
rect 130698 579204 130756 579221
rect 131010 579204 131048 579221
rect 131356 579204 131414 579221
rect 131768 579204 131806 579221
rect 132014 579204 132072 579221
rect 132526 579204 132564 579221
rect 132654 579210 132730 579221
rect 132672 579204 132730 579210
rect 129382 579170 129532 579204
rect 129584 579170 130290 579204
rect 130342 579170 131048 579204
rect 131100 579170 131806 579204
rect 131858 579170 132564 579204
rect 132616 579170 132730 579204
rect 129382 579154 129440 579170
rect 130040 579154 130098 579170
rect 130698 579154 130756 579170
rect 131356 579154 131414 579170
rect 132014 579154 132072 579170
rect 132672 579154 132730 579170
rect 129382 579139 129397 579154
rect 129394 579102 129428 579136
rect 130052 579102 130086 579136
rect 130710 579102 130744 579136
rect 131368 579102 131402 579136
rect 132026 579102 132060 579154
rect 132715 579139 132730 579154
rect 132684 579102 132718 579136
rect 132798 579102 132832 579221
rect 134239 579102 137863 580282
rect 138468 579554 138930 580192
rect 138526 579470 138876 579504
rect 138526 579102 138560 579470
rect 138618 579440 138652 579470
rect 138658 579456 138702 579470
rect 138658 579440 138748 579454
rect 138618 579402 138756 579440
rect 138618 579364 138652 579402
rect 138684 579368 138756 579402
rect 138730 579364 138748 579368
rect 138618 579332 138658 579364
rect 138664 579360 138686 579364
rect 138730 579360 138740 579364
rect 138758 579336 138776 579470
rect 138758 579332 138768 579336
rect 138618 579318 138652 579332
rect 138664 579318 138674 579329
rect 138717 579318 138762 579329
rect 138618 579254 138674 579318
rect 138640 579242 138674 579254
rect 138728 579242 138762 579318
rect 138640 579204 138686 579242
rect 138716 579204 138774 579242
rect 138640 579170 138774 579204
rect 138640 579156 138686 579170
rect 138628 579154 138686 579156
rect 138716 579154 138774 579170
rect 138628 579142 138674 579154
rect 138628 579136 138668 579142
rect 138734 579136 138774 579154
rect 138628 579130 138674 579136
rect 138640 579126 138674 579130
rect 138728 579130 138774 579136
rect 138728 579126 138762 579130
rect 138650 579102 138752 579126
rect 138842 579102 138876 579470
rect 139346 579266 139380 580282
rect 139460 579324 139505 580282
rect 139346 579242 139416 579266
rect 139460 579242 139500 579324
rect 139346 579170 139364 579242
rect 139448 579204 139506 579242
rect 139518 579210 139528 580282
rect 140118 579324 140179 580282
rect 140776 579324 140821 580282
rect 140892 579324 140937 580282
rect 141434 579324 141479 580282
rect 140118 579266 140168 579324
rect 140118 579242 140174 579266
rect 140776 579242 140810 579324
rect 140892 579266 140926 579324
rect 140886 579254 140926 579266
rect 140886 579242 140932 579254
rect 141434 579242 141468 579324
rect 140106 579204 140158 579242
rect 140184 579204 140214 579210
rect 140764 579204 140822 579242
rect 140864 579210 140932 579242
rect 140830 579204 140932 579210
rect 141422 579204 141480 579242
rect 141510 579210 141538 580282
rect 141566 579210 141594 580282
rect 141650 579324 141695 580282
rect 142092 579324 142137 580282
rect 142408 579324 142453 580282
rect 142750 579324 142795 580282
rect 141650 579254 141684 579324
rect 142092 579242 142126 579324
rect 142408 579254 142442 579324
rect 142750 579242 142784 579324
rect 141622 579204 141660 579242
rect 142080 579204 142138 579242
rect 142380 579204 142418 579242
rect 142738 579204 142796 579242
rect 139448 579182 140158 579204
rect 140180 579182 140932 579204
rect 139448 579170 140152 579182
rect 140180 579170 140186 579182
rect 140196 579170 140902 579182
rect 140954 579170 141660 579204
rect 141712 579170 142418 579204
rect 142470 579170 142796 579204
rect 139346 579102 139380 579170
rect 139448 579154 139506 579170
rect 140106 579154 140152 579170
rect 140764 579154 140822 579170
rect 141422 579154 141480 579170
rect 142080 579154 142138 579170
rect 142738 579154 142796 579170
rect 139448 579139 139463 579154
rect 139460 579102 139494 579136
rect 140118 579102 140152 579154
rect 140776 579102 140810 579136
rect 141434 579102 141468 579154
rect 142781 579139 142796 579154
rect 142092 579102 142126 579136
rect 142750 579102 142784 579136
rect 142864 579102 142898 580282
rect 143160 579242 143206 579266
rect 143918 579242 143964 579266
rect 144676 579242 144722 579266
rect 145434 579254 145474 579266
rect 145434 579242 145480 579254
rect 145554 579164 145588 580282
rect 112140 579012 112167 579098
rect 118760 579068 145492 579102
rect 118760 579032 120395 579068
rect 112102 578498 112129 578660
rect 112140 578536 112167 578622
rect 112222 578384 112842 578806
rect 112892 578754 113458 578788
rect 112892 578726 112926 578754
rect 113424 578726 113458 578754
rect 112858 578723 112926 578726
rect 113390 578723 113492 578726
rect 112892 578660 112926 578723
rect 113263 578674 113274 578685
rect 112892 578636 112932 578660
rect 112947 578654 113028 578659
rect 112940 578636 113028 578654
rect 113087 578640 113274 578674
rect 112892 578432 112926 578636
rect 112947 578612 113028 578636
rect 113275 578612 113356 578659
rect 112994 578574 113028 578612
rect 113322 578574 113356 578612
rect 113263 578546 113274 578557
rect 113087 578512 113274 578546
rect 113424 578432 113458 578723
rect 112892 578398 113458 578432
rect 112222 577908 112842 578330
rect 112892 578278 113458 578312
rect 112892 578206 112926 578278
rect 112892 578188 113064 578206
rect 113263 578198 113274 578209
rect 112892 578098 112926 578188
rect 112947 578178 113028 578183
rect 112940 578160 113036 578178
rect 113087 578164 113274 578198
rect 113286 578188 113394 578190
rect 113275 578162 113356 578183
rect 113275 578160 113366 578162
rect 112940 578105 112942 578160
rect 112947 578136 113028 578160
rect 113275 578136 113356 578160
rect 112994 578111 113028 578136
rect 113322 578111 113356 578136
rect 112978 578099 113075 578111
rect 113275 578099 113372 578111
rect 112978 578098 113372 578099
rect 113424 578098 113458 578278
rect 112892 578065 113458 578098
rect 112892 577956 112926 578065
rect 112940 578058 112942 578059
rect 113087 578053 113263 578065
rect 113087 578036 113274 578053
rect 113424 577956 113458 578065
rect 112892 577922 113458 577956
rect 118212 577938 120217 577966
rect 120263 577938 120276 577966
rect 112068 577522 120284 577533
rect 112079 577510 120273 577522
rect 112068 577499 120284 577510
rect 112095 577453 112129 577499
rect 112720 577490 112728 577499
rect 112914 577490 112920 577499
rect 112884 577441 113538 577462
rect 112188 577395 120164 577441
rect 112188 577385 120175 577395
rect 112095 576789 112129 577379
rect 112904 577364 113558 577385
rect 115918 577190 116366 577200
rect 115910 576988 116366 577190
rect 115910 576978 116358 576988
rect 113750 576794 114022 576821
rect 118854 576794 119310 576798
rect 112177 576783 120175 576794
rect 120223 576789 120257 577379
rect 112188 576773 120175 576783
rect 112188 576727 120164 576773
rect 118892 576713 119348 576727
rect 120189 576713 120291 576733
rect 120325 576713 120359 579032
rect 112095 576699 112129 576703
rect 118295 576679 121751 576713
rect 118295 576669 118329 576679
rect 118518 576676 119870 576679
rect 112057 576649 120295 576669
rect 120325 576649 120359 576679
rect 112057 576635 120359 576649
rect 112086 576550 112095 576584
rect 112068 576539 113602 576550
rect 112079 576527 113602 576539
rect 112068 576516 113602 576527
rect 111993 576342 112058 576454
rect 112095 576342 112096 576516
rect 112176 576448 112610 576495
rect 112768 576448 112815 576495
rect 113426 576448 113473 576495
rect 112200 576414 112815 576448
rect 112858 576414 113473 576448
rect 112100 576367 112129 576393
rect 112138 576367 112172 576376
rect 112100 576366 112176 576367
rect 112100 576342 112183 576366
rect 112785 576355 112830 576366
rect 113443 576355 113488 576366
rect 108862 576308 112414 576342
rect 108862 576108 108896 576308
rect 109172 576256 109218 576287
rect 109160 576240 109218 576256
rect 109038 576206 109218 576240
rect 109160 576159 109218 576206
rect 108965 576147 109010 576158
rect 108976 576108 109010 576147
rect 108720 576046 109016 576108
rect 108862 575716 108896 576046
rect 108976 575865 109010 576046
rect 109172 575877 109206 576159
rect 108964 575818 109023 575865
rect 109144 575818 109191 575865
rect 108964 575784 109191 575818
rect 108964 575768 109022 575784
rect 108964 575753 108979 575768
rect 109286 575716 109320 576308
rect 106390 575682 109320 575716
rect 109670 576154 109674 576159
rect 109670 575968 109698 576154
rect 106390 575646 108348 575682
rect 106410 575640 106444 575646
rect 88508 575574 106382 575608
rect 88508 575528 102756 575574
rect 102794 575528 102828 575574
rect 102856 575528 106382 575574
rect 88508 575492 106382 575528
rect 106384 575492 106390 575640
rect 106410 575492 106446 575640
rect 106722 575492 108348 575646
rect 88508 575458 108348 575492
rect 88508 575390 106382 575458
rect 106384 575448 106390 575458
rect 106410 575448 106446 575458
rect 106410 575390 106444 575448
rect 106722 575390 108348 575458
rect 88508 575356 108348 575390
rect 88508 575340 106382 575356
rect 88506 574876 106382 575340
rect 106410 574876 106444 575356
rect 106722 575136 108348 575356
rect 106722 574938 108372 575136
rect 106848 574876 106893 574938
rect 107466 574876 107500 574938
rect 107506 574876 107538 574938
rect 107580 574876 107614 574938
rect 88506 574100 107676 574876
rect 86640 574034 107676 574100
rect 107946 574846 108348 574882
rect 108862 574846 108896 575682
rect 109670 575282 109674 575968
rect 109938 575220 109972 576308
rect 110052 576271 110099 576287
rect 110040 576240 110099 576271
rect 110264 576240 110311 576287
rect 110710 576256 110757 576287
rect 110698 576240 110757 576256
rect 110922 576240 110969 576287
rect 111124 576240 111516 576308
rect 110040 576206 110311 576240
rect 110354 576206 110969 576240
rect 111012 576206 111516 576240
rect 110040 576159 110098 576206
rect 110698 576159 110756 576206
rect 110052 575381 110086 576159
rect 110281 576147 110326 576158
rect 110292 575369 110326 576147
rect 110710 575381 110744 576159
rect 110939 576148 110984 576158
rect 110926 576012 111004 576148
rect 111124 576012 111516 576206
rect 111630 576172 111648 576274
rect 111658 576200 111704 576246
rect 111993 576240 112058 576308
rect 112095 576287 112183 576308
rect 112095 576240 112185 576287
rect 112238 576240 112285 576287
rect 111993 576206 112285 576240
rect 110926 575960 111516 576012
rect 110950 575866 111516 575960
rect 110950 575369 110984 575866
rect 110280 575322 110339 575369
rect 110682 575322 110729 575369
rect 110938 575322 110997 575369
rect 111124 575364 111516 575866
rect 111340 575322 111387 575364
rect 110114 575288 110729 575322
rect 110772 575288 111387 575322
rect 110280 575272 110338 575288
rect 110938 575272 110996 575288
rect 110292 575220 110332 575272
rect 111482 575220 111516 575364
rect 109938 575186 111516 575220
rect 111993 576088 112058 576206
rect 112095 576159 112184 576206
rect 112095 576131 112129 576159
rect 112104 576115 112129 576131
rect 112138 576103 112172 576159
rect 112255 576147 112300 576158
rect 112266 576103 112300 576147
rect 112380 576103 112414 576308
rect 112784 576115 112785 576116
rect 112783 576114 112784 576115
rect 112796 576103 112830 576355
rect 112841 576115 112842 576116
rect 113442 576115 113443 576116
rect 112842 576114 112843 576115
rect 113441 576114 113442 576115
rect 113454 576103 113488 576355
rect 113568 576103 113602 576516
rect 114128 576548 117680 576552
rect 118295 576548 118329 576635
rect 118424 576611 120176 576635
rect 120223 576611 120257 576635
rect 120325 576611 120359 576635
rect 121584 576617 121616 576630
rect 121640 576617 121644 576658
rect 118471 576577 119086 576611
rect 119129 576577 119744 576611
rect 119787 576584 120359 576611
rect 119787 576577 120367 576584
rect 120223 576552 120257 576577
rect 120294 576571 120367 576577
rect 120433 576571 120516 576584
rect 120964 576571 121025 576584
rect 121091 576571 121168 576584
rect 121616 576571 121640 576584
rect 120325 576552 120359 576571
rect 121584 576552 121616 576571
rect 121640 576552 121644 576571
rect 114128 576518 119468 576548
rect 119714 576518 119770 576529
rect 114128 576103 114162 576518
rect 114872 576450 114919 576497
rect 115530 576450 115577 576497
rect 115910 576450 116358 576518
rect 116574 576514 119468 576518
rect 116574 576450 116608 576514
rect 116846 576450 116893 576497
rect 114304 576416 114919 576450
rect 114962 576416 115577 576450
rect 115620 576446 116893 576450
rect 116920 576450 116936 576493
rect 117504 576450 117551 576497
rect 116920 576446 117551 576450
rect 117646 576493 117680 576514
rect 118295 576493 118329 576514
rect 118409 576496 118454 576514
rect 119067 576496 119112 576514
rect 118409 576493 118443 576496
rect 119067 576493 119101 576496
rect 117646 576446 117693 576493
rect 117976 576446 118023 576493
rect 118295 576446 118342 576493
rect 118409 576462 118456 576493
rect 118397 576446 118456 576462
rect 118634 576446 118681 576493
rect 119067 576462 119114 576493
rect 119055 576446 119114 576462
rect 119292 576446 119339 576493
rect 115620 576416 118023 576446
rect 114231 576357 114276 576368
rect 114889 576357 114934 576368
rect 115547 576357 115592 576368
rect 114242 576103 114276 576357
rect 114287 576115 114288 576116
rect 114888 576115 114889 576116
rect 114288 576114 114289 576115
rect 114887 576114 114888 576115
rect 114900 576103 114934 576357
rect 115558 576196 115592 576357
rect 115910 576312 116358 576416
rect 116192 576196 116270 576312
rect 116290 576196 116320 576248
rect 114945 576115 114946 576116
rect 115546 576115 115547 576116
rect 114946 576114 114947 576115
rect 115545 576114 115546 576115
rect 115558 576109 115598 576196
rect 116192 576192 116290 576196
rect 116320 576192 116346 576196
rect 116192 576178 116270 576192
rect 116290 576178 116320 576192
rect 115603 576115 115604 576116
rect 115604 576114 115605 576115
rect 115558 576103 115592 576109
rect 116190 576103 116358 576178
rect 116574 576166 116608 576416
rect 116750 576412 117365 576416
rect 117408 576412 118023 576416
rect 118066 576412 118681 576446
rect 118724 576412 119339 576446
rect 116862 576365 116920 576369
rect 117520 576365 117578 576369
rect 116677 576353 116722 576364
rect 116863 576357 116908 576365
rect 116574 576148 116644 576166
rect 116574 576110 116608 576148
rect 116574 576103 116644 576110
rect 116688 576103 116722 576353
rect 116874 576103 116908 576357
rect 117335 576353 117380 576364
rect 117521 576357 117566 576365
rect 117346 576103 117380 576353
rect 117532 576103 117566 576357
rect 117646 576103 117680 576412
rect 117993 576353 118038 576364
rect 117992 576115 117993 576116
rect 117991 576114 117992 576115
rect 118004 576103 118038 576353
rect 118040 576109 118044 576196
rect 118126 576148 118182 576166
rect 118049 576115 118050 576116
rect 118050 576114 118051 576115
rect 118126 576103 118182 576110
rect 118295 576103 118329 576412
rect 118397 576365 118455 576412
rect 119055 576365 119113 576412
rect 118409 576103 118443 576365
rect 118651 576353 118696 576364
rect 118662 576103 118696 576353
rect 119067 576108 119101 576365
rect 119309 576353 119354 576364
rect 118868 576103 119164 576108
rect 119320 576103 119354 576353
rect 119434 576103 119468 576514
rect 119725 576496 119770 576518
rect 120086 576518 121664 576552
rect 119713 576115 119714 576116
rect 119712 576114 119713 576115
rect 119725 576103 119759 576496
rect 119770 576115 119771 576116
rect 119771 576114 119772 576115
rect 120086 576103 120120 576518
rect 120223 576496 120304 576518
rect 120325 576497 120359 576518
rect 120383 576497 120393 576518
rect 121616 576515 121664 576518
rect 120223 576450 120257 576496
rect 120322 576450 121535 576497
rect 120223 576416 120877 576450
rect 120920 576416 121535 576450
rect 120223 576391 120257 576416
rect 120223 576368 120268 576391
rect 120189 576357 120268 576368
rect 120200 576131 120268 576357
rect 120200 576115 120245 576131
rect 120164 576103 120175 576114
rect 111993 576041 112129 576088
rect 111993 575430 112058 576041
rect 112095 575473 112129 576041
rect 112104 575457 112129 575473
rect 112138 576069 112183 576103
rect 112188 576069 113602 576103
rect 114094 576069 120180 576103
rect 120200 576088 120234 576115
rect 112138 575445 112172 576069
rect 112266 575445 112300 576069
rect 112380 575445 112414 576069
rect 112783 576057 112784 576058
rect 112784 576056 112785 576057
rect 112784 575457 112785 575458
rect 112783 575456 112784 575457
rect 112796 575445 112830 576069
rect 112842 576057 112843 576058
rect 113441 576057 113442 576058
rect 112841 576056 112842 576057
rect 113442 576056 113443 576057
rect 113010 575866 113260 576012
rect 113074 575752 113228 575866
rect 112841 575457 112842 575458
rect 113442 575457 113443 575458
rect 112842 575456 112843 575457
rect 113441 575456 113442 575457
rect 113454 575445 113488 576069
rect 113568 575445 113602 576069
rect 114128 575445 114162 576069
rect 114242 575445 114276 576069
rect 114288 576057 114289 576058
rect 114887 576057 114888 576058
rect 114287 576056 114288 576057
rect 114888 576056 114889 576057
rect 114287 575457 114288 575458
rect 114888 575457 114889 575458
rect 114288 575456 114289 575457
rect 114887 575456 114888 575457
rect 114900 575445 114934 576069
rect 115558 576063 115592 576069
rect 114946 576057 114947 576058
rect 115545 576057 115546 576058
rect 114945 576056 114946 576057
rect 115546 576056 115547 576057
rect 115558 576018 115598 576063
rect 115604 576057 115605 576058
rect 115603 576056 115604 576057
rect 115558 575940 115592 576018
rect 116190 576010 116358 576069
rect 116176 576008 116358 576010
rect 116574 576046 116644 576069
rect 116574 576018 116608 576046
rect 116176 575992 116210 576008
rect 116144 575972 116210 575982
rect 116216 575972 116250 576008
rect 116256 575992 116320 576008
rect 116574 575990 116644 576018
rect 115598 575940 116250 575972
rect 116256 575964 116320 575982
rect 115558 575878 116250 575940
rect 116264 575958 116320 575964
rect 116574 575958 116608 575990
rect 116688 575958 116722 576069
rect 116264 575936 116834 575958
rect 116268 575924 116834 575936
rect 116268 575878 116302 575924
rect 115558 575829 116366 575878
rect 116574 575844 116608 575924
rect 116688 575861 116722 575924
rect 116800 575865 116834 575924
rect 116874 575956 116908 576069
rect 116874 575865 116919 575956
rect 117346 575877 117380 576069
rect 117532 575865 117566 576069
rect 117646 575865 117680 576069
rect 117991 576057 117992 576058
rect 117992 576056 117993 576057
rect 117986 576002 117996 576012
rect 117982 575982 117996 576002
rect 118004 575877 118038 576069
rect 118040 576012 118044 576063
rect 118050 576057 118051 576058
rect 118049 576056 118050 576057
rect 118126 576046 118182 576069
rect 118040 576002 118058 576012
rect 118040 575982 118062 576002
rect 118126 575990 118182 576018
rect 118295 575865 118329 576069
rect 118409 575874 118443 576069
rect 118662 575877 118696 576069
rect 118868 576046 119164 576069
rect 119067 575874 119101 576046
rect 119320 576002 119354 576069
rect 119310 575932 119362 576002
rect 119194 575876 119362 575932
rect 118409 575865 118454 575874
rect 119067 575865 119112 575874
rect 119194 575865 119330 575876
rect 116639 575844 116650 575855
rect 115558 575744 116404 575829
rect 116463 575810 116650 575844
rect 115558 575718 116394 575744
rect 115558 575666 116366 575718
rect 116574 575716 116608 575810
rect 116651 575782 116732 575829
rect 116800 575818 117024 575865
rect 117318 575818 117365 575865
rect 117520 575818 117579 575865
rect 117646 575818 117693 575865
rect 117976 575818 118023 575865
rect 118282 575818 119339 575865
rect 116734 575784 117365 575818
rect 117408 575784 118023 575818
rect 118066 575784 118681 575818
rect 118724 575784 119339 575818
rect 116698 575728 116732 575782
rect 116639 575716 116650 575727
rect 116800 575716 116834 575784
rect 116862 575768 116920 575784
rect 117520 575768 117578 575784
rect 116874 575716 116919 575768
rect 117532 575716 117566 575768
rect 117646 575716 117680 575784
rect 118295 575716 118329 575784
rect 118397 575768 118455 575784
rect 119055 575768 119113 575784
rect 118409 575716 118454 575768
rect 119067 575716 119112 575768
rect 119434 575716 119468 576069
rect 119712 576057 119713 576058
rect 119713 576056 119714 576057
rect 116463 575682 119468 575716
rect 119725 575874 119759 576069
rect 119771 576057 119772 576058
rect 119770 576056 119771 576057
rect 115558 575550 116250 575666
rect 116268 575602 116302 575666
rect 116800 575602 116834 575682
rect 116268 575568 116834 575602
rect 115558 575458 115603 575550
rect 114945 575457 114946 575458
rect 115546 575457 115547 575458
rect 115558 575457 115604 575458
rect 116204 575457 116205 575458
rect 114946 575456 114947 575457
rect 115545 575456 115546 575457
rect 115456 575445 115546 575456
rect 115558 575445 115592 575457
rect 115604 575456 115605 575457
rect 116203 575456 116204 575457
rect 115604 575445 115674 575456
rect 116216 575445 116250 575550
rect 116874 575458 116919 575682
rect 116261 575457 116262 575458
rect 116862 575457 116863 575458
rect 116874 575457 116920 575458
rect 117520 575457 117521 575458
rect 116262 575456 116263 575457
rect 116861 575456 116862 575457
rect 116802 575445 116862 575456
rect 116874 575445 116908 575457
rect 116920 575456 116921 575457
rect 117519 575456 117520 575457
rect 116920 575445 117024 575456
rect 117532 575445 117566 575682
rect 117646 575445 117680 575682
rect 118295 575445 118329 575682
rect 118409 575458 118454 575682
rect 119050 575466 119120 575682
rect 118409 575457 118455 575458
rect 118409 575445 118443 575457
rect 118455 575456 118456 575457
rect 118876 575456 119332 575466
rect 119725 575458 119770 575874
rect 119713 575457 119714 575458
rect 119725 575457 119771 575458
rect 119712 575456 119713 575457
rect 118455 575445 119713 575456
rect 119725 575445 119759 575457
rect 119771 575456 119772 575457
rect 120086 575456 120120 576069
rect 120187 576041 120257 576088
rect 120200 575874 120268 576041
rect 120200 575473 120304 575874
rect 119771 575445 120175 575456
rect 111993 575383 112129 575430
rect 111993 575218 112058 575383
rect 112095 575252 112129 575383
rect 112138 575411 112183 575445
rect 112188 575422 113602 575445
rect 114094 575424 117680 575445
rect 118261 575424 120175 575445
rect 120200 575430 120245 575473
rect 120187 575428 120304 575430
rect 114094 575422 120175 575424
rect 112188 575411 120175 575422
rect 112138 575379 112172 575411
rect 112200 575405 112236 575411
rect 112138 575363 112163 575379
rect 112200 575372 112204 575405
rect 112266 575367 112300 575411
rect 112380 575367 112414 575411
rect 112734 575405 112890 575411
rect 113388 575405 114236 575411
rect 112783 575399 112784 575400
rect 112784 575398 112785 575399
rect 112790 575367 112836 575405
rect 112842 575399 112843 575400
rect 112841 575398 112842 575399
rect 113426 575378 113520 575405
rect 113428 575370 113518 575378
rect 113448 575367 113494 575370
rect 112200 575344 112232 575366
rect 112254 575320 112313 575367
rect 112380 575320 112427 575367
rect 112768 575366 112815 575367
rect 113426 575366 113473 575367
rect 112762 575339 112864 575366
rect 113398 575350 113548 575366
rect 113400 575342 113546 575350
rect 113420 575339 113522 575342
rect 112768 575320 112815 575339
rect 113426 575320 113473 575339
rect 112200 575286 112815 575320
rect 112858 575286 113473 575320
rect 112254 575270 112312 575286
rect 112086 575218 112129 575252
rect 112266 575218 112300 575270
rect 112380 575218 112414 575286
rect 113568 575218 113602 575405
rect 107946 574812 110218 574846
rect 107946 574070 108348 574812
rect 108798 574448 108820 574658
rect 108862 574070 108896 574812
rect 108964 574744 109044 574791
rect 109384 574744 109431 574791
rect 109634 574760 109681 574791
rect 109622 574744 109681 574760
rect 110042 574744 110089 574791
rect 108964 574710 109431 574744
rect 109474 574710 110089 574744
rect 108964 574663 109022 574710
rect 109622 574663 109680 574710
rect 108976 574070 109021 574663
rect 109401 574651 109446 574662
rect 109412 574374 109446 574651
rect 109634 574374 109668 574663
rect 110059 574651 110104 574662
rect 110070 574374 110104 574651
rect 107946 574034 109058 574070
rect 86640 574000 109058 574034
rect 86640 573931 107676 574000
rect 107946 573931 109058 574000
rect 86640 573894 109058 573931
rect 86640 573860 109320 573894
rect 86640 573792 109058 573860
rect 109144 573792 109191 573839
rect 86640 573758 109191 573792
rect 86640 573616 109058 573758
rect 109161 573699 109206 573710
rect 109172 573663 109206 573699
rect 109172 573616 109219 573663
rect 109286 573616 109320 573860
rect 109412 573842 109457 574374
rect 109634 573842 109679 574374
rect 110070 573898 110115 574374
rect 110184 573898 110218 574812
rect 110292 574732 110332 575186
rect 111993 575184 113602 575218
rect 111993 575152 112027 575184
rect 112095 575152 112129 575184
rect 112266 575152 112300 575184
rect 112380 575152 112414 575184
rect 114128 575152 114162 575405
rect 114242 575152 114276 575411
rect 114282 575405 114342 575411
rect 114838 575405 114894 575411
rect 114288 575399 114289 575400
rect 114887 575399 114888 575400
rect 114287 575398 114288 575399
rect 114888 575398 114889 575399
rect 114900 575152 114934 575411
rect 114940 575405 114992 575411
rect 114936 575366 114940 575405
rect 114946 575399 114947 575400
rect 115545 575399 115546 575400
rect 115558 575399 115592 575411
rect 115604 575399 115605 575400
rect 116203 575399 116204 575400
rect 114945 575398 114946 575399
rect 115546 575398 115547 575399
rect 115558 575398 115604 575399
rect 116204 575398 116205 575399
rect 115558 575202 115603 575398
rect 115558 575152 115592 575202
rect 116216 575182 116250 575411
rect 116816 575405 116868 575411
rect 116262 575399 116263 575400
rect 116261 575398 116262 575399
rect 116292 575370 116308 575405
rect 116264 575312 116308 575370
rect 116320 575312 116364 575405
rect 116861 575399 116862 575400
rect 116874 575399 116908 575411
rect 116914 575405 116970 575411
rect 117466 575405 117526 575411
rect 116920 575399 116921 575400
rect 117519 575399 117520 575400
rect 116862 575398 116863 575399
rect 116874 575398 116920 575399
rect 117520 575398 117521 575399
rect 116874 575184 116919 575398
rect 115910 575152 116358 575182
rect 116874 575152 116908 575184
rect 117532 575152 117566 575411
rect 117572 575405 118268 575411
rect 117646 575152 117680 575405
rect 118212 575349 118268 575368
rect 118295 575152 118329 575411
rect 118409 575399 118443 575411
rect 118455 575399 118456 575400
rect 118409 575398 118455 575399
rect 118409 575152 118454 575398
rect 118876 575396 119332 575411
rect 119712 575399 119713 575400
rect 119725 575399 119759 575411
rect 119771 575399 119772 575400
rect 119713 575398 119714 575399
rect 119725 575398 119771 575399
rect 119050 575246 119120 575396
rect 119067 575152 119112 575246
rect 119725 575152 119770 575398
rect 120086 575220 120120 575411
rect 120176 575381 120304 575428
rect 120223 575369 120304 575381
rect 120325 575369 120359 576416
rect 120371 576369 120429 576416
rect 121029 576369 121087 576416
rect 120383 575369 120428 576369
rect 120847 576357 120903 576368
rect 120858 575381 120903 576357
rect 121041 575369 121086 576369
rect 121505 576357 121561 576368
rect 121516 575381 121561 576357
rect 120215 575322 121535 575369
rect 120223 575288 120877 575322
rect 120920 575288 121535 575322
rect 120223 575233 120304 575288
rect 120176 575220 120304 575233
rect 120325 575220 120359 575288
rect 120371 575272 120429 575288
rect 121029 575272 121087 575288
rect 120383 575220 120393 575272
rect 121584 575220 121616 575230
rect 121630 575220 121664 576515
rect 120086 575186 121664 575220
rect 120223 575152 120304 575186
rect 120325 575152 120359 575186
rect 120383 575152 120393 575186
rect 111980 574758 120400 575152
rect 110270 574720 110278 574732
rect 110266 574468 110278 574720
rect 110270 574456 110278 574468
rect 110272 574446 110278 574456
rect 110292 574446 110326 574732
rect 110292 573898 110332 574446
rect 111980 574430 120417 574758
rect 120424 574468 120455 574720
rect 111980 574059 120400 574430
rect 121584 574059 121616 575186
rect 121640 574059 121644 575186
rect 121699 575058 121733 576518
rect 121813 575058 121847 576617
rect 121882 576586 121883 576749
rect 124452 576718 124486 577146
rect 124566 576718 124600 576752
rect 125224 576718 125258 576752
rect 125338 576718 125372 577146
rect 125642 576718 125676 577146
rect 125756 576718 125790 576752
rect 126414 576718 126448 576752
rect 126528 576718 126562 577146
rect 123462 576684 126822 576718
rect 124452 576588 124486 576684
rect 125218 576654 125220 576658
rect 124554 576588 124806 576654
rect 124820 576616 125270 576654
rect 124858 576588 125270 576616
rect 125338 576588 125372 576684
rect 125642 576588 125676 576684
rect 125744 576588 126122 576654
rect 126136 576616 126460 576654
rect 126174 576588 126460 576616
rect 126528 576588 126562 576684
rect 126952 576588 126972 576772
rect 129280 576767 129314 579068
rect 131368 578672 131402 579068
rect 130926 578434 131640 578672
rect 132026 578434 132060 579068
rect 130918 578062 132098 578434
rect 131368 576768 131402 578062
rect 132026 576768 132060 578062
rect 132650 577236 132674 577526
rect 132684 577236 132708 577526
rect 129382 576767 132730 576768
rect 129280 576749 132730 576767
rect 127838 576588 127872 576606
rect 122136 575148 122137 576586
rect 122882 575354 122884 575382
rect 122882 575340 122956 575354
rect 122966 575340 123038 575354
rect 122882 575284 122928 575326
rect 122994 575284 123038 575326
rect 123330 575148 123786 576586
rect 124240 576584 127872 576588
rect 124060 576576 124122 576584
rect 124188 576576 127872 576584
rect 121699 574354 122080 575058
rect 121699 574059 121733 574354
rect 111980 574025 121745 574059
rect 111980 574004 120400 574025
rect 121584 574004 121616 574025
rect 121640 574004 121644 574025
rect 121699 574004 121733 574025
rect 111980 573957 121733 574004
rect 111980 573945 120400 573957
rect 111980 573932 112450 573945
rect 109938 573864 111516 573898
rect 109412 573675 109446 573842
rect 109634 573663 109668 573842
rect 109384 573616 109431 573663
rect 109622 573616 109681 573663
rect 109938 573616 109972 573864
rect 110070 573842 110115 573864
rect 110184 573843 110218 573864
rect 110292 573843 110332 573864
rect 110070 573796 110104 573842
rect 110171 573796 110546 573843
rect 110682 573796 110729 573843
rect 110937 573796 111387 573843
rect 110070 573762 110729 573796
rect 110772 573766 111387 573796
rect 111482 573766 111516 573864
rect 110772 573762 111516 573766
rect 110070 573714 110104 573762
rect 110041 573703 110104 573714
rect 110052 573675 110104 573703
rect 110052 573663 110097 573675
rect 110042 573659 110097 573663
rect 110042 573616 110089 573659
rect 86640 573582 109431 573616
rect 109474 573582 110089 573616
rect 86640 573514 109058 573582
rect 109172 573514 109206 573582
rect 109286 573514 109320 573582
rect 109622 573566 109680 573582
rect 109670 573514 109674 573566
rect 109938 573514 109972 573582
rect 110052 573514 110086 573582
rect 110184 573514 110218 573762
rect 110280 573715 110338 573762
rect 110938 573715 110996 573762
rect 86640 573480 110218 573514
rect 86640 573428 109058 573480
rect 86640 573398 106382 573428
rect 106390 573398 109058 573428
rect 86640 573392 109058 573398
rect 86640 573370 106382 573392
rect 106390 573370 109058 573392
rect 86640 573364 109058 573370
rect 86640 573348 106382 573364
rect 106390 573348 109058 573364
rect 86640 573314 109058 573348
rect 86640 573270 106382 573314
rect 86640 573088 102756 573270
rect 102794 573088 102828 573270
rect 102856 573152 106382 573270
rect 106390 573278 109058 573314
rect 109172 573306 109206 573480
rect 109286 573306 109320 573480
rect 109670 573306 109674 573480
rect 109938 573306 109972 573480
rect 110052 573306 110086 573480
rect 110292 573418 110337 573715
rect 110699 573703 110744 573714
rect 110292 573310 110326 573418
rect 110710 573310 110744 573703
rect 110950 573358 110995 573715
rect 111124 573358 111516 573762
rect 110950 573310 111516 573358
rect 111980 573728 113638 573932
rect 114092 573930 117824 573945
rect 118094 573930 120400 573945
rect 114092 573898 120400 573930
rect 120405 573898 120423 573957
rect 120433 573923 121060 573957
rect 120433 573917 120451 573923
rect 121007 573917 121025 573923
rect 121035 573898 121053 573923
rect 121063 573898 121081 573957
rect 121091 573923 121733 573957
rect 121091 573917 121109 573923
rect 121584 573898 121616 573917
rect 121640 573898 121644 573917
rect 114092 573864 121664 573898
rect 114092 573843 120400 573864
rect 114092 573796 121428 573843
rect 121488 573796 121535 573843
rect 114092 573762 120877 573796
rect 120920 573762 121535 573796
rect 111980 573714 113894 573728
rect 114092 573715 120429 573762
rect 121029 573715 121087 573762
rect 111980 573310 113638 573714
rect 102856 573102 106384 573152
rect 102856 573088 106382 573102
rect 86640 573064 106382 573088
rect 106390 573064 108896 573278
rect 108942 573164 108962 573278
rect 108976 573211 109010 573278
rect 108964 573182 109022 573211
rect 108964 573164 109023 573182
rect 109060 573164 110086 573306
rect 108964 573130 110086 573164
rect 86640 573062 108896 573064
rect 108942 573062 108962 573130
rect 108964 573114 109022 573130
rect 108964 573099 108996 573114
rect 108976 573062 108996 573099
rect 109060 573062 110086 573130
rect 86640 573030 110086 573062
rect 86640 573000 106382 573030
rect 106390 573028 110086 573030
rect 106390 573000 108896 573028
rect 86640 572992 108896 573000
rect 86640 572962 107088 572992
rect 107102 572962 107746 572992
rect 107760 572962 108404 572992
rect 86640 572928 106444 572962
rect 106482 572928 107088 572962
rect 107140 572928 107746 572962
rect 107798 572928 108404 572962
rect 86640 572838 106382 572928
rect 106410 572889 106444 572928
rect 106410 572838 106465 572889
rect 106618 572838 106652 572928
rect 106720 572890 106778 572928
rect 106732 572838 106777 572890
rect 106848 572838 106893 572928
rect 107378 572890 107436 572928
rect 107494 572890 107572 572928
rect 107067 572878 107123 572889
rect 107078 572838 107123 572878
rect 107390 572838 107435 572890
rect 107504 572838 107572 572890
rect 107725 572878 107781 572889
rect 86640 572804 107614 572838
rect 86640 572774 106382 572804
rect 106410 572774 106465 572804
rect 106618 572774 106652 572804
rect 106732 572774 106777 572804
rect 106848 572774 106893 572804
rect 107078 572774 107123 572804
rect 107390 572774 107435 572804
rect 86640 572702 107476 572774
rect 86640 572222 106382 572702
rect 106408 572664 106466 572702
rect 106410 572356 106465 572664
rect 106490 572460 106548 572594
rect 106550 572460 106608 572594
rect 106410 572222 106454 572356
rect 106618 572222 106652 572702
rect 106732 572356 106777 572702
rect 106848 572356 106893 572702
rect 106732 572222 106766 572356
rect 106848 572222 106882 572356
rect 107078 572222 107123 572702
rect 107390 572222 107435 572702
rect 107504 572663 107572 572804
rect 107455 572652 107572 572663
rect 107466 572222 107572 572652
rect 107580 572222 107614 572804
rect 86640 571858 107676 572222
rect 86300 571548 107676 571858
rect 107736 571548 107781 572878
rect 86300 571410 107781 571548
rect 86640 571380 107781 571410
rect 107928 572228 107962 572928
rect 108030 572890 108088 572928
rect 108042 572356 108087 572890
rect 108164 572356 108209 572928
rect 108042 572228 108076 572356
rect 108164 572228 108198 572356
rect 108278 572228 108312 572928
rect 108383 572878 108439 572889
rect 108394 572356 108439 572878
rect 108394 572228 108428 572356
rect 108508 572228 108542 572992
rect 108694 572228 108696 572992
rect 108826 572228 108896 572992
rect 108942 572356 108962 573028
rect 108976 572322 108996 573028
rect 109060 572727 110086 573028
rect 110220 573274 113638 573310
rect 114092 573418 120428 573715
rect 120847 573703 120892 573714
rect 114092 573310 120417 573418
rect 120858 573310 120892 573703
rect 121041 573310 121075 573715
rect 121505 573703 121550 573714
rect 121516 573310 121550 573703
rect 121584 573310 121616 573864
rect 121630 573802 121664 573864
rect 121630 573310 121672 573802
rect 121699 573310 121733 573923
rect 121813 573518 121847 574354
rect 121882 573932 121883 574186
rect 123366 573932 123400 575148
rect 124138 574712 124172 576532
rect 124240 575920 127872 576576
rect 128264 576272 128274 576630
rect 128407 576611 129076 576749
rect 129244 576734 132730 576749
rect 129244 576700 132507 576734
rect 132650 576704 132674 576724
rect 132684 576704 132718 576734
rect 132650 576700 132718 576704
rect 129244 576676 132718 576700
rect 129244 576666 132507 576676
rect 132656 576672 132718 576676
rect 132650 576666 132718 576672
rect 129244 576632 132718 576666
rect 129094 576617 129122 576630
rect 129150 576617 129178 576630
rect 129244 576611 132507 576632
rect 132650 576626 132668 576632
rect 128407 576577 132507 576611
rect 132678 576598 132718 576632
rect 132678 576586 132680 576598
rect 128407 576529 129076 576577
rect 129122 576571 129150 576577
rect 128264 576058 128292 576272
rect 128264 576052 128274 576058
rect 124240 575850 127864 575920
rect 124208 574864 124230 575340
rect 124240 575216 126954 575850
rect 127016 575668 127020 575850
rect 127794 575668 127828 575850
rect 128407 575842 129078 576529
rect 129094 576528 129122 576571
rect 129150 576528 129178 576571
rect 129244 576529 132507 576577
rect 129204 576518 132507 576529
rect 132654 576528 132680 576586
rect 128443 575668 128477 575842
rect 128557 575668 128591 575702
rect 128919 575668 128953 575842
rect 129033 575668 129078 575842
rect 129215 576010 132507 576518
rect 132684 576048 132718 576598
rect 132656 576010 132718 576048
rect 129215 575976 132718 576010
rect 129215 575908 132507 575976
rect 132684 575908 132718 575976
rect 129215 575874 132730 575908
rect 132736 575874 132752 575908
rect 129215 575668 132507 575874
rect 127006 575634 132507 575668
rect 127006 575534 127040 575634
rect 127135 575566 127726 575613
rect 127058 575534 127062 575541
rect 127006 575478 127062 575534
rect 127182 575532 127726 575566
rect 127668 575485 127726 575532
rect 127794 575507 127828 575634
rect 127006 575216 127040 575478
rect 127056 575216 127062 575478
rect 127084 575216 127090 575478
rect 127109 575473 127165 575484
rect 127120 575216 127165 575473
rect 127680 575216 127725 575485
rect 127772 575216 127776 575485
rect 127794 575216 127846 575507
rect 128360 575484 128374 575526
rect 128402 575470 128416 575484
rect 128443 575473 128477 575634
rect 128919 575613 128953 575634
rect 129033 575613 129078 575634
rect 128545 575600 129080 575613
rect 128498 575532 128515 575566
rect 128545 575532 129100 575600
rect 128545 575485 128603 575532
rect 124138 574682 124178 574712
rect 124240 574700 127908 575216
rect 128372 575208 128374 575454
rect 128400 575208 128402 575426
rect 128436 575400 128477 575473
rect 128557 575400 128602 575485
rect 128408 575222 128752 575400
rect 128436 575208 128477 575222
rect 128557 575208 128602 575222
rect 128919 575208 128953 575532
rect 129021 575485 129079 575532
rect 129033 575208 129078 575485
rect 129083 575473 129139 575484
rect 124204 574684 127908 574700
rect 124198 574682 127908 574684
rect 124138 574064 124172 574682
rect 124204 574574 127908 574682
rect 124204 574444 124210 574574
rect 124240 574266 127908 574574
rect 128084 574485 129078 575208
rect 129094 574497 129139 575473
rect 129150 575144 129190 575340
rect 129150 574694 129162 575144
rect 129094 574485 129134 574490
rect 129150 574485 129162 574490
rect 128084 574472 129079 574485
rect 129094 574472 129122 574485
rect 128084 574404 129122 574472
rect 128084 574388 129079 574404
rect 128084 574336 129078 574388
rect 129094 574336 129122 574404
rect 129150 574336 129178 574485
rect 129208 574409 132507 575634
rect 129204 574398 132507 574409
rect 129208 574336 132507 574398
rect 128084 574302 132507 574336
rect 128084 574266 129078 574302
rect 124240 574064 127872 574266
rect 123468 574030 127872 574064
rect 124138 574000 124172 574030
rect 124240 574000 127872 574030
rect 123504 573996 127872 574000
rect 123502 573962 127872 573996
rect 123502 573932 123520 573962
rect 123530 573932 124178 573962
rect 122136 573518 122137 573932
rect 123330 573928 124178 573932
rect 122920 573532 122938 573708
rect 123330 573518 123786 573928
rect 124104 573922 124122 573928
rect 124132 573894 124178 573928
rect 124188 573928 127872 573962
rect 124188 573922 124206 573928
rect 121790 573494 123786 573518
rect 121813 573462 121847 573494
rect 122136 573462 122137 573494
rect 123330 573462 123786 573494
rect 121790 573438 123786 573462
rect 121813 573310 121847 573438
rect 122136 573310 122137 573438
rect 123330 573310 123786 573438
rect 110220 573240 113808 573274
rect 110220 573210 113638 573240
rect 110220 573138 113670 573210
rect 110220 573128 113638 573138
rect 110220 573112 113728 573128
rect 110220 573028 113638 573112
rect 113654 573099 113700 573100
rect 113649 573088 113700 573099
rect 113654 573084 113700 573088
rect 113648 573040 113649 573041
rect 113647 573039 113648 573040
rect 113654 573034 113656 573084
rect 113660 573028 113694 573084
rect 113774 573028 113808 573240
rect 110220 572994 113808 573028
rect 109060 572566 110052 572727
rect 110220 572668 113638 572994
rect 113647 572982 113648 572983
rect 113648 572981 113649 572982
rect 113654 572896 113656 572988
rect 110114 572634 113638 572668
rect 110220 572566 113638 572634
rect 107928 572192 108896 572228
rect 109020 572192 109040 572564
rect 109060 572532 113638 572566
rect 109060 572192 110052 572532
rect 110220 572494 113638 572532
rect 110220 572462 112450 572494
rect 113002 572462 113036 572494
rect 113660 572462 113694 572994
rect 113774 572462 113808 572994
rect 114092 572992 121883 573310
rect 114092 572462 117716 572992
rect 118076 572462 118110 572992
rect 118190 572462 118224 572992
rect 118228 572896 118246 572988
rect 118259 572462 121883 572992
rect 122136 573274 123786 573310
rect 122136 573240 123956 573274
rect 122136 573210 123786 573240
rect 122136 573138 123818 573210
rect 122136 572494 123786 573138
rect 123797 573088 123842 573099
rect 110220 572428 121883 572462
rect 110220 572370 112450 572428
rect 112936 572392 112996 572406
rect 113002 572388 113036 572428
rect 113042 572392 113102 572406
rect 113600 572392 113654 572406
rect 112884 572370 113538 572388
rect 113648 572382 113649 572383
rect 113647 572381 113648 572382
rect 113660 572370 113694 572428
rect 113774 572370 113808 572428
rect 114092 572370 117716 572428
rect 118076 572370 118110 572428
rect 118190 572370 118224 572428
rect 118228 572376 118230 572428
rect 118235 572382 118236 572383
rect 118236 572381 118237 572382
rect 118259 572370 121883 572428
rect 110220 572314 121883 572370
rect 107928 572158 110218 572192
rect 107928 572090 108896 572158
rect 108970 572156 109040 572158
rect 109060 572112 110052 572158
rect 110184 572112 110218 572158
rect 109038 572090 110218 572112
rect 107928 572078 110218 572090
rect 107928 572056 110052 572078
rect 107928 572010 108896 572056
rect 109060 572031 110052 572056
rect 109060 572010 110138 572031
rect 110184 572010 110218 572078
rect 110220 572010 112450 572314
rect 112920 572290 113574 572314
rect 107928 571976 112450 572010
rect 107928 571512 108884 571976
rect 109060 571800 110068 571976
rect 109060 571512 110052 571800
rect 107928 571478 110052 571512
rect 107928 571457 108884 571478
rect 107928 571416 108944 571457
rect 108946 571416 108993 571457
rect 107928 571380 109058 571416
rect 86640 571370 109058 571380
rect 109060 571370 110052 571478
rect 110064 571418 110068 571800
rect 110184 571620 110218 571976
rect 110220 571940 112450 571976
rect 110220 571620 110254 571940
rect 110256 571620 110290 571940
rect 110370 571792 110404 571940
rect 110370 571676 110410 571792
rect 110370 571656 110432 571676
rect 110370 571620 110404 571656
rect 110164 571600 110432 571620
rect 110070 571370 110096 571396
rect 86640 571366 110108 571370
rect 86640 571346 109058 571366
rect 86640 571277 107781 571346
rect 107844 571277 107868 571332
rect 86640 571266 107868 571277
rect 107878 571277 107902 571332
rect 107928 571314 109058 571346
rect 107946 571277 109058 571314
rect 109060 571362 110052 571366
rect 109060 571286 110062 571362
rect 107878 571266 109058 571277
rect 86640 571232 109058 571266
rect 86640 570910 107781 571232
rect 86640 570860 107676 570910
rect 86640 570819 107708 570860
rect 107736 570819 107781 570910
rect 107844 570819 107868 571232
rect 86640 570808 107868 570819
rect 107878 570819 107902 571232
rect 107946 570980 109058 571232
rect 109088 570980 109122 571286
rect 107946 570946 109122 570980
rect 109208 570980 109242 571286
rect 109322 571141 109367 571286
rect 109376 571272 109390 571286
rect 109412 571272 109446 571286
rect 109450 571272 109495 571286
rect 109564 571272 109598 571286
rect 109348 571129 109362 571141
rect 109376 571129 109728 571272
rect 109337 571094 109728 571129
rect 109337 571082 109474 571094
rect 109384 571072 109474 571082
rect 109358 571016 109474 571072
rect 109358 571009 109458 571016
rect 109358 571008 109448 571009
rect 109350 570994 109462 570996
rect 109564 570980 109598 571094
rect 109208 570969 109411 570980
rect 109447 570969 109598 570980
rect 109208 570968 109400 570969
rect 109458 570968 109598 570969
rect 109988 570968 110012 571002
rect 110036 570974 110062 571286
rect 110070 571005 110096 571366
rect 110016 570971 110062 570974
rect 110016 570968 110040 570971
rect 109208 570966 109598 570968
rect 109208 570957 109400 570966
rect 109458 570957 109598 570966
rect 109208 570946 109411 570957
rect 109447 570946 109598 570957
rect 107946 570896 109058 570946
rect 110184 570922 110218 571600
rect 107946 570819 109136 570896
rect 107878 570808 109136 570819
rect 86640 570790 109136 570808
rect 109190 570790 109612 570896
rect 110220 570790 110254 571600
rect 86640 570774 108576 570790
rect 108584 570786 108642 570790
rect 108716 570774 108818 570790
rect 86219 570534 86264 570724
rect 85834 570502 86264 570534
rect 86640 570694 97688 570774
rect 97785 570724 106386 570774
rect 106410 570724 106454 570774
rect 97785 570694 106382 570724
rect 106410 570694 106465 570724
rect 106848 570694 106916 570774
rect 107002 570760 107392 570774
rect 107002 570758 107123 570760
rect 107034 570738 107123 570758
rect 107040 570724 107123 570738
rect 107078 570708 107123 570724
rect 106962 570694 107064 570708
rect 107078 570694 107152 570708
rect 107198 570694 107232 570760
rect 107358 570694 107392 570760
rect 107482 570758 107588 570774
rect 107506 570724 107588 570758
rect 107506 570708 107551 570724
rect 107438 570694 107628 570708
rect 107674 570694 107708 570774
rect 107736 570694 107781 570774
rect 107844 570724 107868 570774
rect 107878 570724 107902 570774
rect 108164 570694 108209 570774
rect 108278 570694 108312 570774
rect 108320 570698 108334 570768
rect 108348 570712 108390 570768
rect 108388 570698 108390 570712
rect 108320 570694 108388 570698
rect 108394 570694 108428 570774
rect 108508 570754 108542 570774
rect 108434 570712 108548 570754
rect 108508 570698 108542 570712
rect 108434 570694 108576 570698
rect 108750 570694 108784 570774
rect 108832 570768 108848 570790
rect 108858 570724 108890 570790
rect 108892 570724 108924 570758
rect 108954 570756 108958 570758
rect 108988 570756 109022 570790
rect 108940 570724 108942 570741
rect 108988 570724 108989 570756
rect 108830 570694 108932 570708
rect 86640 570686 108951 570694
rect 86640 570660 108998 570686
rect 109016 570660 109022 570756
rect 85834 570500 86253 570502
rect 85834 570002 85868 570500
rect 86037 570479 86071 570500
rect 86037 570432 86084 570479
rect 86010 570398 86084 570432
rect 86037 570350 86071 570398
rect 86076 570350 86105 570355
rect 85937 570339 85982 570350
rect 85948 570163 85982 570339
rect 86037 570339 86110 570350
rect 86114 570346 86142 570500
rect 86170 570346 86253 570500
rect 86037 570151 86071 570339
rect 86076 570163 86110 570339
rect 86076 570151 86105 570163
rect 86037 570147 86105 570151
rect 86190 570150 86253 570346
rect 86037 570104 86084 570147
rect 86010 570070 86084 570104
rect 86037 570002 86071 570070
rect 86114 570002 86142 570150
rect 86170 570002 86253 570150
rect 85834 569968 86253 570002
rect 86037 569918 86071 569968
rect 86114 569918 86142 569968
rect 86170 569918 86198 569968
rect 86219 569918 86253 569968
rect 85820 569374 86253 569918
rect 86640 570344 97688 570660
rect 97785 570624 106382 570660
rect 97785 570616 102756 570624
rect 97762 570344 102756 570616
rect 86640 570272 102756 570344
rect 86640 570204 97688 570272
rect 97762 570204 102756 570272
rect 86640 570181 102756 570204
rect 102794 570181 102828 570624
rect 102856 570572 106382 570624
rect 106410 570572 106465 570660
rect 106848 570600 106916 570660
rect 106996 570600 107041 570660
rect 107078 570600 107129 570660
rect 107198 570600 107232 570660
rect 107358 570600 107392 570660
rect 107472 570600 107551 570660
rect 106618 570572 107551 570600
rect 107560 570572 107605 570660
rect 107674 570572 107708 570660
rect 107736 570572 107781 570660
rect 108164 570608 108209 570660
rect 108278 570608 108312 570660
rect 108394 570608 108428 570660
rect 108508 570608 108542 570660
rect 108750 570608 108784 570660
rect 107928 570574 108784 570608
rect 108827 570574 108848 570608
rect 107928 570572 107962 570574
rect 108164 570572 108209 570574
rect 108278 570572 108312 570574
rect 108394 570572 108428 570574
rect 102856 570506 108462 570572
rect 108508 570506 108542 570574
rect 102856 570472 108672 570506
rect 102856 570280 108462 570472
rect 108508 570280 108542 570472
rect 102856 570194 108542 570280
rect 102856 570181 108462 570194
rect 86640 570170 108462 570181
rect 86640 570134 97685 570170
rect 86640 570111 96492 570134
rect 86640 569802 91268 570111
rect 85820 569298 86264 569374
rect 86037 569156 86082 569298
rect 86037 567688 86071 569156
rect 86114 567635 86142 569298
rect 86170 567635 86198 569298
rect 86219 569156 86264 569298
rect 86219 567688 86253 569156
rect 86640 568614 91261 569802
rect 86640 568311 91268 568614
rect 86640 567629 87537 568311
rect 85123 567595 87537 567629
rect 84351 567527 84385 567561
rect 85009 567527 85043 567561
rect 85123 567527 85157 567595
rect 85444 567582 85472 567589
rect 85500 567582 85528 567589
rect 86114 567582 86142 567589
rect 86170 567582 86198 567589
rect 86640 567527 87537 567595
rect 83473 567493 87537 567527
rect 83035 567338 83069 567372
rect 82368 567304 82758 567338
rect 82368 567276 82402 567304
rect 82368 566868 82436 567276
rect 82582 567236 82629 567283
rect 82544 567202 82629 567236
rect 82471 567143 82516 567154
rect 82599 567143 82644 567154
rect 82482 566967 82516 567143
rect 82610 566967 82644 567143
rect 82582 566908 82629 566955
rect 82544 566874 82629 566908
rect 82368 566806 82402 566868
rect 82724 566806 82758 567304
rect 82368 566772 82758 566806
rect 82844 567304 83234 567338
rect 82844 566806 82878 567304
rect 83035 567270 83082 567283
rect 83035 567258 83092 567270
rect 83014 567202 83092 567258
rect 82924 567150 82942 567183
rect 83014 567159 83088 567202
rect 83014 567155 83103 567159
rect 82952 567154 82970 567155
rect 83014 567154 83116 567155
rect 82947 567143 82992 567154
rect 82958 566967 82992 567143
rect 83014 567148 83120 567154
rect 83014 567144 83126 567148
rect 83014 566967 83120 567144
rect 83014 566964 83116 566967
rect 83014 566955 83126 566964
rect 82966 566954 82992 566955
rect 82994 566951 83103 566955
rect 82994 566942 83088 566951
rect 82994 566926 83092 566942
rect 83014 566898 83092 566926
rect 82994 566874 83092 566898
rect 82994 566834 83088 566874
rect 82978 566820 82994 566822
rect 83014 566806 83088 566834
rect 83100 566806 83102 566951
rect 83200 566806 83234 567304
rect 82844 566772 83234 566806
rect 83014 566722 83088 566772
rect 81685 566138 81708 566212
rect 81713 566110 81736 566212
rect 82350 566102 82772 566722
rect 82826 566102 83248 566722
rect 81685 565848 81708 565970
rect 81713 565876 81736 565998
rect 85123 565789 85157 567493
rect 86640 567457 87537 567493
rect 87637 568002 91268 568311
rect 91290 568214 91335 570111
rect 91766 568214 91811 570111
rect 91836 569802 91864 570111
rect 91866 570070 96492 570111
rect 91866 569932 96442 570070
rect 96458 570002 96492 570070
rect 96558 570002 97685 570134
rect 96458 569968 97685 570002
rect 91892 569802 91920 569932
rect 91948 569882 91993 569932
rect 92062 569882 92096 569932
rect 92193 569882 96442 569932
rect 96558 569918 97685 569968
rect 91924 569848 96442 569882
rect 91924 569368 91993 569848
rect 92062 569818 92096 569848
rect 92062 569746 92154 569818
rect 92062 569707 92096 569746
rect 92193 569718 96442 569848
rect 96444 569718 97685 569918
rect 92027 569696 92096 569707
rect 92115 569696 92171 569707
rect 92038 569520 92096 569696
rect 92126 569520 92171 569696
rect 92193 569668 97685 569718
rect 97762 570147 108462 570170
rect 97762 570111 102756 570147
rect 97762 569690 101409 570111
rect 97752 569682 101409 569690
rect 92193 569658 96442 569668
rect 96444 569658 97685 569668
rect 92193 569576 97685 569658
rect 92062 569508 92096 569520
rect 92062 569436 92154 569508
rect 92062 569368 92096 569436
rect 92193 569368 96442 569576
rect 91924 569334 96442 569368
rect 87637 567652 91261 568002
rect 91290 567702 91324 568214
rect 91766 567702 91800 568214
rect 91836 568002 91864 568614
rect 91892 568002 91920 568614
rect 91948 568214 91993 569334
rect 91948 567702 91982 568214
rect 92062 567652 92096 569334
rect 92193 569329 96442 569334
rect 96444 569329 97685 569576
rect 92193 569298 97685 569329
rect 92193 569248 96504 569298
rect 92193 569180 96460 569248
rect 96476 569214 96504 569248
rect 96476 569180 96494 569214
rect 96558 569180 97685 569298
rect 92193 569146 97685 569180
rect 92193 569096 96442 569146
rect 96558 569096 97685 569146
rect 92193 568624 97685 569096
rect 97762 568894 101409 569682
rect 101668 568894 101713 570111
rect 101914 569150 101959 570111
rect 102326 569702 102371 570111
rect 102292 569560 102318 569702
rect 102326 569560 102360 569702
rect 101876 569036 102068 569150
rect 102326 569048 102371 569560
rect 101896 568894 101970 569036
rect 97762 568826 102174 568894
rect 97762 568668 101702 568826
rect 92193 568476 96644 568624
rect 96698 568476 97120 568624
rect 97174 568476 97685 568624
rect 92193 568334 96332 568476
rect 92193 568326 92608 568334
rect 92708 568326 96332 568334
rect 92193 568292 96332 568326
rect 92193 568242 92608 568292
rect 92708 568242 96332 568292
rect 96750 568278 96766 568476
rect 96822 568458 96968 568476
rect 96822 568394 96915 568458
rect 96822 568384 96896 568394
rect 96844 568356 96877 568384
rect 92193 567652 96332 568242
rect 87637 567618 96332 567652
rect 87637 567550 91261 567618
rect 92062 567602 92096 567618
rect 92062 567591 92073 567602
rect 92085 567591 92096 567602
rect 92193 567612 96332 567618
rect 97264 567652 97685 568476
rect 97785 568311 101702 568668
rect 98072 567690 98106 568311
rect 98696 567690 98728 568311
rect 98730 567690 98764 568311
rect 97716 567652 98764 567690
rect 98922 567690 98956 568311
rect 99036 567690 99070 568311
rect 99168 567690 99202 568311
rect 99282 567702 99316 568311
rect 99388 567690 99422 568311
rect 98922 567652 98960 567690
rect 99036 567652 99074 567690
rect 99168 567652 99206 567690
rect 99388 567652 99426 567690
rect 99694 567652 99728 568311
rect 99940 567702 99974 568311
rect 100046 567690 100080 568311
rect 100046 567652 100084 567690
rect 100352 567652 100386 568311
rect 100598 567702 100632 568311
rect 100704 567690 100738 568311
rect 100704 567652 100742 567690
rect 100818 567652 100852 568311
rect 101010 567698 101044 568311
rect 101236 568256 101702 568311
rect 101712 568256 102174 568826
rect 101256 568206 101290 568256
rect 101256 568172 101640 568206
rect 101256 567702 101324 568172
rect 101482 568104 101520 568142
rect 101448 568070 101520 568104
rect 101393 568020 101438 568031
rect 101481 568020 101526 568031
rect 101404 567844 101438 568020
rect 101492 567844 101526 568020
rect 101482 567794 101520 567832
rect 101448 567760 101520 567794
rect 101010 567690 101055 567698
rect 101290 567692 101324 567702
rect 101606 567692 101640 568172
rect 101290 567690 101640 567692
rect 101668 567698 101702 568256
rect 101914 568206 101948 568256
rect 101766 568172 102116 568206
rect 101668 567690 101713 567698
rect 101766 567692 101800 568172
rect 101914 568138 101948 568172
rect 101890 568104 101948 568138
rect 101958 568104 101996 568142
rect 101914 568070 101996 568104
rect 101914 568031 101948 568070
rect 101968 568031 101982 568036
rect 101869 568020 101948 568031
rect 101957 568020 102002 568031
rect 101880 567844 101948 568020
rect 101914 567828 101948 567844
rect 101968 567844 102002 568020
rect 101968 567832 101982 567844
rect 101890 567794 101948 567828
rect 101958 567794 101996 567832
rect 101914 567760 101996 567794
rect 101914 567702 101948 567760
rect 102082 567692 102116 568172
rect 101766 567690 102116 567692
rect 102326 567690 102360 569048
rect 100906 567652 101266 567690
rect 101280 567658 102120 567690
rect 101280 567652 101924 567658
rect 101938 567652 102120 567658
rect 102314 567652 102372 567690
rect 97264 567618 98106 567652
rect 98134 567618 98764 567652
rect 98776 567618 101266 567652
rect 101318 567618 101924 567652
rect 101976 567618 102372 567652
rect 92193 567595 96358 567612
rect 92193 567550 92608 567595
rect 87637 567527 92608 567550
rect 92708 567527 96332 567595
rect 87637 567516 96332 567527
rect 87637 567480 91261 567516
rect 92193 567493 96332 567516
rect 92193 567480 92608 567493
rect 87637 565829 90264 567480
rect 90381 567068 90402 567150
rect 90419 567030 90440 567188
rect 91070 567058 91123 567112
rect 91191 567058 91225 567480
rect 92708 567457 96332 567493
rect 97264 567550 97685 567618
rect 98072 567550 98106 567618
rect 98696 567554 98728 567618
rect 98730 567550 98764 567618
rect 98922 567550 98956 567618
rect 99036 567554 99070 567618
rect 99036 567550 99081 567554
rect 99168 567550 99202 567618
rect 99388 567554 99422 567618
rect 99694 567554 99728 567618
rect 100046 567554 100080 567618
rect 100352 567554 100386 567618
rect 100704 567554 100738 567618
rect 99388 567550 99433 567554
rect 99694 567550 99739 567554
rect 100046 567550 100091 567554
rect 100352 567550 100397 567554
rect 100704 567550 100749 567554
rect 100818 567550 100852 567618
rect 100998 567602 101056 567618
rect 101656 567602 101714 567618
rect 102314 567602 102372 567618
rect 102357 567587 102372 567602
rect 102440 567550 102474 570111
rect 102578 569560 102606 569702
rect 102612 569560 102640 569702
rect 102794 569628 102828 570147
rect 102856 569876 108462 570147
rect 102856 569550 106382 569876
rect 106410 569702 106454 569876
rect 106410 569550 106444 569702
rect 106482 569618 106491 569652
rect 106618 569550 106652 569876
rect 106732 569690 106777 569876
rect 107078 569804 107123 569876
rect 107052 569748 107123 569804
rect 107390 569748 107435 569876
rect 107504 569748 107538 569876
rect 107736 569748 107770 569876
rect 106828 569690 107290 569748
rect 107304 569702 107770 569748
rect 107304 569690 107766 569702
rect 106720 569618 107766 569690
rect 106720 569602 106778 569618
rect 106720 569587 106766 569602
rect 106732 569550 106766 569587
rect 106828 569550 107290 569618
rect 107304 569550 107766 569618
rect 107928 569550 107962 569876
rect 108042 569690 108087 569876
rect 108374 569772 108462 569876
rect 108322 569696 108472 569772
rect 108030 569630 108404 569690
rect 107980 569618 108404 569630
rect 107980 569612 108088 569618
rect 108030 569602 108088 569612
rect 108030 569587 108045 569602
rect 107980 569556 108036 569574
rect 108042 569550 108076 569584
rect 108082 569556 108136 569574
rect 108508 569550 108542 570194
rect 108694 569638 108704 570434
rect 108725 570312 108746 570434
rect 108750 570346 108784 570574
rect 108814 570346 108848 570574
rect 108852 570486 108902 570660
rect 109050 570626 109056 570790
rect 109066 570764 109076 570790
rect 109066 570520 109100 570764
rect 109226 570616 109260 570764
rect 109340 570616 109374 570650
rect 109428 570616 109462 570650
rect 109542 570616 109576 570764
rect 109192 570582 109920 570616
rect 109066 570408 109130 570520
rect 108750 570312 108800 570346
rect 108814 570312 109004 570346
rect 108694 569612 108696 569638
rect 102856 569516 108542 569550
rect 102856 569496 106382 569516
rect 103664 568894 103698 569496
rect 105428 569286 105462 569496
rect 105542 569438 105587 569496
rect 105620 569426 105694 569496
rect 106200 569438 106245 569496
rect 105566 569388 106210 569426
rect 105604 569354 106210 569388
rect 105620 569286 105694 569354
rect 106314 569348 106364 569496
rect 106314 569286 106342 569348
rect 105428 569252 106342 569286
rect 105620 569238 105694 569252
rect 102586 568474 102612 568614
rect 103104 568466 103566 568894
rect 103580 568466 104042 568894
rect 105660 568746 105672 569094
rect 105698 568784 105710 569056
rect 103104 568460 104042 568466
rect 102764 568258 102780 568360
rect 103104 568334 103566 568460
rect 103580 568334 104042 568460
rect 106376 568408 106386 569048
rect 106410 568466 106444 569516
rect 106618 569348 106652 569516
rect 106732 569438 106766 569516
rect 106828 569388 107290 569516
rect 107304 569480 107766 569516
rect 107304 569388 107574 569480
rect 106828 569354 107574 569388
rect 106828 569216 107290 569354
rect 107304 569216 107574 569354
rect 107304 569110 107544 569216
rect 106882 568814 107264 569052
rect 106996 568698 107030 568814
rect 107084 568698 107118 568814
rect 107928 568756 107962 569516
rect 108036 569256 108046 569364
rect 108814 568756 108848 570312
rect 109096 568764 109130 570408
rect 109226 570346 109260 570582
rect 109328 570486 109474 570552
rect 109346 570480 109456 570486
rect 109384 570442 109418 570448
rect 109384 570414 109456 570442
rect 109542 570388 109576 570582
rect 109542 570368 109798 570388
rect 109542 570346 109576 570368
rect 109226 570312 109576 570346
rect 109594 570183 109595 570368
rect 109778 570183 109798 570368
rect 109594 570182 109798 570183
rect 106410 568408 106420 568466
rect 102792 568258 102808 568332
rect 103268 568312 103422 568332
rect 103580 568314 103820 568334
rect 103580 568312 103898 568314
rect 103580 568256 103820 568312
rect 102780 568058 102956 568084
rect 103312 568062 103354 568084
rect 107844 568044 107868 568738
rect 107878 568044 107902 568704
rect 102586 568002 102612 568028
rect 103830 568020 103844 568028
rect 103748 567844 103782 568020
rect 103830 568002 103870 568020
rect 103836 567844 103870 568002
rect 97264 567516 102624 567550
rect 97264 567457 97685 567516
rect 90648 567024 91038 567058
rect 90648 566526 90682 567024
rect 90777 566956 90909 567003
rect 90824 566922 90909 566956
rect 90751 566863 90807 566874
rect 90879 566863 90935 566874
rect 90762 566687 90807 566863
rect 90890 566687 90935 566863
rect 90777 566662 90909 566675
rect 90777 566642 90912 566662
rect 90777 566628 90909 566642
rect 90824 566594 90909 566628
rect 91004 566526 91038 567024
rect 91099 566996 91123 567058
rect 91090 566962 91123 566996
rect 91099 566642 91123 566962
rect 90648 566492 91038 566526
rect 91090 566492 91123 566642
rect 91124 567024 91177 567058
rect 91191 567024 91418 567058
rect 91124 566526 91158 567024
rect 91191 566526 91225 567024
rect 91226 566675 91279 566875
rect 91250 566642 91388 566662
rect 91284 566608 91354 566628
rect 91124 566492 91177 566526
rect 91191 566492 91418 566526
rect 91090 566460 91111 566492
rect 91088 566442 91123 566460
rect 91191 566442 91225 566492
rect 90630 565829 91052 566442
rect 91088 566406 91261 566442
rect 87510 565826 90391 565829
rect 87510 565818 90424 565826
rect 87637 565795 90424 565818
rect 90481 565822 91052 565829
rect 91106 566232 91261 566406
rect 91106 566032 91279 566232
rect 91106 565822 91261 566032
rect 90481 565795 91049 565822
rect 87637 565680 90264 565795
rect 91191 565789 91225 565822
rect 92708 565680 95817 567457
rect 96228 567116 96250 567457
rect 96262 567116 96284 567457
rect 97156 566456 97618 567094
rect 97300 566406 97334 566456
rect 97414 566406 97448 566440
rect 97300 566372 97560 566406
rect 97300 566220 97334 566372
rect 97414 566342 97448 566372
rect 97402 566304 97448 566342
rect 97352 566270 97448 566304
rect 97402 566232 97448 566270
rect 97414 566220 97448 566232
rect 97312 566044 97334 566220
rect 97412 566044 97448 566220
rect 97022 565680 97032 565960
rect 97050 565652 97060 565960
rect 97300 565892 97334 566044
rect 97414 566032 97448 566044
rect 97402 565994 97448 566032
rect 97352 565960 97448 565994
rect 97402 565929 97448 565960
rect 97414 565902 97448 565929
rect 97526 565892 97560 566372
rect 98072 565902 98106 567516
rect 98922 567106 98956 567516
rect 99036 567258 99081 567516
rect 99388 567246 99433 567516
rect 99694 567258 99739 567516
rect 100046 567246 100091 567516
rect 100352 567258 100397 567516
rect 100704 567246 100749 567516
rect 99060 567208 99704 567246
rect 99718 567208 100362 567246
rect 100376 567208 100750 567246
rect 99098 567174 99704 567208
rect 99756 567174 100362 567208
rect 100414 567174 100750 567208
rect 99376 567158 99434 567174
rect 100034 567158 100092 567174
rect 100692 567158 100750 567174
rect 99388 567106 99422 567140
rect 100046 567106 100080 567158
rect 100704 567143 100750 567158
rect 100704 567106 100738 567143
rect 100818 567106 100852 567516
rect 101010 567486 101044 567516
rect 100902 567174 100982 567188
rect 101378 567174 101540 567188
rect 102440 567168 102474 567516
rect 110256 567168 110290 571600
rect 110370 571474 110404 571600
rect 110370 570620 110410 571474
rect 111680 570620 111704 571940
rect 112016 571598 112050 571940
rect 112118 571718 112152 571940
rect 112344 571712 112378 571940
rect 113002 571712 113036 572290
rect 113660 571712 113694 572314
rect 113774 571712 113808 572314
rect 114092 572222 117716 572314
rect 118076 572228 118110 572314
rect 118190 572228 118224 572314
rect 118228 572244 118230 572308
rect 118259 572228 121883 572314
rect 114092 571712 117824 572222
rect 118076 571712 121883 572228
rect 112080 571628 112152 571666
rect 112202 571656 121883 571712
rect 112331 571644 112332 571645
rect 112332 571643 112333 571644
rect 112118 571602 112152 571628
rect 112080 571598 112152 571602
rect 112344 571598 112378 571656
rect 112390 571644 112391 571645
rect 112989 571644 112990 571645
rect 112389 571643 112390 571644
rect 112990 571643 112991 571644
rect 113002 571598 113036 571656
rect 113048 571644 113049 571645
rect 113647 571644 113648 571645
rect 113047 571643 113048 571644
rect 113648 571643 113649 571644
rect 113660 571598 113694 571656
rect 113774 571598 113808 571656
rect 114092 571598 117824 571656
rect 118076 571598 121883 571656
rect 112016 571564 121883 571598
rect 112016 571454 112050 571564
rect 112118 571510 112152 571564
rect 112118 571454 112190 571510
rect 112016 571368 112190 571454
rect 112016 570970 112050 571368
rect 112118 571126 112190 571368
rect 112344 571126 112378 571564
rect 113002 571180 113036 571564
rect 112118 571092 112706 571126
rect 112118 571060 112192 571092
rect 112158 571008 112192 571060
rect 112332 571044 112333 571045
rect 112331 571043 112332 571044
rect 112344 571032 112378 571092
rect 112672 571064 112706 571092
rect 112389 571044 112390 571045
rect 112390 571043 112391 571044
rect 112638 571032 112740 571064
rect 112756 571050 113394 571180
rect 113600 571116 113654 571130
rect 113654 571074 113656 571116
rect 112756 571043 113546 571050
rect 113648 571044 113649 571045
rect 113647 571043 113648 571044
rect 112756 571032 113548 571043
rect 113660 571032 113694 571564
rect 113774 571032 113808 571564
rect 112080 570970 112192 571008
rect 112202 570998 113808 571032
rect 112016 570892 112192 570970
rect 112222 570968 112294 570998
rect 112331 570986 112332 570987
rect 112332 570985 112333 570986
rect 112260 570934 112294 570968
rect 112344 570978 112531 570998
rect 112016 570620 112050 570892
rect 112118 570810 112192 570892
rect 112344 570924 112378 570978
rect 112532 570968 112604 570998
rect 112520 570924 112531 570935
rect 112570 570934 112604 570968
rect 112344 570890 112531 570924
rect 112344 570810 112378 570890
rect 112672 570810 112706 570998
rect 112118 570776 112706 570810
rect 112756 570976 113546 570998
rect 113647 570986 113648 570987
rect 113648 570985 113649 570986
rect 112118 570650 112190 570776
rect 112344 570650 112378 570776
rect 112756 570718 113394 570976
rect 113654 570906 113656 570966
rect 113002 570704 113036 570718
rect 112118 570624 112706 570650
rect 112080 570620 112706 570624
rect 112756 570620 113394 570704
rect 113660 570620 113694 570998
rect 113774 570620 113808 570998
rect 110358 570586 113808 570620
rect 110370 570580 110410 570586
rect 110364 570524 110410 570580
rect 111028 570556 111062 570586
rect 111680 570580 111720 570586
rect 111680 570556 111726 570580
rect 112016 570556 112050 570586
rect 112118 570556 112192 570586
rect 112344 570556 112378 570586
rect 112672 570556 112706 570586
rect 112756 570556 113394 570586
rect 113660 570556 113694 570586
rect 110370 570478 110410 570524
rect 110420 570518 110438 570524
rect 111000 570518 111062 570556
rect 111142 570518 112198 570556
rect 112316 570552 112378 570556
rect 112482 570552 112536 570556
rect 112316 570536 112536 570552
rect 112298 570518 112536 570536
rect 112672 570518 112710 570556
rect 112756 570518 113548 570556
rect 113632 570518 113694 570556
rect 110416 570484 111062 570518
rect 111074 570484 111726 570518
rect 110420 570478 110438 570484
rect 110364 570440 110410 570478
rect 110370 570380 110436 570440
rect 110460 570380 110464 570468
rect 110370 570180 110404 570380
rect 110370 570034 110436 570180
rect 110370 569924 110410 570034
rect 110460 570006 110464 570180
rect 110364 569868 110410 569924
rect 111028 569900 111062 570484
rect 111652 570478 111670 570484
rect 111680 570422 111726 570484
rect 111736 570502 113694 570518
rect 111736 570484 112378 570502
rect 112390 570484 113694 570502
rect 111736 570478 111754 570484
rect 111686 570094 111720 570422
rect 111680 569924 111720 570094
rect 111680 569900 111726 569924
rect 112016 569900 112050 570484
rect 112118 570402 112192 570484
rect 112260 570458 112294 570484
rect 112304 570458 112338 570482
rect 112332 570408 112338 570454
rect 112344 570448 112378 570484
rect 112384 570458 112438 570482
rect 112384 570448 112438 570454
rect 112520 570448 112531 570459
rect 112570 570458 112604 570484
rect 112344 570414 112531 570448
rect 112158 570350 112192 570402
rect 112332 570386 112333 570387
rect 112331 570385 112332 570386
rect 112344 570374 112378 570414
rect 112384 570402 112438 570414
rect 112389 570386 112390 570387
rect 112390 570385 112391 570386
rect 112672 570374 112706 570484
rect 112756 570385 113394 570484
rect 113648 570386 113649 570387
rect 113647 570385 113648 570386
rect 112756 570374 113548 570385
rect 113654 570380 113656 570432
rect 113660 570374 113694 570484
rect 113774 570374 113808 570586
rect 112202 570368 113808 570374
rect 112080 570334 112192 570350
rect 112198 570340 113808 570368
rect 112344 570334 112378 570340
rect 112672 570334 112706 570340
rect 112080 570312 112706 570334
rect 112118 570300 112706 570312
rect 112118 570296 112190 570300
rect 110370 569822 110410 569868
rect 110420 569862 110438 569868
rect 111000 569862 111062 569900
rect 111142 569862 112054 569900
rect 112118 569862 112152 570296
rect 112344 569900 112378 570300
rect 112756 570242 113394 570340
rect 113647 570328 113648 570329
rect 113648 570327 113649 570328
rect 113654 570242 113656 570334
rect 113002 569900 113036 570242
rect 113660 569900 113694 570340
rect 112316 569862 112378 569900
rect 112974 569862 113036 569900
rect 113632 569862 113694 569900
rect 110416 569828 111062 569862
rect 111074 569828 111726 569862
rect 110420 569822 110438 569828
rect 110364 569766 110410 569822
rect 110370 569760 110410 569766
rect 111028 569760 111062 569828
rect 111652 569822 111670 569828
rect 111680 569766 111726 569828
rect 111736 569828 112378 569862
rect 112390 569828 113036 569862
rect 113048 569828 113694 569862
rect 111736 569822 111754 569828
rect 111680 569760 111720 569766
rect 112016 569760 112050 569828
rect 112118 569770 112152 569828
rect 112344 569770 112378 569828
rect 113002 569770 113036 569828
rect 113660 569770 113694 569828
rect 112118 569760 112190 569770
rect 112344 569760 112389 569770
rect 113002 569760 113047 569770
rect 113660 569760 113705 569770
rect 113774 569760 113808 570340
rect 110352 569726 113808 569760
rect 110404 568930 110410 569726
rect 111082 569258 111126 569274
rect 111116 569232 111126 569240
rect 111088 568986 111102 569232
rect 111116 568930 111158 569232
rect 111680 569186 111704 569726
rect 112016 568944 112050 569726
rect 112191 569716 112332 569726
rect 112344 569716 112378 569726
rect 112390 569716 112990 569726
rect 113002 569716 113036 569726
rect 113048 569716 113648 569726
rect 113660 569716 113694 569726
rect 113774 569716 113808 569726
rect 114092 570784 117824 571564
rect 118076 571426 121883 571564
rect 118040 571416 121883 571426
rect 118076 571314 121883 571416
rect 118094 570790 121883 571314
rect 114092 570374 117716 570784
rect 118259 570620 121883 570790
rect 122492 570620 122526 572494
rect 122546 572028 122580 572494
rect 122666 572434 122776 572472
rect 122704 572400 122776 572434
rect 122649 572350 122705 572361
rect 122737 572350 122793 572361
rect 122660 572174 122705 572350
rect 122748 572174 122793 572350
rect 122666 572124 122776 572162
rect 122704 572090 122776 572124
rect 122542 572022 122580 572028
rect 122862 572022 122896 572494
rect 123058 572358 123084 572462
rect 123114 572358 123140 572462
rect 122542 571988 122896 572022
rect 122542 571810 122560 571988
rect 123058 571006 123084 571810
rect 123114 571006 123140 571810
rect 123150 571006 123184 572494
rect 123366 571006 123400 572494
rect 123480 571006 123525 572494
rect 123808 571870 123842 573088
rect 123922 571870 123956 573240
rect 124094 572360 124116 573234
rect 124138 572058 124172 573894
rect 124240 573828 127872 573928
rect 124240 573782 127964 573828
rect 128264 573792 128274 574266
rect 128407 574059 129078 574266
rect 129094 574059 129122 574302
rect 129150 574059 129178 574302
rect 129215 574059 132507 574302
rect 128407 574025 132507 574059
rect 128407 574004 129078 574025
rect 129094 574004 129122 574025
rect 128407 573991 129122 574004
rect 129150 574004 129178 574025
rect 129215 574004 132507 574025
rect 132650 574022 132674 575128
rect 129150 574000 132507 574004
rect 129150 573991 132662 574000
rect 128407 573923 132662 573991
rect 128407 573922 129078 573923
rect 128407 573917 129150 573922
rect 128407 573907 129122 573917
rect 129150 573907 129178 573917
rect 129215 573907 132662 573923
rect 128407 573860 132662 573907
rect 128407 573792 129122 573860
rect 129126 573826 132662 573860
rect 129126 573820 129178 573826
rect 128056 573782 129122 573792
rect 124240 573772 127872 573782
rect 124240 573754 127908 573772
rect 128264 573764 128274 573782
rect 128407 573776 129122 573782
rect 129150 573776 129178 573820
rect 128407 573764 129140 573776
rect 128084 573754 129140 573764
rect 124240 573502 127872 573754
rect 128264 573618 128274 573754
rect 128264 573502 128292 573618
rect 128407 573536 129140 573754
rect 129150 573536 129168 573776
rect 124208 572210 124230 573314
rect 124240 573196 127908 573502
rect 124240 572742 126964 573196
rect 126972 573014 127020 573196
rect 127022 573014 127056 573196
rect 127538 573014 127572 573196
rect 127600 573014 127614 573196
rect 127628 573014 127670 573196
rect 127680 573014 127714 573196
rect 127794 573102 127828 573196
rect 128084 573188 128380 573502
rect 128407 573188 129122 573536
rect 129150 573480 129196 573536
rect 129150 573264 129178 573480
rect 129215 573356 132662 573826
rect 132678 573394 132680 575340
rect 132684 573988 132708 575162
rect 132684 573390 132718 573412
rect 132674 573356 132752 573378
rect 129215 573322 132672 573356
rect 127744 573074 127964 573102
rect 127744 573056 127864 573074
rect 127744 573040 127920 573056
rect 127794 573014 127828 573040
rect 127864 573038 127920 573040
rect 128310 573014 128344 573182
rect 128407 573050 128634 573188
rect 128443 573014 128477 573050
rect 128919 573014 128953 573188
rect 128962 573014 128996 573188
rect 129033 573014 129067 573188
rect 129076 573014 129122 573188
rect 129215 573242 132662 573322
rect 132674 573288 132706 573356
rect 132798 573316 132832 579068
rect 134239 579032 137863 579068
rect 138526 579052 138560 579068
rect 138842 579052 138876 579068
rect 134275 576962 134309 579032
rect 133248 576928 136704 576962
rect 133152 573478 133186 576866
rect 133232 576724 133252 576817
rect 133266 576690 133286 576783
rect 133924 576779 133958 576783
rect 133918 576754 133958 576779
rect 133960 576754 133964 576779
rect 134275 576754 134309 576928
rect 134389 576891 134436 576907
rect 134377 576860 134436 576891
rect 134554 576860 134601 576907
rect 135047 576876 135094 576907
rect 135035 576860 135094 576876
rect 135212 576860 135259 576907
rect 135705 576876 135752 576907
rect 135693 576860 135752 576876
rect 135870 576860 135917 576907
rect 136363 576876 136410 576907
rect 136351 576860 136410 576876
rect 136528 576860 136575 576907
rect 134377 576826 134601 576860
rect 134644 576826 135259 576860
rect 135302 576826 135917 576860
rect 135960 576826 136575 576860
rect 134377 576779 134435 576826
rect 134389 576754 134423 576779
rect 134582 576778 134616 576783
rect 135035 576779 135093 576826
rect 134571 576767 134616 576778
rect 134582 576754 134616 576767
rect 135047 576754 135081 576779
rect 135240 576778 135274 576783
rect 135693 576779 135751 576826
rect 135229 576767 135274 576778
rect 135240 576754 135274 576767
rect 135705 576754 135739 576779
rect 135898 576778 135932 576783
rect 136351 576779 136409 576826
rect 135887 576767 135932 576778
rect 135898 576754 135932 576767
rect 136363 576754 136397 576779
rect 136468 576754 136490 576820
rect 136496 576778 136546 576820
rect 136556 576778 136590 576783
rect 136496 576767 136590 576778
rect 136496 576754 136546 576767
rect 136556 576754 136590 576767
rect 136670 576754 136704 576928
rect 133478 575279 137578 576754
rect 139346 576749 139380 579068
rect 141434 576749 141468 579068
rect 142864 576749 142898 579068
rect 146196 577424 146230 580282
rect 156922 580244 156956 582118
rect 157710 582008 157714 582118
rect 158590 582116 160240 583554
rect 160694 583552 164318 583556
rect 164861 583552 168485 583567
rect 169688 583554 169714 583846
rect 169716 583554 169770 583846
rect 169830 583818 169854 583920
rect 169858 583886 169882 583892
rect 171054 583886 171088 583954
rect 171156 583886 171334 583924
rect 171348 583886 171872 583924
rect 169858 583852 170538 583886
rect 170628 583852 171334 583886
rect 171386 583852 171872 583886
rect 169858 583846 169882 583852
rect 170566 583686 170600 583802
rect 171054 583686 171088 583852
rect 171156 583814 171214 583852
rect 171814 583814 171872 583852
rect 171168 583686 171213 583814
rect 171313 583802 171369 583813
rect 171324 583686 171369 583802
rect 171826 583686 171871 583814
rect 171940 583686 171974 583954
rect 172244 583686 172278 583954
rect 172346 583852 172850 583924
rect 172954 583892 172988 583954
rect 172346 583814 172404 583852
rect 172358 583686 172403 583814
rect 172829 583802 172885 583813
rect 172840 583686 172885 583802
rect 172954 583702 173006 583892
rect 173016 583720 173022 583926
rect 172954 583686 172988 583702
rect 173016 583686 173050 583720
rect 173130 583686 173164 584114
rect 169968 583652 173424 583686
rect 169968 583554 170002 583652
rect 170566 583622 170600 583652
rect 170698 583622 170718 583652
rect 171054 583622 171088 583652
rect 171168 583622 171213 583652
rect 171324 583622 171369 583652
rect 171826 583622 171871 583652
rect 171940 583622 171974 583652
rect 172244 583622 172278 583652
rect 172358 583622 172403 583652
rect 172840 583622 172885 583652
rect 172954 583622 172988 583652
rect 173016 583622 173022 583652
rect 170106 583584 170750 583622
rect 170764 583584 171408 583622
rect 171422 583584 172066 583622
rect 172080 583584 172724 583622
rect 172738 583584 173062 583622
rect 170144 583554 170750 583584
rect 160694 582614 168485 583552
rect 157744 582008 157748 582086
rect 160694 582084 164318 582614
rect 164861 582084 168485 582614
rect 168738 583550 170750 583554
rect 170802 583556 171408 583584
rect 171460 583556 172066 583584
rect 172082 583556 172724 583584
rect 172776 583556 173062 583584
rect 173130 583556 173164 583652
rect 173554 583556 173574 583740
rect 177970 583717 178004 585030
rect 178628 583717 178662 585030
rect 190092 584962 190126 588654
rect 190092 584874 190150 584962
rect 174440 583556 174474 583574
rect 170802 583550 174474 583556
rect 168738 582116 170388 583550
rect 170554 583512 170612 583550
rect 170566 583464 170611 583512
rect 158618 582050 168485 582084
rect 158618 580244 158652 582050
rect 159060 581976 159086 582034
rect 159088 581976 159114 582006
rect 159196 581970 159230 582050
rect 159954 581970 159988 582050
rect 160694 581970 164318 582050
rect 164502 581970 164536 582050
rect 164861 581970 168485 582050
rect 158682 581908 158754 581946
rect 158804 581936 168485 581970
rect 158720 581340 158754 581908
rect 159060 581870 159086 581930
rect 159088 581898 159114 581930
rect 159183 581924 159184 581925
rect 159184 581923 159185 581924
rect 159184 581324 159185 581325
rect 159183 581323 159184 581324
rect 159196 581312 159230 581936
rect 159242 581924 159243 581925
rect 159941 581924 159942 581925
rect 159241 581923 159242 581924
rect 159942 581923 159943 581924
rect 159241 581324 159242 581325
rect 159942 581324 159943 581325
rect 159242 581323 159243 581324
rect 159941 581323 159942 581324
rect 159954 581312 159988 581936
rect 160000 581924 160001 581925
rect 159999 581923 160000 581924
rect 160694 581844 164318 581936
rect 164489 581924 164490 581925
rect 164490 581923 164491 581924
rect 159999 581324 160000 581325
rect 160000 581323 160001 581324
rect 160694 581312 164426 581844
rect 164490 581324 164491 581325
rect 164489 581323 164490 581324
rect 164502 581312 164536 581936
rect 164548 581924 164549 581925
rect 164547 581923 164548 581924
rect 164861 581850 168485 581936
rect 164547 581324 164548 581325
rect 164548 581323 164549 581324
rect 164696 581312 168485 581850
rect 158682 581250 158754 581288
rect 158804 581278 168485 581312
rect 159183 581266 159184 581267
rect 159184 581265 159185 581266
rect 158720 580682 158754 581250
rect 159066 580660 159086 580724
rect 159094 580660 159114 580696
rect 159184 580666 159185 580667
rect 159183 580665 159184 580666
rect 159196 580654 159230 581278
rect 159242 581266 159243 581267
rect 159941 581266 159942 581267
rect 159241 581265 159242 581266
rect 159942 581265 159943 581266
rect 159241 580666 159242 580667
rect 159942 580666 159943 580667
rect 159242 580665 159243 580666
rect 159941 580665 159942 580666
rect 159954 580654 159988 581278
rect 160000 581266 160001 581267
rect 159999 581265 160000 581266
rect 159999 580666 160000 580667
rect 160000 580665 160001 580666
rect 160694 580654 164426 581278
rect 164489 581266 164490 581267
rect 164490 581265 164491 581266
rect 164452 580660 164460 580738
rect 164490 580666 164491 580667
rect 164489 580665 164490 580666
rect 164502 580654 164536 581278
rect 164548 581266 164549 581267
rect 164547 581265 164548 581266
rect 164547 580666 164548 580667
rect 164548 580665 164549 580666
rect 164696 580654 168485 581278
rect 158682 580592 158754 580630
rect 158804 580620 168485 580654
rect 158720 580246 158754 580592
rect 159066 580560 159086 580614
rect 159094 580588 159114 580614
rect 159183 580608 159184 580609
rect 159184 580607 159185 580608
rect 158682 580244 158754 580246
rect 159196 580244 159230 580620
rect 159242 580608 159243 580609
rect 159941 580608 159942 580609
rect 159241 580607 159242 580608
rect 159942 580607 159943 580608
rect 159954 580244 159988 580620
rect 160000 580608 160001 580609
rect 159999 580607 160000 580608
rect 160694 580406 164426 580620
rect 164452 580528 164460 580614
rect 164489 580608 164490 580609
rect 164490 580607 164491 580608
rect 160694 580244 164318 580406
rect 164502 580244 164536 580620
rect 164548 580608 164549 580609
rect 164547 580607 164548 580608
rect 164696 580412 168485 580620
rect 164861 580244 168485 580412
rect 169688 580346 169714 582116
rect 169716 580346 169770 582116
rect 169808 580244 169842 582116
rect 169890 580244 169900 580346
rect 169968 580244 170002 582116
rect 170082 580244 170127 582116
rect 170566 580244 170600 583464
rect 170642 582992 170662 583544
rect 170640 581982 170662 582992
rect 170698 582936 170718 583544
rect 170729 583500 170785 583511
rect 170696 581982 170718 582936
rect 170740 583464 170785 583500
rect 170740 582696 170774 583464
rect 170842 582888 174474 583550
rect 174866 583240 174876 583598
rect 175009 583579 175678 583717
rect 175696 583585 175724 583598
rect 175752 583585 175780 583598
rect 175846 583579 179109 583717
rect 179252 583644 179276 584750
rect 179286 583610 179310 584784
rect 175009 583545 179109 583579
rect 175009 583497 175678 583545
rect 174866 583026 174894 583240
rect 174866 583020 174876 583026
rect 170842 582818 174466 582888
rect 170740 581848 170785 582696
rect 170740 581836 170788 581848
rect 170642 580244 170662 581782
rect 170698 580244 170718 581782
rect 170740 581188 170785 581836
rect 170792 581798 170800 581836
rect 170842 581668 173556 582818
rect 173618 582636 173622 582818
rect 174396 582636 174430 582818
rect 175009 582810 175680 583497
rect 175045 582636 175079 582810
rect 175159 582636 175193 582670
rect 175521 582636 175555 582810
rect 175635 582636 175680 582810
rect 175696 582636 175724 583539
rect 175752 582886 175780 583539
rect 175846 583497 179109 583545
rect 175806 583486 179109 583497
rect 175817 582806 179109 583486
rect 179280 583016 179282 583598
rect 175817 582636 175862 582806
rect 170806 581542 173556 581668
rect 170806 581412 170812 581542
rect 170740 580244 170774 581188
rect 170842 580434 173556 581542
rect 173608 582602 175862 582636
rect 173608 582502 173642 582602
rect 173737 582534 174328 582581
rect 173660 582502 173664 582509
rect 173608 582446 173664 582502
rect 173784 582500 174328 582534
rect 174270 582453 174328 582500
rect 174396 582475 174430 582602
rect 173608 581304 173642 582446
rect 173658 582122 173664 582446
rect 173686 582150 173692 582446
rect 173711 582441 173767 582452
rect 173660 581397 173664 582122
rect 173722 581465 173767 582441
rect 173862 581916 174054 581968
rect 174282 581916 174327 582453
rect 173838 581848 174327 581916
rect 174282 581453 174327 581848
rect 174374 581668 174378 582453
rect 174348 581458 174378 581668
rect 174396 581499 174448 582475
rect 174380 581465 174448 581499
rect 174374 581453 174378 581458
rect 173737 581406 174328 581453
rect 173784 581372 174328 581406
rect 174270 581356 174328 581372
rect 174313 581341 174328 581356
rect 174396 581304 174430 581465
rect 175045 581304 175079 582602
rect 175521 582581 175555 582602
rect 175635 582581 175680 582602
rect 175147 582568 175682 582581
rect 175696 582568 175724 582602
rect 175100 582500 175117 582534
rect 175147 582500 175724 582568
rect 175147 582453 175205 582500
rect 175159 581453 175204 582453
rect 175521 581453 175555 582500
rect 175623 582453 175681 582500
rect 175696 582453 175724 582500
rect 175810 582574 175862 582602
rect 175635 581453 175680 582453
rect 175696 582452 175736 582453
rect 175685 582441 175741 582452
rect 175696 581465 175741 582441
rect 175752 581662 175764 582481
rect 175696 581453 175736 581458
rect 175147 581440 175682 581453
rect 175696 581440 175724 581453
rect 175100 581372 175117 581406
rect 175147 581372 175724 581440
rect 175752 581425 175764 581458
rect 175810 581377 175878 582574
rect 175147 581356 175205 581372
rect 175147 581341 175162 581356
rect 175159 581304 175193 581338
rect 175521 581304 175555 581372
rect 175623 581356 175681 581372
rect 175635 581304 175680 581356
rect 175696 581304 175724 581372
rect 175806 581366 175878 581377
rect 176293 582032 176327 582806
rect 175810 581304 175862 581366
rect 173608 581270 175862 581304
rect 173618 580434 173622 581270
rect 174396 580434 174430 581270
rect 175045 580724 175079 581270
rect 175159 580724 175193 581270
rect 170842 580400 174850 580434
rect 170842 580379 173556 580400
rect 173618 580379 173622 580400
rect 170842 580332 174328 580379
rect 170842 580298 174159 580332
rect 174202 580298 174328 580332
rect 170842 580292 173556 580298
rect 173612 580292 173670 580298
rect 174270 580292 174328 580298
rect 170842 580244 173566 580292
rect 146298 580210 173566 580244
rect 146310 580180 146344 580210
rect 147068 580180 147102 580210
rect 147826 580180 147860 580210
rect 148584 580180 148618 580210
rect 149342 580180 149376 580210
rect 150100 580180 150134 580210
rect 150858 580180 150892 580210
rect 151616 580180 151650 580210
rect 152030 580188 152950 580210
rect 152030 580180 152064 580188
rect 152916 580180 152950 580188
rect 153132 580180 153166 580210
rect 153220 580188 154140 580210
rect 153220 580180 153254 580188
rect 154106 580180 154140 580188
rect 154530 580196 155450 580210
rect 154530 580180 154564 580196
rect 154648 580180 154682 580196
rect 155406 580180 155450 580196
rect 155698 580204 156618 580210
rect 146310 580158 152384 580180
rect 152398 580158 153900 580180
rect 153914 580158 155564 580180
rect 146310 580142 155564 580158
rect 155698 580142 155732 580204
rect 156158 580180 156204 580204
rect 156136 580152 156204 580180
rect 156210 580152 156226 580174
rect 156136 580148 156226 580152
rect 156130 580142 156232 580148
rect 156584 580142 156618 580204
rect 156858 580208 160410 580210
rect 156858 580142 156892 580208
rect 156922 580180 156956 580208
rect 157710 580180 157714 580208
rect 156894 580142 156956 580180
rect 157652 580176 157690 580180
rect 157704 580176 157714 580180
rect 157744 580180 157748 580208
rect 158618 580180 158652 580208
rect 157744 580178 158448 580180
rect 158462 580178 158656 580180
rect 157652 580156 157714 580176
rect 157726 580156 157742 580178
rect 157652 580142 157742 580156
rect 157744 580142 158656 580178
rect 158720 580142 158754 580208
rect 159196 580180 159230 580208
rect 159954 580180 159988 580208
rect 159168 580178 159230 580180
rect 159926 580178 159988 580180
rect 159168 580156 159234 580178
rect 159242 580156 159258 580178
rect 159168 580142 159258 580156
rect 159926 580156 159992 580178
rect 160000 580156 160016 580178
rect 159926 580142 160016 580156
rect 160376 580142 160410 580208
rect 160694 580180 164318 580210
rect 164502 580180 164536 580210
rect 160684 580142 164318 580180
rect 164474 580142 164536 580180
rect 164678 580208 170558 580210
rect 164678 580196 168485 580208
rect 164678 580142 164712 580196
rect 164861 580142 168485 580196
rect 169090 580180 169552 580192
rect 169808 580180 169842 580208
rect 169890 580180 169900 580208
rect 169968 580180 170002 580208
rect 170082 580180 170127 580208
rect 169022 580178 169060 580180
rect 169074 580178 169084 580180
rect 169022 580174 169088 580178
rect 169090 580174 170306 580180
rect 169022 580142 170306 580174
rect 170524 580142 170558 580208
rect 146310 579266 146344 580142
rect 146372 580108 147108 580142
rect 147034 580102 147052 580108
rect 147062 580074 147108 580108
rect 147118 580108 147860 580142
rect 147888 580108 148624 580142
rect 147118 580102 147136 580108
rect 146304 579242 146350 579266
rect 147068 579242 147102 580074
rect 147826 579266 147860 580108
rect 148550 580102 148568 580108
rect 148578 580074 148624 580108
rect 148634 580108 149376 580142
rect 149404 580108 150140 580142
rect 148634 580102 148652 580108
rect 147820 579242 147866 579266
rect 148584 579242 148618 580074
rect 149342 579266 149376 580108
rect 150066 580102 150084 580108
rect 150094 580074 150140 580108
rect 150150 580108 150892 580142
rect 150920 580108 151656 580142
rect 150150 580102 150168 580108
rect 149336 579242 149382 579266
rect 150100 579242 150134 580074
rect 150858 579266 150892 580108
rect 151582 580102 151600 580108
rect 151610 580074 151656 580108
rect 151666 580108 153172 580142
rect 151666 580102 151684 580108
rect 150852 579242 150898 579266
rect 151616 579242 151650 580074
rect 146304 579204 148474 579242
rect 148556 579204 148618 579242
rect 149314 579210 149382 579242
rect 149308 579204 149382 579210
rect 149392 579204 149410 579210
rect 150072 579204 150134 579242
rect 150830 579210 150898 579242
rect 150824 579204 150898 579210
rect 150908 579204 150926 579210
rect 151588 579204 151650 579242
rect 151736 579210 151752 579264
rect 152030 579204 152064 580108
rect 152206 580086 152812 580108
rect 152133 580036 152189 580047
rect 152144 579324 152189 580036
rect 152144 579242 152178 579324
rect 152144 579204 152182 579242
rect 152190 579210 152240 580080
rect 152246 579210 152268 580080
rect 152362 580048 152420 580086
rect 152374 579324 152419 580048
rect 152791 580036 152847 580047
rect 152802 579324 152847 580036
rect 152374 579242 152408 579324
rect 152346 579204 152408 579242
rect 152802 579242 152836 579324
rect 152802 579204 152840 579242
rect 152916 579204 152950 580108
rect 153098 580102 153116 580108
rect 153126 580074 153172 580108
rect 153182 580128 155450 580142
rect 153182 580108 154688 580128
rect 153182 580102 153200 580108
rect 153076 579210 153078 579912
rect 153132 579242 153166 580074
rect 153104 579204 153166 579242
rect 153220 579204 153254 580108
rect 153396 580086 154002 580108
rect 153878 580048 153936 580086
rect 153323 580036 153379 580047
rect 153334 579324 153379 580036
rect 153334 579242 153368 579324
rect 153890 579266 153935 580048
rect 153958 579450 153976 580076
rect 153986 580047 154032 580048
rect 154034 580047 154060 580076
rect 153981 580036 154060 580047
rect 153986 579394 154060 580036
rect 153992 579382 154060 579394
rect 153884 579242 153935 579266
rect 153956 579242 153986 579382
rect 153992 579242 154037 579382
rect 154106 579242 154140 580108
rect 153334 579204 153372 579242
rect 153556 579204 154470 579242
rect 154530 579204 154564 580108
rect 154614 580102 154632 580108
rect 154642 580074 154688 580108
rect 154648 580060 154688 580074
rect 154690 580108 155450 580128
rect 155468 580108 156956 580142
rect 156968 580108 164536 580142
rect 164548 580108 170558 580142
rect 154690 580102 155398 580108
rect 154690 580094 155312 580102
rect 154690 580088 154716 580094
rect 154648 580056 154682 580060
rect 154690 580056 154694 580088
rect 154633 580044 154636 580055
rect 154648 580052 154688 580056
rect 154690 580052 154693 580056
rect 155338 580055 155342 580056
rect 154648 580044 154700 580052
rect 155291 580044 155347 580055
rect 154644 579954 154700 580044
rect 154644 579242 154728 579954
rect 154620 579210 154728 579242
rect 154738 579210 154756 579982
rect 155302 579324 155347 580044
rect 155366 579466 155398 580102
rect 155302 579242 155336 579324
rect 155406 579266 155450 580108
rect 155400 579242 155450 579266
rect 154620 579204 154682 579210
rect 146304 579182 146350 579204
rect 146360 579182 147102 579204
rect 146310 579102 146344 579182
rect 146372 579170 147102 579182
rect 147130 579182 147866 579204
rect 147876 579182 148618 579204
rect 147130 579170 147860 579182
rect 147888 579170 148618 579182
rect 148630 579182 149382 579204
rect 148630 579170 149376 579182
rect 149388 579170 150134 579204
rect 150146 579182 150898 579204
rect 150146 579170 150892 579182
rect 150904 579170 151650 579204
rect 151662 579170 152408 579204
rect 152420 579170 153166 579204
rect 153178 579170 153935 579204
rect 153940 579182 154682 579204
rect 153952 579170 154682 579182
rect 147068 579102 147102 579170
rect 147826 579102 147860 579170
rect 148584 579102 148618 579170
rect 149342 579102 149376 579170
rect 150020 579102 150028 579164
rect 150048 579102 150084 579164
rect 150100 579102 150134 579170
rect 150858 579102 150892 579170
rect 151616 579102 151650 579170
rect 152030 579102 152064 579170
rect 152144 579102 152178 579170
rect 152374 579102 152408 579170
rect 152802 579102 152836 579170
rect 152916 579102 152950 579170
rect 153132 579102 153166 579170
rect 153220 579102 153254 579170
rect 153334 579102 153368 579170
rect 153890 579102 153935 579170
rect 153992 579102 154037 579170
rect 154106 579102 154140 579170
rect 154530 579102 154564 579170
rect 154644 579102 154682 579170
rect 154690 579102 154693 579210
rect 155302 579204 155340 579242
rect 155378 579210 155450 579242
rect 155372 579204 155450 579210
rect 155456 579204 155474 579210
rect 155698 579204 155732 580108
rect 155874 580102 156480 580108
rect 156152 580064 156210 580102
rect 155801 580052 155846 580063
rect 155812 579242 155846 580052
rect 156164 579242 156198 580064
rect 156459 580052 156504 580063
rect 155812 579204 155850 579242
rect 156136 579204 156198 579242
rect 156470 579242 156504 580052
rect 156470 579204 156508 579242
rect 156584 579204 156618 580108
rect 156858 579210 156892 580108
rect 156922 579454 156956 580108
rect 157034 580106 157640 580108
rect 157676 580106 158298 580108
rect 158322 580106 158956 580108
rect 159008 580106 159614 580108
rect 159666 580106 160272 580108
rect 156994 580100 156996 580102
rect 157022 580100 157024 580102
rect 156966 580068 156996 580100
rect 156966 580062 157012 580068
rect 156966 580056 157038 580062
rect 156972 579656 157038 580056
rect 156972 579454 157012 579656
rect 157056 579628 157066 580090
rect 157646 580067 157664 580072
rect 157619 580056 157664 580067
rect 156922 579266 156962 579454
rect 156916 579242 156962 579266
rect 156894 579238 156962 579242
rect 156966 579238 157012 579454
rect 156894 579210 157012 579238
rect 157630 579242 157664 580056
rect 157676 580068 157726 580106
rect 157630 579238 157668 579242
rect 157676 579238 157714 580068
rect 156858 579204 157006 579210
rect 157630 579204 157714 579238
rect 157744 579242 157748 580106
rect 158322 580102 158384 580106
rect 158310 580072 158322 580102
rect 158338 580100 158384 580102
rect 158322 580067 158328 580068
rect 158277 580056 158333 580067
rect 158288 580044 158333 580056
rect 158382 580044 158408 580100
rect 158426 580068 158484 580106
rect 158288 579716 158352 580044
rect 158288 579242 158333 579716
rect 158382 579242 158384 579716
rect 158438 579242 158483 580068
rect 158618 579242 158652 580106
rect 158720 580024 158754 580106
rect 159184 580068 159242 580106
rect 159942 580068 160000 580106
rect 158935 580056 158980 580067
rect 158946 579996 158980 580056
rect 159196 579996 159230 580068
rect 159593 580056 159638 580067
rect 159604 579996 159638 580056
rect 159954 579996 159988 580068
rect 160251 580056 160296 580067
rect 160262 579996 160296 580056
rect 160376 579996 160410 580108
rect 160694 579996 164318 580108
rect 164452 580002 164460 580080
rect 164490 580008 164491 580009
rect 164489 580007 164490 580008
rect 164502 579996 164536 580108
rect 164547 580008 164548 580009
rect 164548 580007 164549 580008
rect 164678 579996 164712 580108
rect 164854 580094 168485 580108
rect 168498 580106 169762 580108
rect 169798 580106 170420 580108
rect 164781 580044 164826 580055
rect 164792 579996 164826 580044
rect 164861 579996 168485 580094
rect 169038 580068 169084 580106
rect 158682 579934 158754 579972
rect 158804 579962 168485 579996
rect 158720 579366 158754 579934
rect 158946 579338 158980 579962
rect 159196 579338 159230 579962
rect 159604 579338 159638 579962
rect 159954 579338 159988 579962
rect 160262 579338 160296 579962
rect 160376 579338 160410 579962
rect 160638 579956 164318 579962
rect 160694 579954 164318 579956
rect 160666 579928 164318 579954
rect 160694 579338 164318 579928
rect 164452 579864 164460 579956
rect 164489 579950 164490 579951
rect 164490 579949 164491 579950
rect 164490 579350 164491 579351
rect 164489 579349 164490 579350
rect 164502 579338 164536 579962
rect 164548 579950 164549 579951
rect 164547 579949 164548 579950
rect 164547 579350 164548 579351
rect 164548 579349 164549 579350
rect 164678 579338 164712 579962
rect 164792 579338 164826 579962
rect 164861 579338 168485 579962
rect 158682 579276 158754 579314
rect 158804 579304 168485 579338
rect 157744 579204 158656 579242
rect 158720 579204 158754 579276
rect 158946 579242 158980 579304
rect 159196 579242 159230 579304
rect 158946 579204 158984 579242
rect 159168 579204 159230 579242
rect 159604 579242 159638 579304
rect 159954 579242 159988 579304
rect 159604 579204 159642 579242
rect 159926 579204 159988 579242
rect 160262 579242 160296 579304
rect 160262 579204 160300 579242
rect 160376 579204 160410 579304
rect 160694 579242 164318 579304
rect 164489 579292 164490 579293
rect 164490 579291 164491 579292
rect 164502 579242 164536 579304
rect 164548 579292 164549 579293
rect 164547 579291 164548 579292
rect 160684 579204 164318 579242
rect 164474 579204 164536 579242
rect 164678 579204 164712 579304
rect 164792 579242 164826 579304
rect 164792 579204 164830 579242
rect 164861 579204 168485 579304
rect 169050 579242 169084 580068
rect 169090 579554 169552 580106
rect 169798 580068 169854 580106
rect 169741 580056 169796 580067
rect 169752 579772 169796 580056
rect 169688 579736 169714 579772
rect 169716 579764 169796 579772
rect 169690 579630 169714 579736
rect 169746 579630 169796 579764
rect 169022 579238 169084 579242
rect 169094 579238 169128 579554
rect 169022 579204 169128 579238
rect 169148 579470 169498 579504
rect 169148 579204 169182 579470
rect 169268 579402 169378 579440
rect 169306 579368 169378 579402
rect 169251 579318 169307 579329
rect 169339 579318 169395 579329
rect 169262 579242 169307 579318
rect 169350 579242 169395 579318
rect 169464 579242 169498 579470
rect 169752 579430 169796 579630
rect 169690 579326 169714 579430
rect 169746 579326 169796 579430
rect 169752 579242 169796 579326
rect 169226 579238 169796 579242
rect 169798 579242 169853 580068
rect 169968 579242 170002 580106
rect 170082 579242 170127 580106
rect 170399 580056 170444 580067
rect 170410 579242 170444 580056
rect 169798 579238 170306 579242
rect 169226 579204 170306 579238
rect 170410 579204 170448 579242
rect 170524 579204 170558 580108
rect 154694 579170 155450 579204
rect 155452 579170 156198 579204
rect 156210 579182 156962 579204
rect 156966 579182 157714 579204
rect 156210 579170 156956 579182
rect 156968 579170 157714 579182
rect 157726 579170 158483 579204
rect 158500 579170 159230 579204
rect 159242 579170 159988 579204
rect 160000 579170 164536 579204
rect 164548 579170 169084 579204
rect 155302 579102 155336 579170
rect 155406 579102 155450 579170
rect 155698 579102 155732 579170
rect 155812 579102 155846 579170
rect 156164 579102 156198 579170
rect 156470 579102 156504 579170
rect 156584 579102 156618 579170
rect 156858 579102 156892 579170
rect 156922 579102 156956 579170
rect 156972 579102 157006 579170
rect 157630 579102 157664 579170
rect 157676 579102 157714 579170
rect 157744 579102 157748 579170
rect 158288 579102 158333 579170
rect 158438 579102 158483 579170
rect 158618 579102 158652 579170
rect 158720 579106 158754 579170
rect 158682 579102 158792 579106
rect 158946 579102 158980 579170
rect 159196 579102 159230 579170
rect 159604 579102 159638 579170
rect 159954 579102 159988 579170
rect 160262 579102 160296 579170
rect 160376 579102 160410 579170
rect 160694 579118 164318 579170
rect 160712 579102 160746 579118
rect 161470 579102 161504 579118
rect 162178 579102 162212 579118
rect 162228 579102 162262 579118
rect 162292 579102 162326 579118
rect 162950 579102 162984 579118
rect 162986 579102 163020 579118
rect 163064 579102 163098 579118
rect 163368 579102 163402 579118
rect 163482 579102 163516 579118
rect 163744 579102 163778 579118
rect 164140 579102 164174 579118
rect 164254 579102 164288 579118
rect 164502 579102 164536 579170
rect 164678 579102 164712 579170
rect 164792 579102 164826 579170
rect 164861 579102 168485 579170
rect 169050 579102 169084 579170
rect 169094 579170 169853 579204
rect 169870 579170 170558 579204
rect 169094 579102 169128 579170
rect 169148 579102 169182 579170
rect 169262 579142 169307 579170
rect 169350 579142 169395 579170
rect 169272 579106 169374 579126
rect 169268 579102 169378 579106
rect 169464 579102 169498 579170
rect 169752 579102 169796 579170
rect 169798 579102 169853 579170
rect 169968 579102 170002 579170
rect 170082 579102 170127 579170
rect 170410 579102 170444 579170
rect 170524 579102 170558 579170
rect 170566 579102 170600 580210
rect 170642 580148 170662 580210
rect 170698 580148 170718 580210
rect 170740 580180 170774 580210
rect 170740 580142 170778 580180
rect 170842 580142 173566 580210
rect 170612 580108 173566 580142
rect 170642 579210 170662 580102
rect 170698 579210 170718 580102
rect 170740 579242 170774 580108
rect 170842 579751 173566 580108
rect 173574 580251 173670 580292
rect 173574 579751 173622 580251
rect 173624 579751 173669 580251
rect 174129 580239 174185 580250
rect 174140 579763 174185 580239
rect 174202 579751 174216 580292
rect 174230 580251 174328 580292
rect 174230 579751 174272 580251
rect 174282 579751 174327 580251
rect 174396 580070 174430 580400
rect 174346 580042 174522 580070
rect 174346 580024 174466 580042
rect 174346 580008 174522 580024
rect 170842 579704 174328 579751
rect 170842 579670 174159 579704
rect 174202 579670 174328 579704
rect 170842 579602 173556 579670
rect 173612 579654 173670 579670
rect 174270 579654 174328 579670
rect 173618 579602 173622 579654
rect 174313 579639 174328 579654
rect 174396 579602 174430 580008
rect 174466 580006 174522 580008
rect 170842 579568 174850 579602
rect 170740 579204 170778 579242
rect 170842 579204 173556 579568
rect 173618 579550 173622 579568
rect 173596 579342 173622 579550
rect 173618 579337 173622 579342
rect 174396 579250 174430 579568
rect 175009 579532 175236 580724
rect 170612 579170 173556 579204
rect 170642 579102 170662 579164
rect 170698 579102 170718 579164
rect 170740 579102 170774 579170
rect 170842 579118 173556 579170
rect 171324 579102 171358 579118
rect 171398 579102 171438 579118
rect 171458 579102 171494 579118
rect 172056 579102 172127 579118
rect 172714 579102 172759 579118
rect 172840 579102 172885 579118
rect 172954 579102 172988 579118
rect 146292 579068 172988 579102
rect 147068 577424 147102 579068
rect 147826 577424 147860 579068
rect 150020 578536 150028 579068
rect 150048 578564 150084 579068
rect 152030 578908 152064 579068
rect 152144 579060 152189 579068
rect 152374 579048 152419 579068
rect 152802 579060 152847 579068
rect 152168 579010 152812 579048
rect 152206 578976 152812 579010
rect 152362 578960 152420 578976
rect 152374 578908 152408 578960
rect 152916 578908 152950 579068
rect 152030 578874 152950 578908
rect 145192 577406 148760 577424
rect 145192 577404 145736 577406
rect 146074 577396 148760 577406
rect 146196 577368 146230 577396
rect 147068 577368 147102 577396
rect 147826 577368 147860 577396
rect 145192 577350 148760 577368
rect 145192 577348 145792 577350
rect 146018 577340 148760 577350
rect 139310 576713 142934 576749
rect 143626 576718 144999 576749
rect 146196 576718 146230 577340
rect 146310 576718 146344 576778
rect 147068 576740 147102 577340
rect 147826 576740 147860 577340
rect 152374 576749 152408 578874
rect 153132 576749 153166 579068
rect 153220 578908 153254 579068
rect 153334 579060 153379 579068
rect 153890 579048 153935 579068
rect 153992 579060 154037 579068
rect 153358 579010 154002 579048
rect 153396 578976 154002 579010
rect 153878 578960 153936 578976
rect 153890 578908 153924 578960
rect 154106 578908 154140 579068
rect 153220 578874 154140 578908
rect 153484 578436 153824 578472
rect 153852 578436 153866 578674
rect 153446 578398 153786 578434
rect 153890 576749 153924 578874
rect 154530 578316 154564 579068
rect 154644 578468 154682 579068
rect 154648 578456 154682 578468
rect 154690 578456 154693 579068
rect 155302 578468 155347 579068
rect 154648 578418 155312 578456
rect 154648 578316 154682 578418
rect 154690 578368 154694 578418
rect 154706 578384 155312 578418
rect 155416 578316 155450 579068
rect 154530 578282 155450 578316
rect 155698 578324 155732 579068
rect 155812 578476 155857 579068
rect 156164 578464 156209 579068
rect 156470 578476 156515 579068
rect 155836 578426 156480 578464
rect 155874 578392 156480 578426
rect 156152 578376 156210 578392
rect 156164 578324 156198 578376
rect 156584 578324 156618 579068
rect 155698 578290 156618 578324
rect 146348 576718 147860 576740
rect 143626 576713 150034 576718
rect 139310 576684 150034 576713
rect 139310 576679 144999 576684
rect 133478 574308 136770 575279
rect 133254 574274 136770 574308
rect 133266 573478 133300 574274
rect 133478 574206 136770 574274
rect 133312 574172 136770 574206
rect 133478 574064 136770 574172
rect 136782 574064 136804 575279
rect 136862 574970 136890 575279
rect 136918 574064 136963 575279
rect 137032 574064 137066 575279
rect 133478 574030 137440 574064
rect 133478 574000 136770 574030
rect 136782 574000 136804 574030
rect 136918 574000 136963 574030
rect 137032 574000 137066 574030
rect 137394 574000 137428 574030
rect 133478 573962 136774 574000
rect 136782 573962 137428 574000
rect 133478 573928 137428 573962
rect 129215 573224 132832 573242
rect 133116 573224 133352 573478
rect 129215 573184 132868 573224
rect 133112 573188 133352 573224
rect 133478 573188 136770 573928
rect 129215 573076 129249 573184
rect 129215 573048 129260 573076
rect 129691 573048 129725 573184
rect 129734 573052 129780 573184
rect 129808 573108 129836 573184
rect 129808 573052 129852 573108
rect 129734 573048 129796 573052
rect 129198 573014 129268 573048
rect 126972 572980 129268 573014
rect 126972 572783 127056 572980
rect 127538 572959 127572 572980
rect 127538 572912 127585 572959
rect 127600 572918 127614 572980
rect 127628 572918 127670 572980
rect 127680 572959 127714 572980
rect 127794 572959 127828 572980
rect 127680 572912 127727 572959
rect 127750 572912 127828 572959
rect 128196 572928 128242 572959
rect 128184 572912 128242 572928
rect 127182 572878 127828 572912
rect 127840 572878 128242 572912
rect 127109 572819 127154 572830
rect 127120 572783 127154 572819
rect 127538 572795 127572 572878
rect 127680 572783 127714 572878
rect 127794 572853 127828 572878
rect 127794 572830 127846 572853
rect 128184 572831 128242 572878
rect 127767 572819 127846 572830
rect 127778 572783 127846 572819
rect 128196 572795 128230 572831
rect 126972 572742 127068 572783
rect 124240 572736 126954 572742
rect 127006 572736 127068 572742
rect 127120 572736 127167 572783
rect 127510 572736 127557 572783
rect 127668 572736 127726 572783
rect 127766 572736 127846 572783
rect 128168 572736 128215 572783
rect 124240 572702 127557 572736
rect 127600 572702 128215 572736
rect 124240 572634 126954 572702
rect 127006 572686 127068 572702
rect 127006 572634 127062 572686
rect 127084 572634 127090 572696
rect 127120 572652 127154 572702
rect 127668 572686 127726 572702
rect 127766 572686 127846 572702
rect 127680 572652 127714 572686
rect 127120 572634 127165 572652
rect 127680 572634 127725 572652
rect 127772 572634 127776 572686
rect 127794 572668 127846 572686
rect 127778 572634 127846 572668
rect 128310 572634 128344 572980
rect 128409 572878 128424 572912
rect 124240 572600 128344 572634
rect 124240 572369 126954 572600
rect 127006 572582 127062 572600
rect 127084 572582 127090 572600
rect 126994 572374 127056 572582
rect 127058 572374 127090 572528
rect 127006 572369 127062 572374
rect 127114 572369 127118 572528
rect 127120 572369 127165 572600
rect 127680 572369 127725 572600
rect 124240 572322 127725 572369
rect 124240 572288 127062 572322
rect 124240 572220 126954 572288
rect 126988 572282 127062 572288
rect 127072 572288 127725 572322
rect 127072 572282 127090 572288
rect 127006 572226 127062 572282
rect 127006 572220 127056 572226
rect 127058 572220 127062 572226
rect 127120 572220 127165 572288
rect 127236 572226 127725 572288
rect 127680 572220 127725 572226
rect 127772 572220 127776 572600
rect 127794 572220 127846 572600
rect 124240 572186 127846 572220
rect 124138 572028 124178 572058
rect 124240 572046 126954 572186
rect 124204 572030 126954 572046
rect 124198 572028 126954 572030
rect 123668 571848 123990 571870
rect 122530 570984 123622 571006
rect 122530 570980 123582 570984
rect 123058 570786 123084 570980
rect 123114 570786 123140 570980
rect 123150 570626 123184 570980
rect 123150 570620 123246 570626
rect 123366 570620 123400 570980
rect 123480 570620 123525 570980
rect 123808 570786 123842 571848
rect 123808 570620 123853 570786
rect 123922 570620 123956 571848
rect 118259 570608 123956 570620
rect 124138 570608 124172 572028
rect 124204 571920 126954 572028
rect 124204 571790 124210 571920
rect 124240 570812 126954 571920
rect 127006 571682 127040 572186
rect 127058 571775 127062 572186
rect 127120 572120 127165 572186
rect 127680 572120 127725 572186
rect 127120 571843 127154 572120
rect 127680 571831 127714 572120
rect 127716 572046 127748 572120
rect 127772 572046 127776 572186
rect 127716 571836 127776 572046
rect 127794 571877 127846 572186
rect 127778 571843 127846 571877
rect 127716 571831 127748 571836
rect 127772 571831 127776 571836
rect 127668 571784 127748 571831
rect 127182 571750 127726 571784
rect 127668 571734 127748 571750
rect 127682 571719 127748 571734
rect 127682 571682 127714 571719
rect 127716 571682 127748 571719
rect 127794 571682 127828 571843
rect 128443 571682 128477 572980
rect 128557 572943 128591 572980
rect 128545 572928 128591 572943
rect 128545 572912 128603 572928
rect 128919 572912 128953 572980
rect 128962 572959 128996 572980
rect 128962 572912 129009 572959
rect 129033 572912 129067 572980
rect 129076 572912 129122 572980
rect 128482 572878 128515 572912
rect 128545 572878 129122 572912
rect 128545 572831 128603 572878
rect 128557 572652 128591 572831
rect 128919 572720 128953 572878
rect 128962 572720 128996 572878
rect 128557 571831 128602 572652
rect 128776 572630 128996 572720
rect 129033 572652 129067 572878
rect 129076 572831 129122 572878
rect 129076 572775 129134 572831
rect 129094 572738 129134 572775
rect 129150 572738 129162 572859
rect 129198 572779 129268 572980
rect 129674 572784 129796 573048
rect 129808 572784 129824 573052
rect 129094 572732 129128 572738
rect 129198 572732 129570 572779
rect 129674 572738 129780 572784
rect 129808 572738 129852 572784
rect 129674 572732 129744 572738
rect 129094 572698 129744 572732
rect 129094 572692 129128 572698
rect 129094 572652 129134 572692
rect 129033 572630 129078 572652
rect 129094 572630 129139 572652
rect 129150 572630 129162 572692
rect 129198 572630 129664 572698
rect 129674 572692 129744 572698
rect 129756 572692 129780 572738
rect 129784 572732 129852 572738
rect 129873 572732 129907 573184
rect 130349 572779 130383 573184
rect 130337 572732 130383 572779
rect 130392 572775 130442 573184
rect 129784 572698 130383 572732
rect 129784 572692 129836 572698
rect 129674 572636 129780 572692
rect 129674 572630 129744 572636
rect 129752 572630 129780 572636
rect 129808 572630 129836 572692
rect 129873 572652 129907 572698
rect 129873 572630 129918 572652
rect 129928 572630 130310 572698
rect 130337 572682 130383 572698
rect 130349 572652 130383 572682
rect 130349 572630 130394 572652
rect 130414 572630 130442 572775
rect 130470 572630 130498 573184
rect 130506 573032 130565 573184
rect 131007 573032 131041 573184
rect 131048 573032 131082 573184
rect 130506 572720 130580 573032
rect 130506 572630 130786 572720
rect 130986 572712 131082 573032
rect 128776 572596 130786 572630
rect 128776 572288 128988 572596
rect 128642 572272 128988 572288
rect 128642 572226 128953 572272
rect 128919 571831 128953 572226
rect 129033 571831 129078 572596
rect 129094 571843 129139 572596
rect 129150 572040 129162 572596
rect 129198 572592 129664 572596
rect 129674 572592 129744 572596
rect 129208 572272 129664 572592
rect 128498 571750 128515 571784
rect 128545 571750 129078 571831
rect 128545 571734 128603 571750
rect 128545 571719 128591 571734
rect 128557 571682 128591 571719
rect 128919 571682 128953 571750
rect 129033 571682 129078 571750
rect 129094 571831 129134 571836
rect 129094 571682 129122 571831
rect 129150 571803 129162 571836
rect 129208 571682 129260 572272
rect 129452 572264 129664 572272
rect 129480 572184 129648 572264
rect 127006 571648 129260 571682
rect 127016 570812 127020 571648
rect 127682 571200 127714 571648
rect 127716 571234 127748 571648
rect 127794 570812 127828 571648
rect 128443 571102 128477 571648
rect 128557 571102 128591 571648
rect 124240 570778 128248 570812
rect 124240 570710 126954 570778
rect 127016 570726 127020 570778
rect 127022 570726 127069 570757
rect 127010 570710 127069 570726
rect 127510 570710 127557 570757
rect 127680 570726 127726 570757
rect 127668 570710 127726 570726
rect 124240 570676 127557 570710
rect 127600 570676 127726 570710
rect 124240 570670 126954 570676
rect 127010 570670 127068 570676
rect 127668 570670 127726 570676
rect 124240 570608 126964 570670
rect 118076 570574 126964 570608
rect 118076 570374 118110 570574
rect 118259 570544 126964 570574
rect 118214 570506 126964 570544
rect 118252 570472 126964 570506
rect 118156 570458 118258 570462
rect 118184 570433 118230 570434
rect 118179 570430 118235 570433
rect 118179 570422 118246 570430
rect 118190 570386 118246 570422
rect 118190 570374 118224 570386
rect 118228 570385 118246 570386
rect 118259 570385 126964 570472
rect 118228 570380 126964 570385
rect 118236 570374 126964 570380
rect 114092 570340 117720 570374
rect 118042 570340 126964 570374
rect 114092 569716 117716 570340
rect 118076 569716 118110 570340
rect 118190 570328 118224 570340
rect 118228 570328 118246 570334
rect 118190 570242 118246 570328
rect 118190 569729 118235 570242
rect 118259 570088 126964 570340
rect 126972 570629 127068 570670
rect 126972 570129 127020 570629
rect 127022 570129 127056 570629
rect 127527 570617 127572 570628
rect 127538 570141 127572 570617
rect 126972 570088 127069 570129
rect 118259 570082 126954 570088
rect 127010 570082 127069 570088
rect 127510 570082 127557 570129
rect 127600 570088 127614 570670
rect 127628 570629 127726 570670
rect 127628 570129 127670 570629
rect 127680 570129 127714 570629
rect 127794 570448 127828 570778
rect 127744 570386 128040 570448
rect 127628 570088 127726 570129
rect 127668 570082 127726 570088
rect 118259 570048 127557 570082
rect 127600 570048 127726 570082
rect 118259 569980 126954 570048
rect 127010 570032 127068 570048
rect 127668 570032 127726 570048
rect 127016 569980 127020 570032
rect 127711 570017 127726 570032
rect 127794 569980 127828 570386
rect 127864 569980 128380 570002
rect 118259 569946 128380 569980
rect 118190 569728 118236 569729
rect 118190 569716 118224 569728
rect 118228 569722 118230 569728
rect 118236 569727 118237 569728
rect 118259 569727 126954 569946
rect 127016 569928 127020 569946
rect 126994 569902 127020 569928
rect 127022 569727 127056 569946
rect 118236 569716 126954 569727
rect 112080 569658 112190 569692
rect 112202 569682 113842 569716
rect 114092 569682 117720 569716
rect 118042 569714 126954 569716
rect 127668 569715 127726 569766
rect 118042 569682 121883 569714
rect 112331 569670 112332 569671
rect 112344 569670 112378 569682
rect 112390 569670 112391 569671
rect 112989 569670 112990 569671
rect 113002 569670 113036 569682
rect 113048 569670 113049 569671
rect 113647 569670 113648 569671
rect 113660 569670 113694 569682
rect 112332 569669 112333 569670
rect 112344 569669 112390 569670
rect 112990 569669 112991 569670
rect 113002 569669 113048 569670
rect 113648 569669 113649 569670
rect 112080 569654 112212 569658
rect 112118 569644 112212 569654
rect 112118 569258 112190 569644
rect 112344 569258 112389 569669
rect 113002 569258 113047 569669
rect 113660 569258 113705 569670
rect 112118 569086 112152 569258
rect 112332 569070 112333 569071
rect 112331 569069 112332 569070
rect 112344 569058 112378 569258
rect 112389 569070 112390 569071
rect 112990 569070 112991 569071
rect 112390 569069 112391 569070
rect 112989 569069 112990 569070
rect 113002 569058 113036 569258
rect 113047 569070 113048 569071
rect 113648 569070 113649 569071
rect 113048 569069 113049 569070
rect 113647 569069 113648 569070
rect 113660 569058 113694 569258
rect 113774 569058 113808 569682
rect 114092 569496 117716 569682
rect 115576 569286 115610 569496
rect 115690 569438 115735 569496
rect 116348 569438 116393 569496
rect 115714 569388 116358 569426
rect 115752 569354 116358 569388
rect 116462 569286 116496 569496
rect 115576 569252 116496 569286
rect 116766 569286 116800 569496
rect 116880 569438 116925 569496
rect 117538 569438 117583 569496
rect 116904 569388 117548 569426
rect 116942 569354 117548 569388
rect 117652 569286 117686 569496
rect 116766 569252 117686 569286
rect 116938 569142 117488 569144
rect 116966 569114 117460 569116
rect 118076 569058 118110 569682
rect 118190 569670 118224 569682
rect 118228 569670 118230 569676
rect 118236 569670 118237 569671
rect 118190 569669 118236 569670
rect 118190 569258 118235 569669
rect 118190 569058 118224 569258
rect 118228 569064 118230 569142
rect 118235 569070 118236 569071
rect 118236 569069 118237 569070
rect 118259 569058 121883 569682
rect 112202 569024 113808 569058
rect 114976 569024 121883 569058
rect 112344 568944 112378 569024
rect 113002 568944 113036 569024
rect 113660 568944 113694 569024
rect 113774 568944 113808 569024
rect 118076 568944 118110 569024
rect 118190 568944 118224 569024
rect 118228 568944 118230 569018
rect 118259 568944 121883 569024
rect 112016 568910 121883 568944
rect 112918 568526 112936 568910
rect 112974 568526 112992 568858
rect 112158 568438 112706 568472
rect 112158 568156 112192 568438
rect 112344 568358 112378 568438
rect 112520 568358 112531 568369
rect 112222 568314 112294 568352
rect 112260 568280 112294 568314
rect 112344 568324 112531 568358
rect 112331 568312 112332 568313
rect 112332 568311 112333 568312
rect 112332 568282 112333 568283
rect 112331 568281 112332 568282
rect 112344 568270 112378 568324
rect 112532 568314 112604 568352
rect 112390 568312 112391 568313
rect 112389 568311 112390 568312
rect 112389 568282 112390 568283
rect 112390 568281 112391 568282
rect 112520 568270 112531 568281
rect 112570 568280 112604 568314
rect 112344 568236 112531 568270
rect 112344 568156 112378 568236
rect 112672 568156 112706 568438
rect 112158 568122 112706 568156
rect 112756 568064 113394 568526
rect 112918 568050 112936 568064
rect 112974 568050 112992 568064
rect 112158 567962 112706 567996
rect 112158 567680 112192 567962
rect 112344 567882 112378 567962
rect 112520 567882 112531 567893
rect 112222 567842 112294 567876
rect 112344 567848 112531 567882
rect 112222 567838 112302 567842
rect 112260 567804 112302 567838
rect 112331 567836 112332 567837
rect 112332 567835 112333 567836
rect 112332 567806 112333 567807
rect 112331 567805 112332 567806
rect 112276 567788 112302 567804
rect 112332 567786 112338 567800
rect 112344 567794 112378 567848
rect 112532 567838 112604 567876
rect 112390 567836 112391 567837
rect 112389 567835 112390 567836
rect 112389 567806 112390 567807
rect 112390 567805 112391 567806
rect 112384 567794 112438 567800
rect 112520 567794 112531 567805
rect 112570 567804 112604 567838
rect 112344 567760 112531 567794
rect 112344 567680 112378 567760
rect 112672 567680 112706 567962
rect 112158 567646 112706 567680
rect 112756 567588 113394 568050
rect 113654 567860 113656 568874
rect 113774 567168 113808 568910
rect 118076 568756 118110 568910
rect 118228 568834 118230 568910
rect 118259 568874 121883 568910
rect 118259 568624 119032 568874
rect 100940 567136 101020 567150
rect 101416 567136 101502 567150
rect 98922 567072 102378 567106
rect 100046 565902 100080 567072
rect 100704 565902 100738 567072
rect 97300 565858 97560 565892
rect 97300 565812 97334 565858
rect 100818 565812 100852 567072
rect 101236 567036 101698 567072
rect 101712 567036 102174 567072
rect 101712 566456 101952 567036
rect 118295 565789 118329 568624
rect 118409 568530 118443 568624
rect 119033 568530 119038 568704
rect 119067 568530 119101 568874
rect 119208 568632 120200 568874
rect 119725 568530 119759 568632
rect 120368 568530 121883 568874
rect 118409 568489 119038 568530
rect 119039 568517 119101 568530
rect 119039 568489 119107 568517
rect 118409 568483 119107 568489
rect 119117 568483 119135 568489
rect 119198 568483 120210 568530
rect 120355 568489 121883 568530
rect 120349 568483 121883 568489
rect 118409 568482 118443 568483
rect 118471 568482 119107 568483
rect 118409 568415 118449 568482
rect 118459 568449 119107 568482
rect 119113 568449 119759 568483
rect 119787 568449 121883 568483
rect 118459 568443 118477 568449
rect 119033 568443 119051 568449
rect 118409 568381 118443 568415
rect 119033 568381 119038 568443
rect 119061 568415 119107 568449
rect 119117 568443 119135 568449
rect 119067 568381 119101 568415
rect 119725 568381 119759 568449
rect 120349 568443 120367 568449
rect 120368 568381 121883 568449
rect 118391 568347 121883 568381
rect 118409 567258 118443 568347
rect 119033 567116 119038 568347
rect 119067 567116 119072 568347
rect 119725 567258 119759 568347
rect 120368 567954 121883 568347
rect 122492 568582 122526 569714
rect 122546 569368 122580 569714
rect 122649 569696 122705 569707
rect 122737 569696 122793 569707
rect 122660 569520 122705 569696
rect 122748 569520 122793 569696
rect 122666 569470 122776 569508
rect 122704 569436 122776 569470
rect 122862 569368 122896 569714
rect 122546 569334 122896 569368
rect 122542 569156 122560 569258
rect 122492 568326 122532 568582
rect 122540 568354 122560 568554
rect 122492 567954 122526 568326
rect 123060 568132 123084 569156
rect 123116 568916 123140 569156
rect 123150 567954 123184 569714
rect 123366 568404 123400 569714
rect 123480 568544 123525 569714
rect 123808 569258 123853 569714
rect 123808 568544 123842 569258
rect 123480 568506 123704 568544
rect 123808 568506 123846 568544
rect 123922 568506 123956 569714
rect 124138 568544 124172 569714
rect 124240 569566 126954 569714
rect 127338 569690 127726 569712
rect 127338 569678 127690 569690
rect 127338 569618 127372 569678
rect 127476 569634 127590 569648
rect 127794 569628 127828 569946
rect 127864 569910 128380 569946
rect 128407 569910 128634 571102
rect 127338 569616 127349 569618
rect 127361 569616 127372 569618
rect 127338 569566 127372 569616
rect 127514 569596 127552 569610
rect 127694 569566 127728 569616
rect 124240 569532 127732 569566
rect 124240 569496 126954 569532
rect 124796 568544 124830 569496
rect 125454 568544 125488 569496
rect 126112 568544 126146 569496
rect 126770 568544 126804 569496
rect 124110 568540 124172 568544
rect 124768 568540 124830 568544
rect 125426 568540 125488 568544
rect 126084 568540 126146 568544
rect 124110 568512 124178 568540
rect 124768 568512 124836 568540
rect 125426 568512 125494 568540
rect 126084 568512 126152 568540
rect 126742 568512 126804 568544
rect 124104 568506 124178 568512
rect 124188 568506 124206 568512
rect 124762 568506 124836 568512
rect 124846 568506 124864 568512
rect 125420 568506 125494 568512
rect 125504 568506 125522 568512
rect 126078 568506 126152 568512
rect 126162 568506 126180 568512
rect 126736 568506 126804 568512
rect 123480 568404 123525 568506
rect 123542 568472 124178 568506
rect 124184 568472 124836 568506
rect 124842 568472 125494 568506
rect 125500 568472 126152 568506
rect 126158 568472 126804 568506
rect 123808 568408 123842 568472
rect 123808 568404 123853 568408
rect 123922 568404 123956 568472
rect 124104 568466 124122 568472
rect 124132 568438 124178 568472
rect 124188 568466 124206 568472
rect 124762 568466 124780 568472
rect 124790 568438 124836 568472
rect 124846 568466 124864 568472
rect 125420 568466 125438 568472
rect 125448 568438 125494 568472
rect 125504 568466 125522 568472
rect 126078 568466 126096 568472
rect 126106 568438 126152 568472
rect 126162 568466 126180 568472
rect 126736 568466 126754 568472
rect 126764 568438 126804 568472
rect 124138 568404 124172 568438
rect 124796 568404 124830 568438
rect 125454 568404 125488 568438
rect 126112 568404 126146 568438
rect 126770 568404 126804 568438
rect 123366 568370 126838 568404
rect 123366 567954 123400 568370
rect 123480 567954 123525 568370
rect 123808 567954 123853 568370
rect 123922 567954 123956 568370
rect 124138 567954 124172 568370
rect 120368 567880 124428 567954
rect 120368 567560 124512 567880
rect 120368 567060 124428 567560
rect 120368 567036 121883 567060
rect 123366 565812 123400 567060
rect 123480 565902 123514 567060
rect 124138 565902 124172 567060
rect 126884 565812 126918 569496
rect 127338 569242 127372 569532
rect 127440 569507 127498 569529
rect 127568 569507 127626 569529
rect 127694 569242 127728 569532
rect 127472 569194 127592 569214
rect 127778 569196 128018 569496
rect 127778 569194 128068 569196
rect 127466 569166 127620 569186
rect 127778 569168 128018 569194
rect 127778 569166 128096 569168
rect 127778 569110 128018 569166
rect 128407 569110 128494 569910
rect 128443 567348 128477 569110
rect 128557 568517 128591 569910
rect 128557 568415 128597 568517
rect 128607 568483 128625 568489
rect 128919 568483 128953 571648
rect 129033 571308 129078 571648
rect 129094 571308 129122 571648
rect 129215 571308 129260 571648
rect 129691 571308 129736 572592
rect 129752 571308 129780 572596
rect 129808 571308 129836 572596
rect 129873 571308 129918 572596
rect 129928 572272 130310 572596
rect 129928 572264 130140 572272
rect 130349 572120 130394 572596
rect 130349 571308 130383 572120
rect 130414 571308 130442 572596
rect 130470 571308 130498 572596
rect 130510 572576 130786 572596
rect 130531 572272 130786 572576
rect 130794 572632 131082 572712
rect 131084 572632 131112 573184
rect 131140 572793 131223 573184
rect 131140 572632 131168 572793
rect 131189 572734 131223 572793
rect 131665 572781 131699 573184
rect 131653 572734 131711 572781
rect 131736 572740 131764 573184
rect 131792 573010 131881 573184
rect 131792 572790 131902 573010
rect 131792 572781 131820 572790
rect 131832 572781 131902 572790
rect 131792 572734 131902 572781
rect 131961 572734 131995 573184
rect 132323 572781 132357 573184
rect 132311 572734 132369 572781
rect 131189 572700 132369 572734
rect 131189 572652 131223 572700
rect 131189 572632 131234 572652
rect 131270 572632 131652 572700
rect 131653 572684 131711 572700
rect 131665 572652 131699 572684
rect 131665 572632 131710 572652
rect 131792 572632 131820 572694
rect 131832 572632 131902 572700
rect 131916 572632 132128 572700
rect 132311 572684 132369 572700
rect 132240 572644 132254 572650
rect 132280 572644 132282 572678
rect 132323 572669 132369 572684
rect 132437 572743 132471 573184
rect 132478 572777 132505 573184
rect 132437 572700 132466 572743
rect 132240 572638 132280 572644
rect 132323 572632 132357 572669
rect 132437 572644 132471 572700
rect 132514 572650 132518 572694
rect 132408 572638 132518 572644
rect 132437 572632 132471 572638
rect 130794 572598 132530 572632
rect 132672 572622 132680 573184
rect 133112 573154 136770 573188
rect 133112 573086 133352 573154
rect 133362 573086 133409 573133
rect 133112 573052 133409 573086
rect 133112 572758 133352 573052
rect 133379 572993 133424 573004
rect 133390 572817 133424 572993
rect 133362 572758 133409 572805
rect 133112 572732 133409 572758
rect 133478 572732 136770 573154
rect 133112 572698 136770 572732
rect 132808 572670 132928 572672
rect 133112 572656 133352 572698
rect 133478 572656 136770 572698
rect 133112 572652 136770 572656
rect 136782 572652 136804 573928
rect 132780 572642 132956 572644
rect 130794 572576 131056 572598
rect 130531 572120 130576 572272
rect 130794 572264 131006 572576
rect 131007 572120 131052 572576
rect 130531 571308 130565 572120
rect 128962 571274 130565 571308
rect 128962 569976 128996 571274
rect 129033 571268 129078 571274
rect 129094 571268 129122 571274
rect 129033 571253 129122 571268
rect 129215 571253 129260 571274
rect 129691 571268 129736 571274
rect 129752 571268 129780 571274
rect 129691 571253 129780 571268
rect 129808 571253 129836 571274
rect 129873 571253 129918 571274
rect 129033 571234 130166 571253
rect 129033 571124 129067 571234
rect 129070 571212 130166 571234
rect 129076 571206 129736 571212
rect 129749 571206 130166 571212
rect 130349 571206 130383 571274
rect 129076 571166 129122 571206
rect 129126 571172 129736 571206
rect 129126 571166 129150 571172
rect 129070 571124 129122 571166
rect 129033 571122 129122 571124
rect 129033 571113 129140 571122
rect 129033 569998 129067 571113
rect 129076 570882 129140 571113
rect 129076 570137 129122 570882
rect 129150 570854 129168 571150
rect 129215 571092 129260 571172
rect 129691 571166 129736 571172
rect 129756 571166 129780 571206
rect 129784 571172 130383 571206
rect 129784 571166 129836 571172
rect 129691 571092 129780 571166
rect 129070 570084 129122 570137
rect 129098 570038 129122 570084
rect 129126 570078 129150 570084
rect 129215 570078 129249 571092
rect 129691 570078 129725 571092
rect 129734 570398 129780 571092
rect 129808 570454 129836 571166
rect 129873 571092 129918 571172
rect 130349 571124 130383 571172
rect 130414 571129 130442 571274
rect 130392 571124 130442 571129
rect 130349 571122 130442 571124
rect 130470 571178 130498 571274
rect 130506 571178 130565 571274
rect 130470 571122 130565 571178
rect 130349 571113 130464 571122
rect 129808 570398 129852 570454
rect 129734 570137 129796 570398
rect 129728 570130 129796 570137
rect 129808 570130 129824 570398
rect 129728 570084 129780 570130
rect 129808 570084 129852 570130
rect 129126 570044 129725 570078
rect 129126 570038 129150 570044
rect 129070 569998 129122 570038
rect 129033 569982 129122 569998
rect 129033 569976 129078 569982
rect 129094 569976 129122 569982
rect 129215 569998 129249 570044
rect 129252 569998 129664 570044
rect 129215 569976 129664 569998
rect 129691 569998 129725 570044
rect 129756 570038 129780 570084
rect 129784 570078 129852 570084
rect 129873 570078 129907 571092
rect 130349 570078 130383 571113
rect 130392 570774 130464 571113
rect 130470 570774 130492 571122
rect 130506 570774 130565 571122
rect 130392 570121 130442 570774
rect 129784 570044 130383 570078
rect 129784 570038 129836 570044
rect 129728 569998 129780 570038
rect 129691 569982 129780 569998
rect 129691 569976 129736 569982
rect 129752 569976 129780 569982
rect 129808 569976 129836 570038
rect 129873 569998 129907 570044
rect 129873 569976 129918 569998
rect 129928 569976 130310 570044
rect 130349 569998 130383 570044
rect 130349 569976 130394 569998
rect 130414 569976 130442 570121
rect 130470 570718 130565 570774
rect 130470 569976 130498 570718
rect 130506 569998 130565 570718
rect 130782 570058 130786 570066
rect 130506 569976 130576 569998
rect 128962 569942 130576 569976
rect 129033 569466 129078 569942
rect 129033 568530 129067 569466
rect 129021 568483 129080 568530
rect 129094 568489 129122 569942
rect 129215 569618 129664 569942
rect 129215 569466 129260 569618
rect 129452 569610 129664 569618
rect 129691 569466 129736 569942
rect 129215 568530 129249 569466
rect 129691 568530 129725 569466
rect 129215 568483 129262 568530
rect 129679 568483 129738 568530
rect 129752 568489 129780 569942
rect 129808 568489 129836 569942
rect 129873 569466 129918 569942
rect 129928 569618 130310 569942
rect 129928 569610 130140 569618
rect 130349 569466 130394 569942
rect 129873 568530 129907 569466
rect 130349 568530 130383 569466
rect 129873 568483 129920 568530
rect 130337 568483 130396 568530
rect 130414 568489 130442 569942
rect 130470 568489 130498 569942
rect 130531 569466 130576 569942
rect 130794 569618 130798 570058
rect 131007 569998 131041 572120
rect 131084 571310 131112 572598
rect 131140 571310 131168 572598
rect 131189 572120 131234 572598
rect 131270 572264 131652 572598
rect 131665 572120 131710 572598
rect 131189 571310 131223 572120
rect 131665 571310 131699 572120
rect 131792 571310 131820 572598
rect 131832 572554 131902 572598
rect 131847 572120 131892 572554
rect 131916 572488 132214 572598
rect 131916 572264 132128 572488
rect 132252 572450 132254 572458
rect 132280 572422 132282 572458
rect 131847 571310 131881 572120
rect 131961 571310 131995 572264
rect 132323 571310 132357 572598
rect 132437 571310 132471 572598
rect 133112 572596 136781 572652
rect 133112 572586 133352 572596
rect 133152 572572 133186 572586
rect 133478 572572 136781 572596
rect 132658 572562 132662 572572
rect 132832 572392 132908 572394
rect 132804 572364 132936 572366
rect 132814 572142 132924 572162
rect 132852 572104 132886 572124
rect 133134 572120 136781 572572
rect 133134 571952 136770 572120
rect 131048 571276 132530 571310
rect 131048 569998 131082 571276
rect 131084 571122 131112 571276
rect 131140 571126 131168 571276
rect 131189 571208 131223 571276
rect 131665 571208 131699 571276
rect 131792 571255 131820 571276
rect 131792 571208 131839 571255
rect 131189 571174 131839 571208
rect 131847 571208 131881 571276
rect 131961 571208 131995 571276
rect 132323 571239 132357 571276
rect 132323 571224 132369 571239
rect 132311 571208 132369 571224
rect 131847 571174 132369 571208
rect 131189 571126 131223 571174
rect 131140 571122 131223 571126
rect 131151 571115 131223 571122
rect 131162 570866 131223 571115
rect 131007 569978 131082 569998
rect 131084 569978 131112 570866
rect 131140 570139 131223 570866
rect 131140 569978 131168 570139
rect 131189 570080 131223 570139
rect 131665 570080 131699 571174
rect 131736 570086 131764 571168
rect 131792 571126 131820 571168
rect 131847 571126 131881 571174
rect 131792 570139 131881 571126
rect 131792 570127 131820 570139
rect 131792 570080 131839 570127
rect 131189 570046 131839 570080
rect 131847 570080 131881 570139
rect 131961 570080 131995 571174
rect 132311 571127 132369 571174
rect 132437 571208 132471 571276
rect 132437 571165 132466 571208
rect 132323 570127 132357 571127
rect 132311 570080 132369 570127
rect 131847 570046 132369 570080
rect 131189 569998 131223 570046
rect 131189 569978 131234 569998
rect 131270 569978 131652 570046
rect 131665 569998 131699 570046
rect 131665 569978 131710 569998
rect 131792 569978 131820 570040
rect 131847 569998 131881 570046
rect 131847 569978 131892 569998
rect 131916 569978 132128 570046
rect 132311 570030 132369 570046
rect 132323 570015 132369 570030
rect 132437 570089 132471 571165
rect 132478 570123 132505 571131
rect 132650 570952 132662 571208
rect 132678 571006 132718 571238
rect 133152 571006 133186 571952
rect 133266 571870 133372 571952
rect 133266 571006 133300 571870
rect 133478 571006 136770 571952
rect 132678 570980 136770 571006
rect 133152 570824 133186 570980
rect 133266 570824 133300 570980
rect 132618 570534 132626 570588
rect 133116 570570 133352 570824
rect 133112 570534 133352 570570
rect 133478 570534 136770 570980
rect 132437 570046 132466 570089
rect 132240 569990 132254 569996
rect 132240 569984 132317 569990
rect 132323 569978 132357 570015
rect 132437 569990 132471 570046
rect 132514 569996 132518 570040
rect 132363 569984 132518 569990
rect 132437 569978 132471 569984
rect 131007 569944 132530 569978
rect 132672 569968 132680 570534
rect 133112 570500 136770 570534
rect 133112 570432 133352 570500
rect 133362 570432 133409 570479
rect 133112 570398 133409 570432
rect 133112 570151 133352 570398
rect 133379 570339 133424 570350
rect 133390 570163 133424 570339
rect 133112 570125 133409 570151
rect 133112 570104 133352 570125
rect 133112 570078 133362 570104
rect 133478 570078 136770 570500
rect 133112 570044 136770 570078
rect 132808 570016 132928 570018
rect 133112 570002 133352 570044
rect 133402 570016 133404 570036
rect 133402 570002 133410 570008
rect 132780 569988 132956 569990
rect 133112 569976 133442 570002
rect 133478 569998 136770 570044
rect 136782 569998 136804 572120
rect 133478 569976 136781 569998
rect 131007 569466 131052 569944
rect 130531 568530 130565 569466
rect 131007 568530 131041 569466
rect 130531 568483 130578 568530
rect 130995 568483 131054 568530
rect 131084 568489 131112 569944
rect 131140 568489 131168 569944
rect 131189 569466 131234 569944
rect 131270 569892 131652 569944
rect 131665 569892 131710 569944
rect 131270 569610 131718 569892
rect 131189 568530 131223 569466
rect 131644 569238 131718 569610
rect 131665 568530 131699 569238
rect 131189 568483 131236 568530
rect 131653 568483 131712 568530
rect 131792 568489 131820 569944
rect 131847 569466 131892 569944
rect 131916 569834 132214 569944
rect 131916 569610 132128 569834
rect 131847 568530 131881 569466
rect 131847 568483 131894 568530
rect 131961 568483 131995 569610
rect 132323 568530 132357 569944
rect 132295 568489 132357 568530
rect 132289 568483 132357 568489
rect 128603 568449 132357 568483
rect 128607 568443 128625 568449
rect 128557 568381 128591 568415
rect 128919 568381 128953 568449
rect 129021 568433 129079 568449
rect 129033 568381 129067 568433
rect 129094 568381 129122 568443
rect 129215 568381 129249 568449
rect 129679 568433 129737 568449
rect 129691 568381 129725 568433
rect 129752 568381 129780 568443
rect 129808 568381 129836 568443
rect 129873 568381 129907 568449
rect 130337 568433 130395 568449
rect 130349 568381 130383 568433
rect 130414 568381 130442 568443
rect 130470 568381 130498 568443
rect 130531 568381 130565 568449
rect 130995 568433 131053 568449
rect 131007 568381 131041 568433
rect 131084 568381 131112 568443
rect 131140 568381 131168 568443
rect 131189 568381 131223 568449
rect 131653 568433 131711 568449
rect 131665 568381 131699 568433
rect 131792 568381 131820 568443
rect 131847 568381 131881 568449
rect 131961 568381 131995 568449
rect 132289 568443 132307 568449
rect 132317 568415 132357 568449
rect 132323 568381 132357 568415
rect 128539 568347 132369 568381
rect 132375 568347 132391 568381
rect 127472 566540 127592 566560
rect 127778 566542 128018 567094
rect 127778 566540 128068 566542
rect 127466 566512 127620 566532
rect 127778 566514 128018 566540
rect 127778 566512 128096 566514
rect 127778 566456 128018 566512
rect 128407 566456 128494 567348
rect 128443 565789 128477 566456
rect 128919 565829 128953 568347
rect 129033 565888 129067 568347
rect 129094 568002 129122 568347
rect 129094 565835 129122 566814
rect 129215 565888 129249 568347
rect 129691 565888 129725 568347
rect 129752 568002 129780 568347
rect 129808 568002 129836 568347
rect 129752 565835 129780 566814
rect 129808 565835 129836 566814
rect 129873 565888 129907 568347
rect 130349 565888 130383 568347
rect 130414 568002 130442 568347
rect 130470 568002 130498 568347
rect 130414 565835 130442 566814
rect 130470 565835 130498 566814
rect 130531 565888 130565 568347
rect 131007 565888 131041 568347
rect 131084 568002 131112 568347
rect 131140 568002 131168 568347
rect 131084 565835 131112 566814
rect 131140 565835 131168 566814
rect 131189 565888 131223 568347
rect 131665 565888 131699 568347
rect 131792 568002 131820 568347
rect 131792 565835 131820 566814
rect 131847 565888 131881 568347
rect 131961 565829 131995 568347
rect 128919 565795 131995 565829
rect 128919 565779 128953 565795
rect 129094 565782 129122 565789
rect 129752 565782 129780 565789
rect 129808 565782 129836 565789
rect 130414 565782 130442 565789
rect 130470 565782 130498 565789
rect 131084 565782 131112 565789
rect 131140 565782 131168 565789
rect 131792 565782 131820 565789
rect 128919 565768 128930 565779
rect 128942 565768 128953 565779
rect 131961 565779 131995 565795
rect 132437 565789 132471 569944
rect 133112 569942 136781 569976
rect 133112 569932 133352 569942
rect 133478 569918 136781 569942
rect 132658 569908 132662 569918
rect 133134 569906 136781 569918
rect 133514 569786 133548 569906
rect 132832 569738 132908 569740
rect 132804 569710 132936 569712
rect 132774 569582 133046 569702
rect 132724 569488 133046 569582
rect 132852 569450 132886 569470
rect 133486 569430 133548 569786
rect 133514 565812 133548 569430
rect 133628 568540 133662 569906
rect 133694 569706 133700 569808
rect 133722 569734 133728 569808
rect 133628 568438 133668 568540
rect 133678 568506 133696 568512
rect 133990 568506 134024 569906
rect 134088 569590 134096 569906
rect 134104 569466 134149 569906
rect 134180 569534 134208 569734
rect 134286 569466 134331 569906
rect 134348 569590 134750 569906
rect 134538 569586 134750 569590
rect 134762 569466 134807 569906
rect 134104 568544 134138 569466
rect 134092 568506 134150 568544
rect 134180 568512 134208 569334
rect 134286 568544 134320 569466
rect 134762 568544 134796 569466
rect 134286 568506 134324 568544
rect 134750 568506 134808 568544
rect 134832 568512 134860 569906
rect 134888 568512 134916 569906
rect 134944 569466 134989 569906
rect 135136 569590 135398 569906
rect 135402 569590 135410 569900
rect 135136 569586 135226 569590
rect 135420 569466 135465 569906
rect 134944 568544 134978 569466
rect 135420 568544 135454 569466
rect 134944 568506 134982 568544
rect 135408 568506 135466 568544
rect 135490 568512 135518 569906
rect 135546 568512 135574 569906
rect 135602 569466 135647 569906
rect 135662 569590 136066 569906
rect 135854 569584 136066 569590
rect 136078 569466 136123 569906
rect 135602 568544 135636 569466
rect 136078 568544 136112 569466
rect 135602 568506 135640 568544
rect 136066 568506 136124 568544
rect 136154 568512 136182 569906
rect 136210 568512 136238 569906
rect 136260 569466 136305 569906
rect 136330 569584 136710 569906
rect 136498 569572 136710 569584
rect 136718 569572 136722 569892
rect 136736 569466 136781 569906
rect 136260 568544 136294 569466
rect 136736 568544 136770 569466
rect 136782 569430 136804 569466
rect 136260 568506 136298 568544
rect 136724 568506 136782 568544
rect 136862 568512 136890 573782
rect 136918 572908 136963 573928
rect 136894 572674 136986 572908
rect 137032 572674 137066 573928
rect 136894 572450 137186 572674
rect 136918 569430 136963 572450
rect 136974 572226 137186 572450
rect 136918 568544 136952 569430
rect 136918 568506 136956 568544
rect 137032 568506 137066 572226
rect 137394 568544 137428 573928
rect 137508 573182 137542 575279
rect 138591 570002 138625 576617
rect 138755 576584 138758 576604
rect 139310 576584 142934 576679
rect 143414 576649 143612 576679
rect 143626 576649 144999 576679
rect 143318 576646 144999 576649
rect 143318 576618 143352 576646
rect 143284 576611 143386 576618
rect 143576 576617 143596 576646
rect 138727 576550 138730 576576
rect 138755 576571 138822 576584
rect 139270 576571 142934 576584
rect 139310 575302 142934 576571
rect 143318 576148 143352 576611
rect 143456 576577 143471 576611
rect 143487 576578 143512 576611
rect 143514 576578 143545 576611
rect 143494 576568 143509 576578
rect 143523 576568 143532 576578
rect 143561 576577 143570 576611
rect 143626 576584 144999 576646
rect 146196 576616 146230 576684
rect 146310 576654 146344 576684
rect 146348 576654 147860 576684
rect 146298 576616 147922 576654
rect 147936 576616 148474 576654
rect 148542 576650 148580 576654
rect 148542 576616 148582 576650
rect 145812 576584 147922 576616
rect 143596 576571 144999 576584
rect 145008 576576 145076 576584
rect 145142 576576 145218 576584
rect 145666 576576 145734 576584
rect 145800 576582 147922 576584
rect 147974 576582 148582 576616
rect 145800 576576 145882 576582
rect 143478 576544 143548 576568
rect 143499 576530 143533 576534
rect 143465 576496 143466 576501
rect 143487 576497 143545 576530
rect 143576 576528 143596 576571
rect 143421 576485 143466 576496
rect 143432 576309 143466 576485
rect 143465 576293 143466 576309
rect 143499 576297 143533 576497
rect 143560 576496 143567 576501
rect 143549 576485 143594 576496
rect 143560 576309 143594 576485
rect 143487 576284 143546 576297
rect 143560 576293 143567 576309
rect 143487 576216 143566 576284
rect 143487 576200 143545 576216
rect 143499 576148 143533 576182
rect 143626 576148 144999 576571
rect 143318 576114 144999 576148
rect 143626 576064 144999 576114
rect 143300 575444 144999 576064
rect 145666 575574 145802 575684
rect 145666 575548 145818 575574
rect 140021 574848 140055 575302
rect 140021 574528 140492 574848
rect 140021 574059 140055 574528
rect 141337 574059 141371 575302
rect 141411 574059 141445 575302
rect 141525 574059 141570 575302
rect 141995 574059 142040 575302
rect 142109 574970 142146 575302
rect 142109 574059 142143 574970
rect 142807 574532 142822 574742
rect 142835 574504 142850 574770
rect 142807 574059 142822 574424
rect 142835 574059 142878 574480
rect 143499 574059 143533 575444
rect 143576 574878 143578 575302
rect 143626 574064 144999 575444
rect 145726 575116 145818 575548
rect 146196 575358 146230 576582
rect 146298 576544 147872 576582
rect 148486 576576 148554 576582
rect 148578 576548 148582 576582
rect 148584 576632 148618 576684
rect 149222 576654 149226 576678
rect 148584 576584 148630 576632
rect 149200 576616 149238 576654
rect 149342 576632 149380 576654
rect 149330 576616 149388 576632
rect 149858 576616 149896 576654
rect 148632 576584 149238 576616
rect 149290 576584 149896 576616
rect 148584 576582 149238 576584
rect 149278 576582 149896 576584
rect 148584 576576 148702 576582
rect 149278 576576 149298 576582
rect 148584 576544 148630 576576
rect 149330 576544 149388 576582
rect 146310 576420 147871 576544
rect 147901 576532 147957 576543
rect 148559 576532 148572 576543
rect 148584 576532 148618 576544
rect 149242 576543 149268 576544
rect 149217 576532 149268 576543
rect 146272 576412 147871 576420
rect 146272 576272 147904 576412
rect 146310 576264 147904 576272
rect 146310 575510 147871 576264
rect 146348 575498 147830 575510
rect 147912 575498 147957 576532
rect 148570 575510 148618 576532
rect 149228 576528 149268 576532
rect 148570 575498 148604 575510
rect 149228 575498 149262 576528
rect 149342 575510 149376 576544
rect 149875 576532 149920 576543
rect 149886 575498 149920 576532
rect 146334 575460 147836 575498
rect 147850 575460 148474 575498
rect 148556 575460 148604 575498
rect 149216 575460 149274 575498
rect 149314 575460 149352 575498
rect 149874 575460 149932 575498
rect 146348 575426 147836 575460
rect 147888 575426 148604 575460
rect 148630 575426 148638 575460
rect 148646 575426 149352 575460
rect 149404 575426 149932 575460
rect 146348 575358 147830 575426
rect 147900 575410 147958 575426
rect 148558 575410 148604 575426
rect 149216 575410 149274 575426
rect 149874 575410 149932 575426
rect 147912 575358 147946 575392
rect 148570 575358 148604 575410
rect 149917 575395 149932 575410
rect 149228 575358 149262 575392
rect 149886 575358 149920 575392
rect 150000 575358 150034 576684
rect 150571 575358 154195 576749
rect 154648 575510 154682 578282
rect 156164 576718 156198 578290
rect 156858 576728 156892 579068
rect 156922 576738 156926 579068
rect 156934 577994 156956 579068
rect 156972 577994 157017 579068
rect 157630 577994 157668 579068
rect 157676 577994 157725 579068
rect 156934 577100 156962 577994
rect 156966 577526 157017 577994
rect 156966 577100 157006 577526
rect 157624 577134 157670 577994
rect 157674 577526 157725 577994
rect 158288 578672 158333 579068
rect 158438 578672 158483 579068
rect 158618 578672 158652 579068
rect 158720 578708 158792 579068
rect 158946 578691 158991 579068
rect 159196 578691 159241 579068
rect 159604 578691 159649 579068
rect 159954 578691 159999 579068
rect 160262 578691 160307 579068
rect 160376 578691 160410 579068
rect 160712 578693 160757 579068
rect 161470 578693 161515 579068
rect 162178 578908 162212 579068
rect 162228 578908 162273 579068
rect 162292 579060 162337 579068
rect 162950 579060 163031 579068
rect 162316 579010 162960 579048
rect 162354 578976 162960 579010
rect 162986 578908 163031 579060
rect 163064 578908 163098 579068
rect 162178 578874 163098 578908
rect 163368 578908 163402 579068
rect 163482 579060 163527 579068
rect 163744 579048 163789 579068
rect 164140 579060 164185 579068
rect 163506 579010 164150 579048
rect 163544 578976 164150 579010
rect 163732 578960 163790 578976
rect 163744 578908 163789 578960
rect 164254 578908 164288 579068
rect 163368 578874 164288 578908
rect 162228 578693 162273 578874
rect 162986 578693 163031 578874
rect 163634 578764 163692 578766
rect 163634 578708 163692 578738
rect 163744 578693 163789 578874
rect 163816 578764 163900 578766
rect 163816 578708 163900 578738
rect 164502 578693 164547 579068
rect 160700 578692 160701 578693
rect 160712 578692 160758 578693
rect 161458 578692 161459 578693
rect 161470 578692 161516 578693
rect 162216 578692 162217 578693
rect 162228 578692 162274 578693
rect 162974 578692 162975 578693
rect 162986 578692 163032 578693
rect 163732 578692 163733 578693
rect 163744 578692 163790 578693
rect 164490 578692 164491 578693
rect 164502 578692 164548 578693
rect 160699 578691 160700 578692
rect 158793 578680 160700 578691
rect 160712 578680 160746 578692
rect 160758 578691 160759 578692
rect 161457 578691 161458 578692
rect 160758 578680 161458 578691
rect 161470 578680 161504 578692
rect 161516 578691 161517 578692
rect 162215 578691 162216 578692
rect 161516 578680 162216 578691
rect 162228 578680 162262 578692
rect 162274 578691 162275 578692
rect 162973 578691 162974 578692
rect 162274 578680 162974 578691
rect 162986 578680 163020 578692
rect 163032 578691 163033 578692
rect 163731 578691 163732 578692
rect 163032 578680 163732 578691
rect 163744 578680 163778 578692
rect 163790 578691 163791 578692
rect 164489 578691 164490 578692
rect 163790 578680 164490 578691
rect 164502 578680 164536 578692
rect 164548 578691 164549 578692
rect 164678 578691 164712 579068
rect 164792 578691 164837 579068
rect 164861 578691 168485 579068
rect 164548 578680 168485 578691
rect 158804 578672 168485 578680
rect 158288 578646 168485 578672
rect 158288 578566 159040 578646
rect 159196 578566 159241 578646
rect 159604 578566 159649 578646
rect 159954 578566 159999 578646
rect 160262 578566 160307 578646
rect 160376 578566 160410 578646
rect 160712 578566 160746 578646
rect 161470 578566 161504 578646
rect 162228 578566 162262 578646
rect 162986 578566 163020 578646
rect 163744 578566 163778 578646
rect 164502 578566 164536 578646
rect 164678 578566 164712 578646
rect 164792 578566 164837 578646
rect 164861 578566 168485 578646
rect 158288 578532 168485 578566
rect 169050 578538 169084 579068
rect 158288 578114 159040 578532
rect 158288 577526 158333 578114
rect 157674 577134 157714 577526
rect 156934 576842 156956 577100
rect 156972 576880 157006 577100
rect 157630 576880 157664 577134
rect 156972 576864 156990 576880
rect 157646 576872 157664 576880
rect 157676 576872 157714 577134
rect 158288 576880 158322 577526
rect 157624 576868 157670 576872
rect 157674 576868 157714 576872
rect 158326 576868 158328 577526
rect 156938 576830 156956 576842
rect 156994 576762 156996 576864
rect 157022 576790 157024 576836
rect 157602 576830 157640 576868
rect 157646 576864 157664 576868
rect 157674 576864 157726 576868
rect 157658 576830 157726 576864
rect 158260 576830 158298 576868
rect 157034 576796 157640 576830
rect 157676 576796 158298 576830
rect 157676 576780 157726 576796
rect 158310 576790 158322 576864
rect 158382 576836 158384 577994
rect 158438 577526 158483 578114
rect 158946 578094 158991 578114
rect 159196 578094 159241 578532
rect 159604 578148 159649 578532
rect 159954 578444 159999 578532
rect 159954 578358 160052 578444
rect 159954 578148 159999 578358
rect 158760 578060 159308 578094
rect 158760 577778 158794 578060
rect 158946 577991 158991 578060
rect 158824 577936 158934 577974
rect 158862 577902 158934 577936
rect 158946 577946 159133 577991
rect 159196 577974 159241 578060
rect 158946 577903 158991 577946
rect 159134 577936 159241 577974
rect 158946 577858 159133 577903
rect 159172 577902 159241 577936
rect 158946 577778 158991 577858
rect 159196 577778 159241 577902
rect 159274 577778 159308 578060
rect 158760 577744 159308 577778
rect 159358 577968 159999 578148
rect 159358 577882 160052 577968
rect 158946 577618 158991 577744
rect 159196 577618 159241 577744
rect 159358 577686 159999 577882
rect 159398 577672 159720 577686
rect 159954 577672 159999 577686
rect 158760 577584 159308 577618
rect 158438 576868 158472 577526
rect 158760 577302 158794 577584
rect 158946 577538 158991 577584
rect 158896 577526 159172 577538
rect 159196 577526 159241 577584
rect 158946 577504 158980 577526
rect 159122 577504 159133 577515
rect 158930 577498 159138 577504
rect 159196 577498 159230 577526
rect 158824 577460 158896 577498
rect 158930 577494 159234 577498
rect 158930 577492 159240 577494
rect 158862 577426 158896 577460
rect 158946 577470 159133 577492
rect 158946 577416 158980 577470
rect 159134 577460 159240 577492
rect 159122 577416 159133 577427
rect 159172 577426 159240 577460
rect 158946 577382 159133 577416
rect 158946 577302 158980 577382
rect 159196 577302 159230 577426
rect 159274 577302 159308 577584
rect 158760 577268 159308 577302
rect 158946 576880 158980 577268
rect 159196 576868 159230 577268
rect 159358 577248 159999 577672
rect 160262 577526 160307 578532
rect 159358 577210 159996 577248
rect 159604 576880 159638 577210
rect 159954 576868 159988 577210
rect 160262 576880 160296 577526
rect 158338 576830 158384 576836
rect 158426 576830 158484 576868
rect 158918 576830 158956 576868
rect 159184 576830 159242 576868
rect 159576 576830 159614 576868
rect 159942 576830 160000 576868
rect 160234 576830 160272 576868
rect 158338 576796 158956 576830
rect 159008 576796 159614 576830
rect 159666 576796 160272 576830
rect 158338 576790 158378 576796
rect 158282 576734 158322 576790
rect 158426 576780 158484 576796
rect 159184 576780 159242 576796
rect 159942 576780 160000 576796
rect 158438 576728 158472 576780
rect 160376 576728 160410 578532
rect 156858 576718 160410 576728
rect 155678 576694 160410 576718
rect 155678 576684 159230 576694
rect 155678 575358 155712 576684
rect 156164 576654 156198 576684
rect 157056 576654 157080 576684
rect 158438 576654 158472 576684
rect 155816 576616 156460 576654
rect 156474 576616 157118 576654
rect 157132 576616 157776 576654
rect 157790 576616 158434 576654
rect 155854 576582 156460 576616
rect 156512 576582 157118 576616
rect 157170 576582 157776 576616
rect 156152 576544 156210 576582
rect 156910 576544 156968 576582
rect 157024 576576 157056 576582
rect 157668 576576 157750 576582
rect 157816 576576 157818 576584
rect 157828 576582 158434 576616
rect 158438 576582 159092 576654
rect 158346 576576 158396 576582
rect 155781 576532 155837 576543
rect 155792 576226 155837 576532
rect 156164 576226 156209 576544
rect 156439 576532 156495 576543
rect 156450 576226 156495 576532
rect 156922 576226 156967 576544
rect 157000 576528 157024 576576
rect 157056 576528 157080 576576
rect 157668 576544 157726 576576
rect 157097 576532 157153 576543
rect 157108 576226 157153 576532
rect 157680 576226 157725 576544
rect 157760 576543 157776 576544
rect 157790 576543 157806 576544
rect 157755 576532 157811 576543
rect 157760 576528 157811 576532
rect 157818 576528 157834 576572
rect 158340 576528 158346 576576
rect 158413 576532 158426 576543
rect 158438 576532 158814 576582
rect 159071 576532 159127 576543
rect 157766 576226 157811 576528
rect 158424 576440 158814 576532
rect 158400 576352 158814 576440
rect 158424 576226 158483 576352
rect 159082 576226 159127 576532
rect 155792 575498 155826 576226
rect 156164 575510 156198 576226
rect 156450 575498 156484 576226
rect 156922 575510 156956 576226
rect 157108 575498 157142 576226
rect 157680 575510 157714 576226
rect 157766 575498 157800 576226
rect 158424 575510 158472 576226
rect 158424 575498 158458 575510
rect 159082 575498 159116 576226
rect 155780 575460 155838 575498
rect 156136 575460 156174 575498
rect 156438 575460 156496 575498
rect 156894 575460 156932 575498
rect 157096 575460 157154 575498
rect 157652 575460 157690 575498
rect 157754 575460 157812 575498
rect 158410 575460 158458 575498
rect 159070 575460 159128 575498
rect 155780 575426 156174 575460
rect 156226 575426 156932 575460
rect 156984 575426 157690 575460
rect 157742 575426 158458 575460
rect 158484 575426 158492 575460
rect 158500 575426 159128 575460
rect 159162 575426 159184 575460
rect 155780 575410 155838 575426
rect 156438 575410 156496 575426
rect 157096 575410 157154 575426
rect 157754 575410 157812 575426
rect 158412 575410 158458 575426
rect 159070 575410 159128 575426
rect 155780 575395 155795 575410
rect 155792 575358 155826 575392
rect 156450 575358 156484 575392
rect 157108 575358 157142 575392
rect 157766 575358 157800 575392
rect 158424 575358 158458 575410
rect 159113 575395 159128 575410
rect 159082 575358 159116 575392
rect 159196 575358 159230 576684
rect 163744 575510 163778 578532
rect 164678 578316 164712 578532
rect 164792 578468 164837 578532
rect 164861 578456 168485 578532
rect 164816 578418 168485 578456
rect 164854 578384 168485 578418
rect 164861 578316 168485 578384
rect 164678 578282 168485 578316
rect 164861 577576 168485 578282
rect 169016 577754 169028 578538
rect 169044 577754 169084 578538
rect 168512 577584 168834 577588
rect 169050 577576 169084 577754
rect 169094 577576 169139 579068
rect 169148 578990 169182 579068
rect 169306 579058 169378 579068
rect 169464 578990 169498 579068
rect 169148 578956 169498 578990
rect 169752 578924 169796 579068
rect 169798 578924 169853 579068
rect 169740 578838 169853 578924
rect 169752 578778 169796 578838
rect 169142 577976 169162 578176
rect 169198 578066 169316 578136
rect 169198 578014 169622 578066
rect 169300 577576 169622 578014
rect 169662 577754 169714 578778
rect 169718 578538 169796 578778
rect 169718 577754 169742 578538
rect 169752 577576 169796 578538
rect 169798 577576 169853 578838
rect 169968 577576 170002 579068
rect 170082 577576 170127 579068
rect 170410 577576 170455 579068
rect 170524 577576 170558 579068
rect 170566 577576 170611 579068
rect 170642 577754 170662 579068
rect 170698 577754 170718 579068
rect 170740 577576 170785 579068
rect 171324 578546 171369 579068
rect 170792 577584 171042 577588
rect 164861 576682 171030 577576
rect 171290 577272 171314 578546
rect 159246 575460 159292 575466
rect 159242 575442 159292 575460
rect 159242 575426 159280 575442
rect 159246 575420 159280 575426
rect 164861 575358 168485 576682
rect 168978 576330 168992 576534
rect 169006 576302 169020 576534
rect 169050 575510 169084 576682
rect 169124 576348 169130 576534
rect 169152 576376 169158 576534
rect 169690 575466 169714 576534
rect 169718 575466 169742 576534
rect 169808 575510 169842 576682
rect 169830 575392 169856 575494
rect 169858 575420 169884 575466
rect 169968 575460 170002 576682
rect 170082 576226 170127 576682
rect 170566 576226 170611 576682
rect 170082 575524 170116 576226
rect 170566 575512 170600 576226
rect 170642 575524 170662 576534
rect 170698 575512 170718 576534
rect 170740 576226 170785 576682
rect 170740 575524 170774 576226
rect 171262 575758 171314 577272
rect 171290 575540 171314 575758
rect 171318 577526 171369 578546
rect 171398 577526 171443 579068
rect 171458 578490 171494 579068
rect 171318 577216 171364 577526
rect 171398 577216 171438 577526
rect 171458 577216 171466 578490
rect 172056 577526 172127 579068
rect 172292 577540 172614 578048
rect 171318 575814 171370 577216
rect 171398 575814 171432 577216
rect 171318 575512 171364 575814
rect 171398 575524 171438 575814
rect 171430 575512 171438 575524
rect 171458 575512 171466 575814
rect 172056 575524 172116 577526
rect 172352 577366 172504 577540
rect 172714 577526 172759 579068
rect 172840 577526 172885 579068
rect 172160 575722 172162 577112
rect 172188 575694 172190 577140
rect 172714 575524 172748 577526
rect 172778 575778 172786 576686
rect 172082 575512 172116 575524
rect 172840 575512 172874 577526
rect 170106 575498 170750 575512
rect 170764 575498 171408 575512
rect 171422 575498 172066 575512
rect 172082 575510 172724 575512
rect 172080 575508 172724 575510
rect 172078 575498 172724 575508
rect 172738 575498 172886 575512
rect 170566 575494 170600 575498
rect 170698 575480 170718 575498
rect 171324 575494 171358 575498
rect 171458 575484 171466 575498
rect 172082 575494 172116 575498
rect 172840 575494 172874 575498
rect 172102 575480 172112 575494
rect 171290 575474 171382 575480
rect 172102 575474 172150 575480
rect 172778 575474 172840 575480
rect 172954 575474 172988 579068
rect 173386 576749 173412 577076
rect 175045 576814 175079 579532
rect 175159 576880 175193 579532
rect 175140 576814 175214 576880
rect 170144 575460 170712 575474
rect 170802 575460 171404 575474
rect 171460 575460 172028 575474
rect 172102 575460 172686 575474
rect 172776 575460 172988 575474
rect 169968 575440 171370 575460
rect 169968 575426 170538 575440
rect 170628 575426 171296 575440
rect 171386 575426 172054 575460
rect 172068 575426 172070 575460
rect 169968 575410 170002 575426
rect 172102 575424 172112 575460
rect 172118 575440 172988 575460
rect 172144 575434 172812 575440
rect 172144 575426 172824 575434
rect 172784 575420 172824 575426
rect 172840 575422 172852 575434
rect 172954 575424 172988 575440
rect 172954 575413 172965 575424
rect 172977 575413 172988 575424
rect 173005 576713 173556 576749
rect 174084 576740 174170 576772
rect 174976 576740 175214 576814
rect 173748 576713 175230 576740
rect 175521 576713 175555 581270
rect 175635 580964 175680 581270
rect 175626 580930 175680 580964
rect 175696 580930 175724 581270
rect 175817 580930 175862 581270
rect 176293 580930 176338 582032
rect 176354 580930 176382 582806
rect 176410 580930 176438 582806
rect 176475 582032 176509 582806
rect 176475 580930 176520 582032
rect 176951 580930 176985 582806
rect 177016 580930 177044 582806
rect 177072 580930 177100 582806
rect 177133 580930 177167 582806
rect 175564 580896 177167 580930
rect 175564 579598 175598 580896
rect 175635 580890 175680 580896
rect 175696 580890 175724 580896
rect 175635 580875 175724 580890
rect 175817 580875 175862 580896
rect 176293 580890 176338 580896
rect 176354 580890 176382 580896
rect 176293 580875 176382 580890
rect 176410 580875 176438 580896
rect 176475 580875 176520 580896
rect 176951 580875 176985 580896
rect 175635 580834 176768 580875
rect 176951 580862 176998 580875
rect 176951 580844 177000 580862
rect 175635 580788 175680 580834
rect 175693 580828 176342 580834
rect 176351 580828 176768 580834
rect 176939 580828 177000 580844
rect 175700 580788 175724 580828
rect 175728 580794 176342 580828
rect 175728 580788 175752 580794
rect 175635 580744 175724 580788
rect 175635 580504 175742 580744
rect 175635 579747 175724 580504
rect 175752 580476 175770 580772
rect 175817 579747 175862 580794
rect 176281 580788 176338 580794
rect 176358 580788 176382 580828
rect 176386 580794 177000 580828
rect 176386 580788 176438 580794
rect 176281 580747 176382 580788
rect 176293 580714 176382 580747
rect 176293 579747 176327 580714
rect 176336 580020 176382 580714
rect 176410 580076 176438 580788
rect 176475 580714 176520 580794
rect 176939 580747 176985 580794
rect 177016 580751 177044 580896
rect 176951 580746 176985 580747
rect 176994 580746 177044 580751
rect 176951 580744 177044 580746
rect 177072 580800 177100 580896
rect 177108 580868 177167 580896
rect 177108 580800 177176 580868
rect 177072 580744 177176 580800
rect 176951 580735 177066 580744
rect 176410 580020 176454 580076
rect 176336 579759 176398 580020
rect 176330 579752 176398 579759
rect 176410 579752 176426 580020
rect 176330 579747 176382 579752
rect 175635 579706 175874 579747
rect 175635 579660 175680 579706
rect 175693 579700 175874 579706
rect 176281 579706 176382 579747
rect 176410 579706 176454 579752
rect 176281 579700 176342 579706
rect 175700 579660 175724 579700
rect 175728 579666 176342 579700
rect 175728 579660 175752 579666
rect 175635 579632 175724 579660
rect 175626 579604 175724 579632
rect 175626 579598 175680 579604
rect 175696 579598 175724 579604
rect 175817 579598 176266 579666
rect 176281 579650 176327 579666
rect 176358 579660 176382 579706
rect 176386 579700 176454 579706
rect 176475 579747 176509 580714
rect 176951 579747 176985 580735
rect 176994 580396 177066 580735
rect 177072 580396 177094 580744
rect 177108 580396 177176 580744
rect 176994 579747 177044 580396
rect 176475 579700 176522 579747
rect 176939 579743 177044 579747
rect 176939 579734 176998 579743
rect 176939 579700 177000 579734
rect 176386 579666 177000 579700
rect 176386 579660 176438 579666
rect 176293 579620 176327 579650
rect 176330 579620 176382 579660
rect 176293 579604 176382 579620
rect 176293 579598 176338 579604
rect 176354 579598 176382 579604
rect 176410 579598 176438 579660
rect 176475 579620 176509 579666
rect 176475 579598 176520 579620
rect 176530 579598 176912 579666
rect 176939 579650 176985 579666
rect 176951 579620 176985 579650
rect 176951 579598 176996 579620
rect 177016 579598 177044 579743
rect 177072 580340 177176 580396
rect 177072 579598 177100 580340
rect 177108 579660 177176 580340
rect 177384 579680 177388 579688
rect 177108 579620 177167 579660
rect 177108 579598 177178 579620
rect 175564 579564 177178 579598
rect 175635 576713 175680 579564
rect 175696 579182 175724 579564
rect 175817 579240 176266 579564
rect 175696 576713 175724 577994
rect 175752 576713 175780 577076
rect 175817 576713 175862 579240
rect 176054 579232 176266 579240
rect 176293 579088 176338 579564
rect 176354 579182 176382 579564
rect 176410 579182 176438 579564
rect 176475 579088 176520 579564
rect 176530 579240 176912 579564
rect 176530 579232 176742 579240
rect 176951 579088 176996 579564
rect 177016 579182 177044 579564
rect 177072 579182 177100 579564
rect 177133 579088 177178 579564
rect 177396 579240 177400 579680
rect 177609 579620 177643 582806
rect 177686 580932 177714 582806
rect 177742 580932 177770 582806
rect 177791 580932 177825 582806
rect 178267 580932 178301 582806
rect 178394 580932 178422 582806
rect 178449 580932 178483 582806
rect 178563 580932 178597 582806
rect 178925 580932 178959 580966
rect 179039 580932 179073 582806
rect 177650 580898 179132 580932
rect 177650 579620 177684 580898
rect 177686 580744 177714 580898
rect 177742 580748 177770 580898
rect 177791 580830 177825 580898
rect 178267 580877 178301 580898
rect 178394 580877 178422 580898
rect 178267 580846 178314 580877
rect 178255 580830 178314 580846
rect 178394 580830 178441 580877
rect 177791 580796 178441 580830
rect 178449 580830 178483 580898
rect 178563 580830 178597 580898
rect 178925 580846 178971 580877
rect 178913 580830 178971 580846
rect 178449 580796 178971 580830
rect 177791 580748 177825 580796
rect 178255 580749 178313 580796
rect 177742 580744 177825 580748
rect 177753 580737 177825 580744
rect 177764 580488 177825 580737
rect 177609 579600 177684 579620
rect 177686 579600 177714 580488
rect 177742 579761 177825 580488
rect 177742 579600 177770 579761
rect 177791 579702 177825 579761
rect 178267 579749 178301 580749
rect 178255 579702 178314 579749
rect 178338 579708 178366 580790
rect 178394 580748 178422 580790
rect 178449 580748 178483 580796
rect 178394 579761 178483 580748
rect 178394 579749 178422 579761
rect 178394 579702 178441 579749
rect 177791 579668 178441 579702
rect 178449 579702 178483 579761
rect 178563 579702 178597 580796
rect 178913 580749 178971 580796
rect 179039 580830 179073 580898
rect 179039 580787 179068 580830
rect 178925 579749 178959 580749
rect 178913 579702 178971 579749
rect 178449 579668 178971 579702
rect 179039 579711 179073 580787
rect 179080 579745 179107 580753
rect 179754 580446 179788 583834
rect 190092 583786 190126 584874
rect 190194 583866 190228 588654
rect 191104 583866 191138 588654
rect 191206 583786 191240 588654
rect 180526 583747 180560 583751
rect 180520 583722 180560 583747
rect 181184 583722 181218 583751
rect 181842 583722 181876 583751
rect 182500 583722 182534 583751
rect 183158 583722 183192 583751
rect 190092 583724 190126 583735
rect 191206 583724 191240 583740
rect 180080 583686 183342 583722
rect 190092 583717 191240 583724
rect 191550 583717 191584 588654
rect 192080 588334 192116 588342
rect 192162 588334 192180 588342
rect 190056 583686 191601 583717
rect 191664 583686 191698 583720
rect 192122 583686 192156 583720
rect 192236 583686 192270 588654
rect 198134 588618 201770 588666
rect 203247 588665 203281 589021
rect 203361 588826 203395 589021
rect 203407 589009 203408 589010
rect 204006 589009 204007 589010
rect 203406 589008 203407 589009
rect 204007 589008 204008 589009
rect 204019 588826 204053 589021
rect 204065 589009 204066 589010
rect 204664 589009 204665 589010
rect 204064 589008 204065 589009
rect 204665 589008 204666 589009
rect 204677 588826 204711 589021
rect 204723 589009 204724 589010
rect 205322 589009 205323 589010
rect 204722 589008 204723 589009
rect 205323 589008 205324 589009
rect 205335 588826 205369 589021
rect 205381 589009 205382 589010
rect 205380 589008 205381 589009
rect 205644 588993 205725 589040
rect 205644 588814 205645 588815
rect 203991 588767 204038 588814
rect 204649 588767 204696 588814
rect 205307 588767 205354 588814
rect 205643 588813 205644 588814
rect 205691 588767 205725 588993
rect 205793 588767 205827 590451
rect 203423 588733 204038 588767
rect 204081 588733 204696 588767
rect 204739 588733 205354 588767
rect 205397 588733 205827 588767
rect 205691 588665 205725 588733
rect 205793 588665 205827 588733
rect 206765 588727 206799 599555
rect 207042 599016 207089 599654
rect 207268 599618 207302 600944
rect 218054 600936 220194 600970
rect 210352 600510 210972 600932
rect 211022 600884 211588 600918
rect 211022 600562 211056 600884
rect 211393 600804 211404 600815
rect 211077 600742 211158 600789
rect 211217 600770 211404 600804
rect 211405 600742 211486 600789
rect 211124 600704 211158 600742
rect 211452 600704 211486 600742
rect 211393 600676 211404 600687
rect 211217 600642 211404 600676
rect 211554 600562 211588 600884
rect 218597 600752 218631 600936
rect 211022 600528 211588 600562
rect 210410 600456 210428 600495
rect 210728 600467 210758 600502
rect 210784 600467 210786 600502
rect 211400 600488 211920 600502
rect 210444 600456 210462 600461
rect 210758 600456 210784 600467
rect 210352 600410 210972 600456
rect 211084 600442 211526 600476
rect 211022 600415 211588 600442
rect 210352 600408 211032 600410
rect 210352 600394 211090 600408
rect 210352 600382 210972 600394
rect 210352 600380 211004 600382
rect 210352 600347 211062 600380
rect 210352 600313 215776 600347
rect 210352 600277 210972 600313
rect 211022 600180 211062 600313
rect 211070 600186 211090 600306
rect 211124 600279 211158 600282
rect 211452 600279 211486 600282
rect 211022 600148 211056 600180
rect 211554 600148 211588 600313
rect 218042 600277 218667 600752
rect 208282 599656 209624 599692
rect 210210 599686 210428 599690
rect 210864 599656 210898 599772
rect 211040 599732 215776 599766
rect 210988 599704 211046 599722
rect 210978 599694 211012 599698
rect 210928 599668 210972 599678
rect 210978 599676 211018 599694
rect 210978 599656 211012 599676
rect 211556 599668 211778 599690
rect 207382 599618 207406 599652
rect 208282 599632 211870 599656
rect 216150 599632 216184 599772
rect 218078 599632 218112 600277
rect 219422 600256 219442 600538
rect 208282 599622 218594 599632
rect 207174 599584 207468 599618
rect 207268 599550 207302 599584
rect 207268 599482 207326 599550
rect 207400 599522 207416 599556
rect 207268 599222 207302 599482
rect 207320 599247 207336 599423
rect 207344 599247 207354 599423
rect 207370 599260 207420 599489
rect 207370 599235 207428 599260
rect 207268 599154 207326 599222
rect 207268 599086 207302 599154
rect 207372 599086 207428 599235
rect 207434 599086 207468 599584
rect 207174 599052 207468 599086
rect 207554 599584 207944 599618
rect 207554 599086 207588 599584
rect 207768 599516 207815 599563
rect 207730 599482 207815 599516
rect 207657 599423 207702 599434
rect 207785 599423 207830 599434
rect 207668 599247 207702 599423
rect 207796 599247 207830 599423
rect 207768 599188 207815 599235
rect 207730 599154 207815 599188
rect 207910 599086 207944 599584
rect 207554 599052 207944 599086
rect 207268 599002 207302 599052
rect 207372 599050 207428 599052
rect 207308 599002 207428 599050
rect 207232 598638 207482 599002
rect 207536 598638 207958 599002
rect 208282 598638 209624 599622
rect 210342 599601 218594 599622
rect 210246 599598 218594 599601
rect 207538 598564 207570 598638
rect 207572 598564 207604 598638
rect 207686 598588 207720 598598
rect 207774 598588 207808 598598
rect 207652 598554 207842 598564
rect 207412 598452 207446 598464
rect 207190 598418 207446 598452
rect 207572 598452 207606 598464
rect 207888 598452 207922 598464
rect 207572 598418 207922 598452
rect 208318 598410 208352 598638
rect 208432 598410 208466 598444
rect 209090 598410 209124 598444
rect 209748 598410 209782 598444
rect 210246 598410 210280 599598
rect 210864 599554 210898 599598
rect 210978 599585 211016 599592
rect 210966 599570 211016 599585
rect 210966 599554 211024 599570
rect 211036 599554 211074 599592
rect 211694 599554 211732 599592
rect 210468 599552 211074 599554
rect 211126 599552 211732 599554
rect 210322 599514 210342 599522
rect 210382 599520 210394 599552
rect 210452 599530 211074 599552
rect 210437 599520 211074 599530
rect 211110 599522 211732 599552
rect 211836 599522 211870 599598
rect 211104 599520 211732 599522
rect 210388 599514 210390 599520
rect 210437 599518 211058 599520
rect 211104 599518 211190 599520
rect 211638 599518 211716 599520
rect 211762 599518 211920 599522
rect 216036 599518 216070 599598
rect 216150 599518 216184 599598
rect 218078 599518 218112 599598
rect 218192 599584 218226 599598
rect 218180 599542 218238 599584
rect 218192 599538 218226 599542
rect 218220 599530 218408 599538
rect 218220 599524 218420 599530
rect 218158 599518 218420 599524
rect 210314 599482 210322 599496
rect 210406 599486 216184 599518
rect 210406 599482 210416 599486
rect 210418 599482 210420 599486
rect 210432 599484 216184 599486
rect 218044 599484 218112 599518
rect 218154 599516 218420 599518
rect 218158 599504 218420 599516
rect 218216 599494 218420 599504
rect 218216 599484 218530 599494
rect 210446 599482 211058 599484
rect 210310 599468 210382 599482
rect 210400 599472 210416 599482
rect 210446 599478 210538 599482
rect 210452 599472 210453 599473
rect 210310 599466 210388 599468
rect 210310 599456 210382 599466
rect 210348 598888 210382 599456
rect 210372 598872 210382 598888
rect 210394 598872 210440 599472
rect 210451 599471 210452 599472
rect 210446 599450 210538 599466
rect 210451 598872 210452 598873
rect 210406 598860 210440 598872
rect 210452 598871 210453 598872
rect 210864 598860 210898 599482
rect 210978 598906 211012 599482
rect 211018 599481 211058 599482
rect 211018 599478 211098 599481
rect 211104 599478 211190 599484
rect 211638 599481 211716 599484
rect 211638 599478 211756 599481
rect 211762 599478 211920 599484
rect 211053 599470 211098 599478
rect 211711 599470 211756 599478
rect 211018 599450 211058 599466
rect 211064 598894 211098 599470
rect 211104 599450 211190 599466
rect 211638 599450 211716 599466
rect 211722 598894 211756 599470
rect 211836 599466 211870 599478
rect 216023 599472 216024 599473
rect 216024 599471 216025 599472
rect 211762 599450 211870 599466
rect 211836 598954 211870 599450
rect 211836 598952 211920 598954
rect 210978 598890 211012 598894
rect 211052 598890 211110 598894
rect 211710 598890 211768 598894
rect 211836 598890 211870 598952
rect 212048 598890 212088 598898
rect 212104 598890 212116 598926
rect 216036 598906 216070 599484
rect 216036 598890 216070 598894
rect 211006 598864 216042 598890
rect 211002 598860 216046 598864
rect 216150 598860 216184 599484
rect 218078 599402 218112 599484
rect 218238 599472 218530 599484
rect 218254 599470 218530 599472
rect 218458 599402 218492 599456
rect 218560 599402 218594 599598
rect 218078 599368 218902 599402
rect 218458 598908 218492 599368
rect 218560 598908 218594 599368
rect 221344 599162 221346 600550
rect 221320 598956 221346 599162
rect 221344 598950 221346 598956
rect 221670 599682 227590 602424
rect 228059 599682 228093 603980
rect 228173 603943 228220 603959
rect 228161 603878 228220 603943
rect 228831 603928 228878 603959
rect 229489 603928 229536 603959
rect 230147 603928 230194 603959
rect 228819 603912 228878 603928
rect 229477 603912 229536 603928
rect 230135 603912 230194 603928
rect 228270 603878 228878 603912
rect 228928 603878 229536 603912
rect 229586 603878 230194 603912
rect 228161 603869 228196 603878
rect 228819 603869 228854 603878
rect 229477 603869 229512 603878
rect 230135 603869 230170 603878
rect 228161 603831 228207 603869
rect 228112 599790 228138 599906
rect 228140 599831 228166 599878
rect 228173 599831 228207 603831
rect 228208 603830 228241 603835
rect 228819 603831 228865 603869
rect 228208 601466 228242 603830
rect 228208 599843 228253 601466
rect 228262 599834 228266 600046
rect 228290 599831 228294 600074
rect 228831 599831 228865 603831
rect 228866 603830 228899 603835
rect 229477 603831 229523 603869
rect 228866 601466 228900 603830
rect 229489 602788 229523 603831
rect 229455 602120 229466 602788
rect 229483 602120 229523 602788
rect 228866 599843 228911 601466
rect 229489 600932 229523 602120
rect 229455 599866 229466 600932
rect 229483 599866 229523 600932
rect 229489 599831 229523 599866
rect 229524 603830 229557 603835
rect 230135 603831 230181 603869
rect 229524 601466 229558 603830
rect 230113 602120 230116 602788
rect 230141 602120 230144 602788
rect 229524 599843 229569 601466
rect 229582 599836 229592 600044
rect 229610 599831 229620 600072
rect 230113 599831 230116 600932
rect 230141 599831 230144 600932
rect 230147 599831 230181 603831
rect 230182 603830 230215 603835
rect 230182 601466 230216 603830
rect 230182 599843 230227 601466
rect 228140 599790 228220 599831
rect 228161 599750 228220 599790
rect 228223 599784 228878 599831
rect 228881 599784 229536 599831
rect 229539 599784 230194 599831
rect 228161 599734 228196 599750
rect 228161 599719 228176 599734
rect 228230 599716 228248 599784
rect 228258 599750 228878 599784
rect 228928 599750 229536 599784
rect 228258 599744 228276 599750
rect 228819 599734 228854 599750
rect 229477 599734 229512 599750
rect 229546 599716 229556 599784
rect 229574 599744 229584 599784
rect 229586 599750 230194 599784
rect 230135 599734 230170 599750
rect 228173 599682 228207 599716
rect 228831 599682 228865 599716
rect 229489 599682 229523 599716
rect 230147 599682 230181 599716
rect 230296 599682 230330 603980
rect 221670 599651 230330 599682
rect 230805 599651 230839 604321
rect 230945 599651 230979 604321
rect 231059 601466 231093 604321
rect 231278 602178 231280 602334
rect 231463 601466 231497 604321
rect 231059 599651 231104 601466
rect 231463 599651 231508 601466
rect 231577 599651 231611 604321
rect 232995 602808 233010 602890
rect 232288 602764 232678 602798
rect 233033 602770 233048 602928
rect 231614 602120 231624 602316
rect 232288 602266 232322 602764
rect 232375 602603 232409 602764
rect 232502 602696 232549 602743
rect 232464 602662 232549 602696
rect 232421 602603 232436 602614
rect 232519 602603 232564 602614
rect 232375 602427 232436 602603
rect 232530 602427 232564 602603
rect 232375 602404 232409 602427
rect 232375 602266 232415 602404
rect 232424 602280 232443 602376
rect 232502 602368 232549 602415
rect 232464 602334 232549 602368
rect 232644 602266 232678 602764
rect 231670 602120 231680 602260
rect 232288 602232 232678 602266
rect 232274 601562 232696 602182
rect 232999 602120 233026 602272
rect 233027 602120 233054 602300
rect 232276 600590 232282 600846
rect 232304 600618 232310 600818
rect 221670 599648 231611 599651
rect 221670 599308 227590 599648
rect 228059 599555 228093 599648
rect 228141 599617 231611 599648
rect 221670 599088 227600 599308
rect 218380 598894 218772 598908
rect 218316 598882 218772 598894
rect 218380 598866 218772 598882
rect 219446 598872 219992 598908
rect 220542 598878 220868 598908
rect 221204 598878 221534 598908
rect 210406 598856 216104 598860
rect 210310 598798 210382 598836
rect 210406 598826 216046 598856
rect 216116 598826 216184 598860
rect 218288 598860 218772 598866
rect 218288 598854 218420 598860
rect 218560 598852 218594 598860
rect 210406 598814 210440 598826
rect 210452 598814 210453 598815
rect 210348 598778 210382 598798
rect 210394 598778 210440 598814
rect 210451 598813 210452 598814
rect 210348 598414 210451 598778
rect 210864 598754 210898 598826
rect 211040 598822 216046 598826
rect 211052 598806 211110 598822
rect 211710 598814 216024 598822
rect 211710 598806 211768 598814
rect 211064 598778 211098 598806
rect 211722 598778 211756 598806
rect 211064 598754 211109 598778
rect 211722 598754 211767 598778
rect 211836 598754 211870 598814
rect 212048 598790 212088 598814
rect 212104 598800 212116 598814
rect 216150 598754 216184 598826
rect 218380 598804 218828 598852
rect 219418 598844 220020 598852
rect 220514 598850 220868 598852
rect 221204 598850 221562 598852
rect 210864 598720 216184 598754
rect 210310 598410 210451 598414
rect 211064 598410 211109 598720
rect 211722 598410 211767 598720
rect 211836 598410 211870 598720
rect 207340 598376 217592 598410
rect 208318 598296 208352 598376
rect 208432 598296 208466 598376
rect 209090 598296 209124 598376
rect 209372 598296 209736 598307
rect 209748 598296 209782 598376
rect 210246 598307 210280 598376
rect 210348 598362 210451 598376
rect 211064 598362 211109 598376
rect 211722 598362 211767 598376
rect 209794 598296 210284 598307
rect 210348 598300 210382 598362
rect 210310 598296 210382 598300
rect 210394 598296 210440 598362
rect 211064 598296 211098 598362
rect 211722 598296 211756 598362
rect 211836 598296 211870 598376
rect 217558 598320 217592 598376
rect 217406 598296 217417 598307
rect 217418 598300 217592 598320
rect 208318 598262 217417 598296
rect 208318 597838 208352 598262
rect 208432 597838 208466 598262
rect 208478 598250 208479 598251
rect 209077 598250 209078 598251
rect 208477 598249 208478 598250
rect 209078 598249 209079 598250
rect 208477 597850 208478 597851
rect 209078 597850 209079 597851
rect 208478 597849 208479 597850
rect 209077 597849 209078 597850
rect 209090 597838 209124 598262
rect 209136 598250 209137 598251
rect 209735 598250 209736 598251
rect 209748 598250 209782 598262
rect 209794 598250 209795 598251
rect 209135 598249 209136 598250
rect 209736 598249 209737 598250
rect 209748 598249 209794 598250
rect 209748 597851 209793 598249
rect 209135 597850 209136 597851
rect 209736 597850 209737 597851
rect 209748 597850 209794 597851
rect 209136 597849 209137 597850
rect 209735 597849 209736 597850
rect 209184 597838 209736 597849
rect 209748 597838 209782 597850
rect 209794 597849 209795 597850
rect 210246 597849 210280 598262
rect 210348 598256 210382 598262
rect 210314 598190 210322 598256
rect 210342 598218 210382 598256
rect 210394 598250 210440 598262
rect 210366 598214 210382 598218
rect 210366 598178 210378 598214
rect 210406 598202 210440 598250
rect 210502 598202 210538 598208
rect 210986 598202 211058 598208
rect 211064 598202 211098 598262
rect 211104 598202 211190 598208
rect 211638 598202 211674 598208
rect 211722 598202 211756 598262
rect 211836 598208 211870 598262
rect 217418 598234 217490 598272
rect 217456 598214 217490 598234
rect 211810 598202 211920 598208
rect 217418 598202 217506 598214
rect 217558 598202 217592 598300
rect 210310 598140 210382 598178
rect 210348 597922 210382 598140
rect 209794 597838 210284 597849
rect 210308 597844 210322 597922
rect 210336 597844 210382 597922
rect 210406 598168 217506 598202
rect 217524 598168 217592 598202
rect 210406 597850 210440 598168
rect 210348 597842 210382 597844
rect 210310 597838 210382 597842
rect 210394 597838 210440 597850
rect 211064 597838 211098 598168
rect 211722 597838 211756 598168
rect 211836 597838 211870 598168
rect 217418 598156 217506 598168
rect 217456 597866 217490 598156
rect 217406 597838 217417 597849
rect 208318 597804 217417 597838
rect 208318 597724 208352 597804
rect 208432 597724 208466 597804
rect 209090 597724 209124 597804
rect 209748 597724 209782 597804
rect 210246 597724 210280 597804
rect 210348 597798 210382 597804
rect 210308 597728 210322 597798
rect 210336 597754 210382 597798
rect 210394 597754 210440 597804
rect 211064 597754 211098 597804
rect 211722 597754 211756 597804
rect 210336 597728 210451 597754
rect 210308 597724 210451 597728
rect 211064 597724 211109 597754
rect 211722 597724 211767 597754
rect 211836 597724 211870 597804
rect 217558 597724 217592 598168
rect 207340 597690 217592 597724
rect 207008 595582 207058 595588
rect 207064 595582 207086 595616
rect 207008 595388 207058 595396
rect 207064 595360 207086 595396
rect 207008 592928 207058 592934
rect 207064 592928 207086 592962
rect 207008 592734 207058 592742
rect 207064 592706 207086 592742
rect 208318 591444 208352 597690
rect 209748 597226 209782 597690
rect 209436 597002 209782 597226
rect 210246 597002 210280 597690
rect 210308 597608 210322 597690
rect 210336 597636 210451 597690
rect 210314 597532 210322 597608
rect 210342 597572 210451 597636
rect 210342 597560 210388 597572
rect 210394 597557 210451 597572
rect 211064 597557 211109 597690
rect 210394 597556 210452 597557
rect 211052 597556 211053 597557
rect 211064 597556 211110 597557
rect 211710 597556 211711 597557
rect 211722 597556 211767 597690
rect 210400 597544 210440 597556
rect 210452 597555 210453 597556
rect 211051 597555 211052 597556
rect 210452 597544 211052 597555
rect 211064 597544 211098 597556
rect 211110 597555 211111 597556
rect 211709 597555 211710 597556
rect 211110 597544 211710 597555
rect 211722 597544 211756 597556
rect 211836 597544 211870 597690
rect 210400 597532 211904 597544
rect 210406 597522 211904 597532
rect 210314 597520 210322 597522
rect 210400 597520 211904 597522
rect 210310 597510 211904 597520
rect 210310 597498 210440 597510
rect 210452 597498 210453 597499
rect 211051 597498 211052 597499
rect 211064 597498 211098 597510
rect 211110 597498 211111 597499
rect 211709 597498 211710 597499
rect 211722 597498 211756 597510
rect 210310 597497 210452 597498
rect 211052 597497 211053 597498
rect 211064 597497 211110 597498
rect 211710 597497 211711 597498
rect 210310 597482 210451 597497
rect 210314 597002 210322 597482
rect 210342 597426 210451 597482
rect 210342 597002 210474 597426
rect 211064 597002 211109 597497
rect 211722 597002 211767 597498
rect 211836 597002 211870 597510
rect 208420 596968 211870 597002
rect 208432 596938 208466 596968
rect 209090 596938 209124 596968
rect 209436 596938 209782 596968
rect 210246 596938 210280 596968
rect 210314 596938 210322 596968
rect 210342 596938 210451 596968
rect 211064 596938 211109 596968
rect 211722 596938 211767 596968
rect 208432 596900 211767 596938
rect 208432 591482 208466 596900
rect 208494 596866 209124 596900
rect 209152 596866 209782 596900
rect 209810 596899 210451 596900
rect 210456 596899 211109 596900
rect 209810 596898 210452 596899
rect 210456 596898 211110 596899
rect 211114 596898 211767 596900
rect 209810 596892 210446 596898
rect 210452 596897 210453 596898
rect 210456 596897 211104 596898
rect 210452 596892 211104 596897
rect 211110 596897 211111 596898
rect 211114 596897 211756 596898
rect 209810 596886 210440 596892
rect 210452 596886 211098 596892
rect 211110 596886 211756 596897
rect 211836 596886 211870 596968
rect 209810 596866 211870 596886
rect 209056 591482 209068 591600
rect 209090 591482 209124 596866
rect 209436 596784 209782 596866
rect 209748 591482 209782 596784
rect 210246 596114 210280 596866
rect 210372 596864 210390 596866
rect 210314 596862 210390 596864
rect 210400 596862 211870 596866
rect 210310 596852 211870 596862
rect 210310 596840 210440 596852
rect 210452 596840 210453 596841
rect 211051 596840 211052 596841
rect 211064 596840 211098 596852
rect 211110 596840 211111 596841
rect 211709 596840 211710 596841
rect 211722 596840 211756 596852
rect 210310 596839 210452 596840
rect 211052 596839 211053 596840
rect 211064 596839 211110 596840
rect 211710 596839 211711 596840
rect 210310 596824 210451 596839
rect 210314 596802 210322 596824
rect 210308 596298 210322 596802
rect 210342 596774 210451 596824
rect 210336 596732 210451 596774
rect 211064 596732 211109 596839
rect 211722 596732 211767 596840
rect 210336 596326 210382 596732
rect 210314 596216 210322 596298
rect 210342 596244 210388 596326
rect 210372 596240 210382 596244
rect 210394 596240 210440 596732
rect 210451 596240 210452 596241
rect 211052 596240 211053 596241
rect 210400 596234 210440 596240
rect 210452 596239 210453 596240
rect 211051 596239 211052 596240
rect 210366 596228 210440 596234
rect 211064 596228 211098 596732
rect 211109 596240 211110 596241
rect 211710 596240 211711 596241
rect 211110 596239 211111 596240
rect 211709 596239 211710 596240
rect 211722 596228 211756 596732
rect 211836 596228 211870 596852
rect 210366 596216 211870 596228
rect 210366 596114 210378 596216
rect 210406 596194 211870 596216
rect 210406 596114 210440 596194
rect 211064 596114 211098 596194
rect 211722 596114 211756 596194
rect 211836 596114 211870 596194
rect 218560 596176 218594 598804
rect 221670 598504 227590 599088
rect 221670 598488 227630 598504
rect 221670 598240 227590 598488
rect 227630 598424 227646 598488
rect 227878 598424 227882 598504
rect 221670 598137 227591 598240
rect 227629 598176 227630 598177
rect 227630 598175 227631 598176
rect 227644 598137 227671 598180
rect 221670 598136 227590 598137
rect 221670 597816 227814 598136
rect 228045 598053 228093 599555
rect 228173 599565 228207 599617
rect 228831 599596 228865 599617
rect 229489 599596 229523 599617
rect 230147 599596 230181 599617
rect 230805 599596 230839 599617
rect 228789 599565 228865 599596
rect 229447 599565 229523 599596
rect 230105 599565 230181 599596
rect 230763 599565 230839 599596
rect 228173 599468 228219 599565
rect 228789 599549 228877 599565
rect 229447 599549 229535 599565
rect 230105 599549 230193 599565
rect 230763 599549 230851 599565
rect 230862 599555 230876 599617
rect 230945 599596 230979 599617
rect 231059 599614 231104 599617
rect 231463 599614 231508 599617
rect 231059 599596 231093 599614
rect 231463 599596 231497 599614
rect 230945 599549 230992 599596
rect 231059 599565 231106 599596
rect 231047 599549 231106 599565
rect 231421 599549 231497 599596
rect 228221 599515 228877 599549
rect 228879 599515 229535 599549
rect 229537 599515 230193 599549
rect 230195 599515 230851 599549
rect 230853 599515 231497 599549
rect 228797 599509 228801 599515
rect 228825 599481 228829 599515
rect 228831 599468 228877 599515
rect 229489 599468 229535 599515
rect 230113 599509 230117 599515
rect 230141 599481 230145 599515
rect 230147 599468 230193 599515
rect 230805 599468 230851 599515
rect 228173 599456 228207 599468
rect 228806 599456 228819 599467
rect 228831 599456 228865 599468
rect 229464 599456 229477 599467
rect 229489 599456 229523 599468
rect 230122 599456 230135 599467
rect 230147 599456 230181 599468
rect 230780 599456 230793 599467
rect 230805 599456 230839 599468
rect 228159 598152 228207 599456
rect 228817 598152 228865 599456
rect 229475 598152 229523 599456
rect 228159 598080 228193 598152
rect 228817 598140 228851 598152
rect 229475 598140 229509 598152
rect 228195 598080 228199 598127
rect 228223 598093 228227 598099
rect 228803 598093 228851 598140
rect 229461 598093 229509 598140
rect 221670 597815 227590 597816
rect 221670 597708 227591 597815
rect 227630 597776 227631 597777
rect 227629 597775 227630 597776
rect 227644 597768 227671 597815
rect 221670 596504 227590 597708
rect 210246 596080 215776 596114
rect 210366 595968 210378 596080
rect 210366 595130 210378 595830
rect 211698 595698 211790 595846
rect 211836 595698 211870 596080
rect 211302 595164 211514 595612
rect 211698 595486 211870 595698
rect 211698 595388 211790 595486
rect 211836 594597 211870 595486
rect 208432 591444 209124 591482
rect 209720 591444 209782 591482
rect 210187 594561 211906 594597
rect 215429 594561 215463 595059
rect 210187 594527 218589 594561
rect 210187 591444 211906 594527
rect 215429 594447 215463 594527
rect 215518 594476 215525 594481
rect 215571 594476 216724 594481
rect 218076 594476 218434 594481
rect 215395 594413 215463 594447
rect 215484 594453 215612 594459
rect 218394 594453 218405 594458
rect 215484 594448 216724 594453
rect 218076 594448 218406 594453
rect 215484 594447 215612 594448
rect 218394 594447 218405 594448
rect 215484 594417 218405 594447
rect 218406 594417 218487 594432
rect 215484 594413 218487 594417
rect 215429 593789 215463 594413
rect 215515 594407 216724 594413
rect 218076 594407 218487 594413
rect 215515 594401 215612 594407
rect 218406 594395 218487 594407
rect 218406 594389 218503 594395
rect 215612 594383 216724 594389
rect 218076 594383 218503 594389
rect 215608 594379 218503 594383
rect 215484 594321 215565 594368
rect 215624 594358 218503 594379
rect 215612 594343 218534 594358
rect 218406 594337 218503 594343
rect 215502 593818 215525 593823
rect 215531 593802 215565 594321
rect 215584 594315 218447 594330
rect 215880 593823 217394 593851
rect 215571 593818 218434 593823
rect 218453 593817 218487 594337
rect 218493 594315 218506 594330
rect 215484 593801 215565 593802
rect 215484 593795 215612 593801
rect 218394 593795 218405 593800
rect 215474 593790 218406 593795
rect 215395 593755 215463 593789
rect 215484 593789 215612 593790
rect 218394 593789 218405 593790
rect 215484 593759 218405 593789
rect 218406 593759 218487 593774
rect 215484 593755 218487 593759
rect 215429 593131 215463 593755
rect 215515 593749 215936 593755
rect 217338 593749 218487 593755
rect 215515 593743 215612 593749
rect 218406 593737 218487 593749
rect 218406 593731 218503 593737
rect 215612 593725 215936 593731
rect 217338 593725 218503 593731
rect 218555 593725 218589 594527
rect 215608 593721 223600 593725
rect 215484 593663 215565 593710
rect 215624 593706 223600 593721
rect 215612 593691 223600 593706
rect 215612 593685 215936 593691
rect 217338 593685 218534 593691
rect 218406 593679 218503 593685
rect 215518 593156 215525 593165
rect 215531 593144 215565 593663
rect 215584 593657 215936 593678
rect 217338 593657 218447 593678
rect 215571 593156 216754 593165
rect 218106 593156 218434 593165
rect 218453 593159 218487 593679
rect 218493 593657 218506 593678
rect 215395 593097 215463 593131
rect 215484 593143 215565 593144
rect 215484 593137 215612 593143
rect 218394 593137 218405 593142
rect 215484 593131 216754 593137
rect 218106 593131 218406 593137
rect 215484 593128 218406 593131
rect 215484 593101 218405 593128
rect 218406 593101 218487 593116
rect 215484 593097 218487 593101
rect 212290 592616 212680 592650
rect 212290 592473 212324 592616
rect 212504 592548 212551 592595
rect 212466 592514 212551 592548
rect 212450 592473 212520 592485
rect 212646 592473 212680 592616
rect 212766 592616 213156 592650
rect 212766 592473 212800 592616
rect 212980 592586 213027 592595
rect 212888 592560 213027 592586
rect 212980 592558 213027 592560
rect 212916 592532 213027 592558
rect 212942 592514 213027 592532
rect 212916 592506 212988 592507
rect 212926 592479 212996 592485
rect 212888 592478 213016 592479
rect 212926 592473 212996 592478
rect 213122 592473 213156 592616
rect 215429 592473 215463 593097
rect 215515 593091 216754 593097
rect 218106 593091 218487 593097
rect 215515 593085 215612 593091
rect 218406 593079 218487 593091
rect 218406 593073 218503 593079
rect 215612 593067 216754 593073
rect 218106 593067 218503 593073
rect 215608 593063 218503 593067
rect 215484 593005 215565 593052
rect 215624 593036 218503 593063
rect 215612 593027 218534 593036
rect 218406 593021 218503 593027
rect 215518 592486 215525 592507
rect 215531 592486 215565 593005
rect 215584 592999 218447 593008
rect 216698 592971 218162 592999
rect 215858 592507 217372 592535
rect 215571 592486 218434 592507
rect 218453 592501 218487 593021
rect 218493 592999 218506 593008
rect 212256 592439 212680 592473
rect 212732 592439 213156 592473
rect 215395 592439 215463 592473
rect 215484 592485 215565 592486
rect 215484 592479 215612 592485
rect 218394 592479 218405 592484
rect 215484 592458 218406 592479
rect 215484 592443 218405 592458
rect 218406 592443 218487 592458
rect 215484 592439 218487 592443
rect 212290 592118 212324 592439
rect 212404 592279 212438 592439
rect 212450 592427 212451 592428
rect 212519 592427 212520 592428
rect 212449 592426 212450 592427
rect 212520 592426 212521 592427
rect 212532 592279 212566 592439
rect 212386 592118 212396 592258
rect 212414 592128 212452 592230
rect 212504 592220 212551 592267
rect 212466 592186 212551 592220
rect 212646 592118 212680 592439
rect 212290 592084 212680 592118
rect 212766 592118 212800 592439
rect 212880 592279 212914 592439
rect 212926 592427 212927 592428
rect 212995 592427 212996 592428
rect 212925 592426 212926 592427
rect 212996 592426 212997 592427
rect 213008 592279 213042 592439
rect 212980 592220 213027 592267
rect 212942 592186 213027 592220
rect 213122 592118 213156 592439
rect 212766 592084 213156 592118
rect 208222 591410 209124 591444
rect 209136 591410 209782 591444
rect 209794 591410 211906 591444
rect 212272 591414 212694 592034
rect 212748 591414 213170 592034
rect 215429 591815 215463 592439
rect 215515 592433 215914 592439
rect 217316 592433 218487 592439
rect 215515 592427 215612 592433
rect 218406 592421 218487 592433
rect 218406 592415 218503 592421
rect 215612 592409 215914 592415
rect 217316 592409 218503 592415
rect 215608 592405 218503 592409
rect 215484 592347 215565 592394
rect 215624 592375 218503 592405
rect 217316 592374 218156 592375
rect 218406 592374 218503 592375
rect 215612 592369 215914 592374
rect 217316 592369 218503 592374
rect 218406 592363 218503 592369
rect 215518 591834 215525 591849
rect 215531 591828 215565 592347
rect 215584 592341 215914 592346
rect 217316 592341 218447 592346
rect 215571 591834 216748 591849
rect 218100 591834 218434 591849
rect 218453 591843 218487 592363
rect 215395 591781 215463 591815
rect 215484 591827 215565 591828
rect 215484 591821 215612 591827
rect 218394 591821 218405 591826
rect 215484 591815 216748 591821
rect 218100 591815 218406 591821
rect 215484 591806 218406 591815
rect 215484 591785 218405 591806
rect 218406 591785 218487 591800
rect 215484 591781 218487 591785
rect 215429 591637 215463 591781
rect 215515 591775 216748 591781
rect 218100 591775 218487 591781
rect 215515 591769 215612 591775
rect 218406 591763 218487 591775
rect 218406 591757 218503 591763
rect 215612 591751 216748 591757
rect 218100 591751 218503 591757
rect 215608 591747 218503 591751
rect 215624 591720 218503 591747
rect 215624 591717 218518 591720
rect 218406 591716 218518 591717
rect 215612 591711 218534 591716
rect 218406 591705 218518 591711
rect 215584 591683 218447 591688
rect 218493 591683 218506 591688
rect 216692 591655 218156 591683
rect 218555 591637 218589 593691
rect 228045 593342 228079 598053
rect 228159 597991 228199 598080
rect 228219 598080 228227 598093
rect 228235 598080 228851 598093
rect 228219 598059 228851 598080
rect 228877 598059 228885 598093
rect 228893 598059 229509 598093
rect 228223 598053 228276 598059
rect 228218 598025 228276 598052
rect 228805 598043 228851 598059
rect 229463 598043 229509 598059
rect 228218 597991 228227 598025
rect 228817 597991 228851 598043
rect 229475 597991 229509 598043
rect 229511 598025 229515 598127
rect 230056 598099 230058 599196
rect 230084 598099 230086 599168
rect 230133 598152 230181 599456
rect 230791 598152 230839 599456
rect 230862 598442 230876 599509
rect 230945 598287 230979 599515
rect 231047 599468 231105 599515
rect 231059 598448 231093 599468
rect 231463 599467 231497 599515
rect 231438 599456 231497 599467
rect 231449 598436 231497 599456
rect 231437 598389 231509 598436
rect 231121 598355 231509 598389
rect 231378 598287 231380 598342
rect 231406 598287 231408 598342
rect 231437 598339 231509 598355
rect 231449 598324 231509 598339
rect 231449 598287 231497 598324
rect 231563 598287 231611 599617
rect 232354 599192 232428 599818
rect 232340 599038 232494 599192
rect 232999 598408 233018 600932
rect 233027 598436 233046 600932
rect 233094 599692 234533 604344
rect 235876 603186 235910 604344
rect 235138 602492 235600 603130
rect 235810 603104 235910 603186
rect 235196 602408 235546 602442
rect 235196 602380 235230 602408
rect 235196 601990 235264 602380
rect 235388 602340 235426 602378
rect 235354 602306 235426 602340
rect 235299 602256 235344 602267
rect 235387 602256 235432 602267
rect 235310 602080 235344 602256
rect 235398 602080 235432 602256
rect 235388 602030 235426 602068
rect 235354 601996 235426 602030
rect 235196 601928 235230 601990
rect 235512 601928 235546 602408
rect 235196 601894 235546 601928
rect 235838 601776 235874 601862
rect 233080 599656 234533 599692
rect 234560 599656 234594 599690
rect 235218 599656 235252 599690
rect 235876 599656 235910 603104
rect 235946 602710 235948 602788
rect 235946 599656 235948 599822
rect 236016 599656 236050 604344
rect 236130 603470 236175 604344
rect 236130 599656 236164 603470
rect 236534 603444 236579 604344
rect 236534 599656 236568 603444
rect 236648 599656 236682 604344
rect 236788 599687 236822 605696
rect 237098 605084 237560 605722
rect 237574 605084 238036 605722
rect 237152 605000 237502 605034
rect 237152 604520 237186 605000
rect 237344 604932 237382 604970
rect 237310 604898 237382 604932
rect 237255 604848 237300 604859
rect 237343 604848 237388 604859
rect 237266 604672 237300 604848
rect 237354 604672 237388 604848
rect 237344 604622 237382 604660
rect 237310 604588 237382 604622
rect 237468 604520 237502 605000
rect 237152 604486 237502 604520
rect 237628 605000 237978 605034
rect 237628 604520 237662 605000
rect 237820 604932 237858 604970
rect 237786 604898 237858 604932
rect 237731 604848 237776 604859
rect 237819 604848 237864 604859
rect 237742 604672 237776 604848
rect 237830 604672 237864 604848
rect 237820 604622 237858 604660
rect 237786 604588 237858 604622
rect 237944 604520 237978 605000
rect 237628 604486 237978 604520
rect 236824 604368 236860 604454
rect 239420 599687 239454 606438
rect 233080 599622 236682 599656
rect 233080 599592 234533 599622
rect 233080 599520 234556 599592
rect 234560 599570 234594 599622
rect 235176 599588 235214 599592
rect 233080 598389 234533 599520
rect 234560 599482 234606 599570
rect 235176 599554 235216 599588
rect 234608 599520 235216 599554
rect 235172 599514 235188 599520
rect 235212 599514 235216 599520
rect 235200 599486 235216 599514
rect 235218 599570 235252 599622
rect 235218 599482 235264 599570
rect 235834 599554 235872 599592
rect 235266 599520 235872 599554
rect 235876 599570 235910 599622
rect 235876 599482 235922 599570
rect 235932 599560 235948 599622
rect 236002 599586 236004 599622
rect 235988 599560 236004 599586
rect 236016 599592 236050 599622
rect 236130 599592 236164 599622
rect 236016 599554 236054 599592
rect 236130 599570 236168 599592
rect 236118 599554 236176 599570
rect 236492 599554 236530 599592
rect 235924 599520 236530 599554
rect 234535 599470 234548 599481
rect 234560 599470 234594 599482
rect 235193 599470 235206 599481
rect 235218 599470 235252 599482
rect 235851 599470 235864 599481
rect 235876 599470 235910 599482
rect 233079 598355 234533 598389
rect 233080 598287 234533 598355
rect 230945 598253 234533 598287
rect 230133 598140 230167 598152
rect 230791 598140 230825 598152
rect 229539 598093 229543 598099
rect 230119 598093 230167 598140
rect 230777 598093 230825 598140
rect 229535 598059 229543 598093
rect 229551 598059 230167 598093
rect 230193 598059 230201 598093
rect 230209 598059 230825 598093
rect 229539 598053 229543 598059
rect 230056 598046 230058 598053
rect 230084 598018 230086 598053
rect 230121 598043 230167 598059
rect 230779 598043 230825 598059
rect 230133 597991 230167 598043
rect 230791 597991 230825 598043
rect 230827 598025 230831 598127
rect 231378 598099 231380 598253
rect 231406 598099 231408 598253
rect 231449 598152 231497 598253
rect 231449 598140 231483 598152
rect 230855 598093 230859 598099
rect 231435 598093 231483 598140
rect 230851 598059 230859 598093
rect 230867 598059 231483 598093
rect 230855 598053 230859 598059
rect 231378 598046 231380 598053
rect 231406 598018 231408 598053
rect 231437 598043 231483 598059
rect 231449 597991 231483 598043
rect 231563 598053 231611 598253
rect 233080 598217 234533 598253
rect 233116 598076 233164 598217
rect 233230 598166 233278 598217
rect 228147 597957 231495 597991
rect 228190 597824 228199 597957
rect 228218 597852 228227 597957
rect 230792 597612 230831 597957
rect 230848 597612 230859 597908
rect 231563 593342 231597 598053
rect 233116 593342 233150 598076
rect 233230 598014 233264 598166
rect 233266 598048 233270 598150
rect 233816 598122 233824 598217
rect 233844 598122 233852 598217
rect 233888 598166 233936 598217
rect 234546 598166 234594 599470
rect 235204 598166 235252 599470
rect 235280 598364 235300 598888
rect 235862 598166 235910 599470
rect 235932 598420 235948 599514
rect 235988 598378 236004 599514
rect 236016 598310 236050 599520
rect 236118 599482 236176 599520
rect 236130 598462 236164 599482
rect 236534 599481 236568 599622
rect 236509 599470 236568 599481
rect 236520 598450 236568 599470
rect 236508 598412 236580 598450
rect 236192 598378 236580 598412
rect 236444 598310 236450 598366
rect 236472 598310 236478 598366
rect 236508 598362 236580 598378
rect 236520 598347 236580 598362
rect 236520 598310 236568 598347
rect 236634 598310 236682 599622
rect 236765 599651 239604 599687
rect 239701 599651 239735 606523
rect 239815 599651 239849 606424
rect 236765 599618 240353 599651
rect 236765 599617 240378 599618
rect 236690 598910 236710 599540
rect 236765 599512 239604 599617
rect 239609 599515 239615 599549
rect 236718 599496 239604 599512
rect 236718 599234 239615 599496
rect 236718 599018 239604 599234
rect 236718 598938 239615 599018
rect 236765 598818 239615 598938
rect 236765 598796 239604 598818
rect 236690 598494 236710 598750
rect 236754 598722 239604 598796
rect 239620 598762 239674 598788
rect 236718 598618 239604 598722
rect 236718 598522 239615 598618
rect 236706 598418 236710 598494
rect 236765 598492 239615 598522
rect 236734 598418 239615 598492
rect 236765 598372 239604 598418
rect 236706 598366 236710 598372
rect 236734 598322 239604 598372
rect 236718 598310 239604 598322
rect 236016 598276 239604 598310
rect 233888 598154 233922 598166
rect 234546 598154 234580 598166
rect 235204 598154 235238 598166
rect 235862 598154 235896 598166
rect 236444 598154 236450 598276
rect 236472 598154 236478 598276
rect 236520 598166 236568 598276
rect 236520 598154 236554 598166
rect 233294 598116 233298 598122
rect 233874 598116 233922 598154
rect 234532 598116 234580 598154
rect 233290 598082 233298 598116
rect 233306 598082 233922 598116
rect 233948 598082 233956 598116
rect 233964 598082 234580 598116
rect 233294 598076 233298 598082
rect 233816 598070 233824 598076
rect 233844 598042 233852 598076
rect 233876 598066 233922 598082
rect 234534 598066 234580 598082
rect 233888 598014 233922 598066
rect 234546 598014 234580 598066
rect 234582 598048 234586 598150
rect 234610 598116 234614 598122
rect 235190 598116 235238 598154
rect 235848 598116 235896 598154
rect 234606 598082 234614 598116
rect 234622 598082 235238 598116
rect 235264 598082 235272 598116
rect 235280 598082 235896 598116
rect 234610 598076 234614 598082
rect 235192 598066 235238 598082
rect 235850 598066 235896 598082
rect 235204 598014 235238 598066
rect 235862 598014 235896 598066
rect 235898 598048 235904 598150
rect 235926 598116 235932 598122
rect 236014 598116 236554 598154
rect 235922 598082 235932 598116
rect 235938 598082 236554 598116
rect 235926 598076 235932 598082
rect 236444 598064 236450 598076
rect 236472 598042 236478 598076
rect 236508 598066 236554 598082
rect 236520 598014 236554 598066
rect 236634 598076 236682 598276
rect 236765 598240 239604 598276
rect 239701 598287 239735 599617
rect 239815 599580 239862 599596
rect 239803 599549 239862 599580
rect 239988 599584 240378 599617
rect 239988 599556 240022 599584
rect 240177 599563 240224 599584
rect 239954 599549 240056 599556
rect 240177 599549 240249 599563
rect 239803 599515 240249 599549
rect 239803 599468 239861 599515
rect 239815 598458 239849 599468
rect 239988 599086 240022 599515
rect 240164 599482 240249 599515
rect 240205 599467 240239 599472
rect 240194 599456 240239 599467
rect 240205 599439 240239 599456
rect 240205 599434 240250 599439
rect 240091 599423 240136 599434
rect 240102 599247 240136 599423
rect 240205 599247 240264 599434
rect 240205 599235 240250 599247
rect 240202 599231 240250 599235
rect 240202 599188 240249 599231
rect 240164 599154 240249 599188
rect 240205 599086 240239 599154
rect 240319 599086 240378 599584
rect 239988 599052 240378 599086
rect 240464 599584 240854 599618
rect 240464 599556 240498 599584
rect 240464 599148 240532 599556
rect 240678 599516 240725 599563
rect 240640 599482 240725 599516
rect 240567 599423 240612 599434
rect 240695 599423 240740 599434
rect 240578 599247 240612 599423
rect 240706 599247 240740 599423
rect 240678 599188 240725 599235
rect 240640 599154 240725 599188
rect 240464 599086 240498 599148
rect 240820 599086 240854 599584
rect 240464 599052 240854 599086
rect 240205 599002 240239 599052
rect 240319 599002 240353 599052
rect 239815 598448 239860 598458
rect 239970 598436 240392 599002
rect 239830 598389 240392 598436
rect 239877 598382 240392 598389
rect 240446 598382 240868 599002
rect 241755 598408 241758 600932
rect 241783 598436 241786 600932
rect 241836 599656 243289 599692
rect 244772 599656 244806 606528
rect 294434 602610 295786 602612
rect 288532 602108 288588 602124
rect 288098 601339 296074 601373
rect 241836 599622 245424 599656
rect 241836 598389 243289 599622
rect 243928 599514 243944 599542
rect 243956 599488 243972 599514
rect 244640 599486 244660 599588
rect 244668 599514 244688 599560
rect 239877 598355 240353 598382
rect 241835 598355 243289 598389
rect 240193 598339 240251 598355
rect 240205 598324 240251 598339
rect 240205 598287 240239 598324
rect 240319 598287 240353 598355
rect 241836 598287 243289 598355
rect 239701 598253 243289 598287
rect 244772 598310 244806 599622
rect 244886 599585 244924 599592
rect 244874 599570 244924 599585
rect 244874 599554 244932 599570
rect 245248 599554 245286 599592
rect 244874 599520 245286 599554
rect 244874 599482 244932 599520
rect 244886 598462 244920 599482
rect 245265 599470 245310 599481
rect 245276 598450 245310 599470
rect 245264 598412 245322 598450
rect 244948 598378 245322 598412
rect 245264 598362 245322 598378
rect 245307 598347 245322 598362
rect 245276 598310 245310 598344
rect 245390 598310 245424 599622
rect 248878 599100 248998 599120
rect 249184 599102 249424 599654
rect 249184 599100 249474 599102
rect 248872 599072 249026 599092
rect 249184 599074 249424 599100
rect 249184 599072 249502 599074
rect 249184 599016 249424 599072
rect 249813 599016 249900 599908
rect 288561 599672 292221 599705
rect 293632 599672 296240 599706
rect 259026 599100 259146 599120
rect 259332 599102 259572 599654
rect 288579 599626 292203 599672
rect 293686 599644 296240 599656
rect 293686 599638 296308 599644
rect 288579 599614 292370 599626
rect 293720 599622 296154 599638
rect 296206 599622 296308 599638
rect 288579 599592 292203 599614
rect 293686 599597 296100 599604
rect 293686 599594 293720 599597
rect 293652 599592 293754 599594
rect 284436 599560 284462 599592
rect 284866 599560 284884 599592
rect 288576 599580 292404 599592
rect 293652 599588 296104 599592
rect 259332 599100 259622 599102
rect 259020 599072 259174 599092
rect 259332 599074 259572 599100
rect 259332 599072 259650 599074
rect 259332 599016 259572 599072
rect 244772 598276 248228 598310
rect 233218 597980 236566 598014
rect 233888 593342 233922 597980
rect 236634 593342 236668 598076
rect 236877 598004 236878 598090
rect 236734 597944 236909 597964
rect 236696 597214 236744 597222
rect 236696 597180 236710 597188
rect 236915 593342 236949 598240
rect 237084 598086 237506 598240
rect 237560 598086 237982 598240
rect 239564 598184 239587 598240
rect 240205 598146 240239 598253
rect 239548 597736 239587 597964
rect 239541 597680 239587 597736
rect 239548 597418 239587 597680
rect 239541 596664 239587 597418
rect 239604 596720 239615 597908
rect 240319 593342 240353 598253
rect 241836 598217 243289 598253
rect 245390 593342 245424 598276
rect 248326 598032 248338 598314
rect 248360 598066 248372 598288
rect 257444 596664 257644 596686
rect 283690 595526 283692 595582
rect 283690 595270 283692 595326
rect 283690 595126 283692 595182
rect 283690 594870 283692 594926
rect 246034 592650 246068 593342
rect 246114 592650 246122 592840
rect 246142 592684 246150 592868
rect 246142 592650 246172 592684
rect 237088 592616 237478 592650
rect 237088 592118 237122 592616
rect 237302 592548 237349 592595
rect 237264 592514 237349 592548
rect 237191 592455 237236 592466
rect 237319 592455 237364 592466
rect 237202 592279 237236 592455
rect 237330 592279 237364 592455
rect 237302 592220 237349 592267
rect 237264 592186 237349 592220
rect 237444 592118 237478 592616
rect 237088 592084 237478 592118
rect 237564 592616 237954 592650
rect 245940 592616 246234 592650
rect 237564 592588 237598 592616
rect 237564 592180 237632 592588
rect 237778 592548 237825 592595
rect 237740 592514 237825 592548
rect 237667 592455 237712 592466
rect 237795 592455 237840 592466
rect 237678 592279 237712 592455
rect 237806 592279 237840 592455
rect 237778 592220 237825 592267
rect 237740 592186 237825 592220
rect 237564 592118 237598 592180
rect 237920 592118 237954 592616
rect 246034 592582 246068 592616
rect 246034 592514 246092 592582
rect 246034 592254 246068 592514
rect 246086 592263 246102 592471
rect 246114 592467 246122 592616
rect 246142 592521 246150 592616
rect 246166 592521 246182 592616
rect 246114 592462 246126 592467
rect 246114 592455 246120 592462
rect 246110 592279 246120 592455
rect 246114 592263 246120 592279
rect 246136 592292 246186 592521
rect 246136 592267 246194 592292
rect 246034 592186 246092 592254
rect 246034 592152 246068 592186
rect 246094 592152 246098 592228
rect 245978 592132 246098 592152
rect 246034 592124 246068 592132
rect 246122 592124 246126 592256
rect 245972 592118 246126 592124
rect 246138 592118 246194 592267
rect 246200 592118 246234 592616
rect 237564 592084 237954 592118
rect 245940 592084 246234 592118
rect 246320 592616 246710 592650
rect 246320 592118 246354 592616
rect 246534 592548 246581 592595
rect 246496 592514 246581 592548
rect 246423 592455 246468 592466
rect 246551 592455 246596 592466
rect 246434 592279 246468 592455
rect 246562 592279 246596 592455
rect 246372 592118 246392 592266
rect 246534 592220 246581 592267
rect 246496 592186 246581 592220
rect 246676 592118 246710 592616
rect 246320 592084 246710 592118
rect 278754 592616 279144 592650
rect 278754 592118 278788 592616
rect 278968 592548 279015 592595
rect 278930 592514 279015 592548
rect 278857 592455 278902 592466
rect 278985 592455 279030 592466
rect 278868 592279 278902 592455
rect 278996 592279 279030 592455
rect 278968 592220 279015 592267
rect 278930 592186 279015 592220
rect 279110 592118 279144 592616
rect 278754 592084 279144 592118
rect 279230 592616 279620 592650
rect 279230 592588 279264 592616
rect 279230 592180 279298 592588
rect 279444 592548 279491 592595
rect 279406 592514 279491 592548
rect 279333 592455 279378 592466
rect 279461 592455 279506 592466
rect 279344 592279 279378 592455
rect 279472 592279 279506 592455
rect 279444 592220 279491 592267
rect 279406 592186 279491 592220
rect 279230 592118 279264 592180
rect 279586 592118 279620 592616
rect 279230 592084 279620 592118
rect 246034 592034 246068 592084
rect 246138 592082 246194 592084
rect 246074 592034 246194 592082
rect 215429 591603 223699 591637
rect 208318 588750 208352 591410
rect 208432 591342 208466 591410
rect 209056 591346 209068 591410
rect 209090 591342 209124 591410
rect 209748 591342 209782 591410
rect 210187 591342 211906 591410
rect 208414 591308 211906 591342
rect 208432 588840 208466 591308
rect 209090 588840 209124 591308
rect 210187 591157 211906 591308
rect 210187 591123 215776 591157
rect 210187 590973 211906 591123
rect 218555 591105 218589 591603
rect 237070 591421 237492 592034
rect 236977 591387 237545 591421
rect 237546 591414 237968 592034
rect 245998 591670 246248 592034
rect 246302 591670 246724 592034
rect 246064 591620 246098 591630
rect 246452 591620 246486 591630
rect 246540 591620 246574 591630
rect 246080 591586 246132 591596
rect 246418 591586 246608 591596
rect 246046 591552 246070 591586
rect 246080 591518 246104 591586
rect 246178 591484 246212 591496
rect 245956 591450 246212 591484
rect 246338 591484 246372 591496
rect 246654 591484 246688 591496
rect 246338 591450 246688 591484
rect 278736 591421 279158 592034
rect 278643 591387 279211 591421
rect 279212 591414 279634 592034
rect 284436 591510 284462 599514
rect 284866 591510 284884 599514
rect 286278 599470 286324 599482
rect 286284 599458 286324 599470
rect 285586 597784 285598 598888
rect 286314 596174 286324 599458
rect 288579 598682 292203 599580
rect 293652 599558 293720 599588
rect 293812 599558 296104 599588
rect 296240 599570 296251 599581
rect 296263 599570 296274 599581
rect 293686 598934 293720 599558
rect 293846 599524 294468 599558
rect 294504 599524 295126 599558
rect 295162 599524 295784 599558
rect 295820 599554 296100 599558
rect 296240 599554 296274 599570
rect 295820 599524 296274 599554
rect 293862 599520 294468 599524
rect 294520 599520 295126 599524
rect 295178 599520 295784 599524
rect 295836 599520 296274 599524
rect 296099 599482 296100 599483
rect 296100 599481 296101 599482
rect 293789 599470 293834 599481
rect 294447 599470 294492 599481
rect 295105 599470 295150 599481
rect 295763 599470 295808 599481
rect 293800 598934 293834 599470
rect 293845 598946 293846 598947
rect 294446 598946 294447 598947
rect 293846 598945 293847 598946
rect 294445 598945 294446 598946
rect 294458 598934 294492 599470
rect 294503 598946 294504 598947
rect 295104 598946 295105 598947
rect 294504 598945 294505 598946
rect 295103 598945 295104 598946
rect 295116 598934 295150 599470
rect 295161 598946 295162 598947
rect 295762 598946 295763 598947
rect 295162 598945 295163 598946
rect 295761 598945 295762 598946
rect 295774 598934 295808 599470
rect 296138 598962 296172 599520
rect 295819 598946 295820 598947
rect 295820 598945 295821 598946
rect 296088 598934 296099 598945
rect 293652 598900 296099 598934
rect 288579 598470 292244 598682
rect 288579 596188 292203 598470
rect 293686 598276 293720 598900
rect 293800 598276 293834 598900
rect 293846 598888 293847 598889
rect 294445 598888 294446 598889
rect 293845 598887 293846 598888
rect 294446 598887 294447 598888
rect 293845 598288 293846 598289
rect 294446 598288 294447 598289
rect 293846 598287 293847 598288
rect 294445 598287 294446 598288
rect 294458 598276 294492 598900
rect 294504 598888 294505 598889
rect 295103 598888 295104 598889
rect 294503 598887 294504 598888
rect 295104 598887 295105 598888
rect 294503 598288 294504 598289
rect 295104 598288 295105 598289
rect 294504 598287 294505 598288
rect 295103 598287 295104 598288
rect 295116 598276 295150 598900
rect 295706 598894 295768 598900
rect 295162 598888 295163 598889
rect 295761 598888 295762 598889
rect 295161 598887 295162 598888
rect 295734 598866 295768 598888
rect 295161 598288 295162 598289
rect 295762 598288 295763 598289
rect 295162 598287 295163 598288
rect 295761 598287 295762 598288
rect 295774 598276 295808 598900
rect 295814 598894 295898 598900
rect 295820 598888 295821 598889
rect 295814 598866 295870 598888
rect 296100 598872 296172 598910
rect 296138 598304 296172 598872
rect 295819 598288 295820 598289
rect 295820 598287 295821 598288
rect 296088 598276 296099 598287
rect 293652 598242 296099 598276
rect 293686 597618 293720 598242
rect 293800 597618 293834 598242
rect 293846 598230 293847 598231
rect 294445 598230 294446 598231
rect 293845 598229 293846 598230
rect 294446 598229 294447 598230
rect 293845 597630 293846 597631
rect 293846 597629 293847 597630
rect 294374 597624 294380 597686
rect 294402 597624 294408 597658
rect 294446 597630 294447 597631
rect 294445 597629 294446 597630
rect 294458 597618 294492 598242
rect 294504 598230 294505 598231
rect 295103 598230 295104 598231
rect 294503 598229 294504 598230
rect 295104 598229 295105 598230
rect 294503 597630 294504 597631
rect 295104 597630 295105 597631
rect 294504 597629 294505 597630
rect 295103 597629 295104 597630
rect 295116 597618 295150 598242
rect 295162 598230 295163 598231
rect 295761 598230 295762 598231
rect 295161 598229 295162 598230
rect 295762 598229 295763 598230
rect 295161 597630 295162 597631
rect 295762 597630 295763 597631
rect 295162 597629 295163 597630
rect 295761 597629 295762 597630
rect 295774 597618 295808 598242
rect 295820 598230 295821 598231
rect 295819 598229 295820 598230
rect 296100 598214 296172 598252
rect 296138 597646 296172 598214
rect 295819 597630 295820 597631
rect 295820 597629 295821 597630
rect 296088 597618 296099 597629
rect 293652 597584 296099 597618
rect 293686 596960 293720 597584
rect 293800 596960 293834 597584
rect 293846 597572 293847 597573
rect 293845 597571 293846 597572
rect 294374 597494 294380 597578
rect 294402 597522 294408 597578
rect 294445 597572 294446 597573
rect 294446 597571 294447 597572
rect 293845 596972 293846 596973
rect 294446 596972 294447 596973
rect 293846 596971 293847 596972
rect 294445 596971 294446 596972
rect 294458 596960 294492 597584
rect 294504 597572 294505 597573
rect 295103 597572 295104 597573
rect 294503 597571 294504 597572
rect 295104 597571 295105 597572
rect 294503 596972 294504 596973
rect 295104 596972 295105 596973
rect 294504 596971 294505 596972
rect 295103 596971 295104 596972
rect 295116 596960 295150 597584
rect 295162 597572 295163 597573
rect 295761 597572 295762 597573
rect 295161 597571 295162 597572
rect 295762 597571 295763 597572
rect 295161 596972 295162 596973
rect 295762 596972 295763 596973
rect 295162 596971 295163 596972
rect 295761 596971 295762 596972
rect 295774 596960 295808 597584
rect 295820 597572 295821 597573
rect 295819 597571 295820 597572
rect 296100 597556 296172 597594
rect 296138 596988 296172 597556
rect 295819 596972 295820 596973
rect 295820 596971 295821 596972
rect 296088 596960 296099 596971
rect 293652 596926 296099 596960
rect 293686 596302 293720 596926
rect 293800 596302 293834 596926
rect 293846 596914 293847 596915
rect 294445 596914 294446 596915
rect 293845 596913 293846 596914
rect 294446 596913 294447 596914
rect 293845 596314 293846 596315
rect 293846 596313 293847 596314
rect 294376 596308 294380 596378
rect 294404 596308 294408 596350
rect 294446 596314 294447 596315
rect 294445 596313 294446 596314
rect 294458 596302 294492 596926
rect 294504 596914 294505 596915
rect 295103 596914 295104 596915
rect 294503 596913 294504 596914
rect 295104 596913 295105 596914
rect 294503 596314 294504 596315
rect 295104 596314 295105 596315
rect 294504 596313 294505 596314
rect 295103 596313 295104 596314
rect 295116 596302 295150 596926
rect 295162 596914 295163 596915
rect 295761 596914 295762 596915
rect 295161 596913 295162 596914
rect 295762 596913 295763 596914
rect 295161 596314 295162 596315
rect 295762 596314 295763 596315
rect 295162 596313 295163 596314
rect 295761 596313 295762 596314
rect 295774 596302 295808 596926
rect 295820 596914 295821 596915
rect 295819 596913 295820 596914
rect 296100 596898 296172 596936
rect 296138 596330 296172 596898
rect 295819 596314 295820 596315
rect 295820 596313 295821 596314
rect 296088 596302 296099 596313
rect 293652 596268 296099 596302
rect 293686 596188 293720 596268
rect 293800 596188 293834 596268
rect 294376 596188 294380 596262
rect 294404 596214 294408 596262
rect 294458 596188 294492 596268
rect 295116 596188 295150 596268
rect 295774 596188 295808 596268
rect 296240 596188 296274 599520
rect 288579 596154 296274 596188
rect 288579 596118 292203 596154
rect 292808 596118 293270 596154
rect 288615 595783 288649 596118
rect 289349 595980 289360 596066
rect 289387 595942 289398 596104
rect 292133 595783 292167 596118
rect 292844 595783 292878 596030
rect 293200 595783 293234 596030
rect 293686 595819 293720 596154
rect 293650 595783 296323 595819
rect 288017 595749 296323 595783
rect 288032 595669 288652 595749
rect 288729 595734 288763 595749
rect 288702 595700 289268 595734
rect 288702 595669 288763 595700
rect 289234 595688 289268 595700
rect 289387 595688 289421 595749
rect 288832 595669 289486 595688
rect 290045 595669 290079 595749
rect 290703 595669 290737 595749
rect 291361 595669 291395 595749
rect 292019 595669 292053 595749
rect 292133 595669 292167 595749
rect 288032 595638 292167 595669
rect 288032 595607 288652 595638
rect 288023 595568 288652 595607
rect 287950 595482 288652 595568
rect 288023 595330 288652 595482
rect 288702 595635 292167 595638
rect 288702 595605 288763 595635
rect 288775 595623 288776 595624
rect 288774 595622 288775 595623
rect 288832 595614 289486 595635
rect 290032 595623 290033 595624
rect 290033 595622 290034 595623
rect 288881 595605 289160 595614
rect 288702 595558 288838 595605
rect 288881 595601 289166 595605
rect 288897 595586 289166 595601
rect 288702 595378 288763 595558
rect 288804 595520 288838 595558
rect 288948 595520 289166 595586
rect 288948 595492 289160 595520
rect 288897 595458 289160 595492
rect 288948 595378 289160 595458
rect 289234 595378 289268 595614
rect 289349 595504 289360 595590
rect 288702 595344 289268 595378
rect 288023 595276 288057 595330
rect 288615 595276 288649 595330
rect 288023 595039 288652 595276
rect 288729 595258 288763 595344
rect 288948 595258 289160 595344
rect 288032 594854 288652 595039
rect 288702 595224 289268 595258
rect 288702 595129 288763 595224
rect 288948 595210 289160 595224
rect 289073 595144 289084 595155
rect 288702 595082 288838 595129
rect 288897 595110 289084 595144
rect 289085 595082 289166 595129
rect 288702 595011 288763 595082
rect 288804 595028 288838 595082
rect 289132 595028 289166 595082
rect 288774 595023 288775 595024
rect 288775 595022 288776 595023
rect 289073 595022 289084 595027
rect 289234 595022 289268 595224
rect 289387 595024 289432 595614
rect 289375 595023 289376 595024
rect 289387 595023 289433 595024
rect 290033 595023 290034 595024
rect 289374 595022 289375 595023
rect 288881 595016 288897 595022
rect 289073 595016 289089 595022
rect 288881 595011 289089 595016
rect 289234 595011 289375 595022
rect 289387 595011 289421 595023
rect 289433 595022 289434 595023
rect 290032 595022 290033 595023
rect 289433 595011 289458 595022
rect 290045 595011 290079 595635
rect 290091 595623 290092 595624
rect 290690 595623 290691 595624
rect 290090 595622 290091 595623
rect 290691 595622 290692 595623
rect 290090 595023 290091 595024
rect 290691 595023 290692 595024
rect 290091 595022 290092 595023
rect 290690 595022 290691 595023
rect 290703 595011 290737 595635
rect 290749 595623 290750 595624
rect 291348 595623 291349 595624
rect 290748 595622 290749 595623
rect 291349 595622 291350 595623
rect 290748 595023 290749 595024
rect 291349 595023 291350 595024
rect 290749 595022 290750 595023
rect 291348 595022 291349 595023
rect 291361 595011 291395 595635
rect 291407 595623 291408 595624
rect 292006 595623 292007 595624
rect 291406 595622 291407 595623
rect 292007 595622 292008 595623
rect 292019 595450 292053 595635
rect 292133 595450 292167 595635
rect 292844 595594 292878 595749
rect 293020 595696 293058 595703
rect 292989 595669 293105 595681
rect 292989 595666 293089 595669
rect 293004 595646 293074 595666
rect 293200 595594 293234 595749
rect 292844 595560 293234 595594
rect 292268 595478 292386 595558
rect 292242 595450 292386 595478
rect 291846 595426 292386 595450
rect 291846 595238 292294 595426
rect 291406 595023 291407 595024
rect 292007 595023 292008 595024
rect 291407 595022 291408 595023
rect 292006 595022 292007 595023
rect 292019 595011 292053 595238
rect 292133 595011 292167 595238
rect 288702 594977 292167 595011
rect 292830 595000 293252 595510
rect 292828 594977 293634 595000
rect 288702 594902 288763 594977
rect 288775 594965 288776 594966
rect 288774 594964 288775 594965
rect 289234 594902 289268 594977
rect 289374 594965 289375 594966
rect 289387 594965 289421 594977
rect 289433 594965 289434 594966
rect 290032 594965 290033 594966
rect 289375 594964 289376 594965
rect 289387 594964 289433 594965
rect 290033 594964 290034 594965
rect 288702 594868 289268 594902
rect 289387 594870 289432 594964
rect 288615 594353 288649 594854
rect 288729 594353 288763 594868
rect 288774 594365 288775 594366
rect 289375 594365 289376 594366
rect 288775 594364 288776 594365
rect 289374 594364 289375 594365
rect 289387 594353 289421 594870
rect 289432 594365 289433 594366
rect 290033 594365 290034 594366
rect 289433 594364 289434 594365
rect 290032 594364 290033 594365
rect 290045 594353 290079 594977
rect 290091 594965 290092 594966
rect 290690 594965 290691 594966
rect 290090 594964 290091 594965
rect 290691 594964 290692 594965
rect 290090 594365 290091 594366
rect 290691 594365 290692 594366
rect 290091 594364 290092 594365
rect 290690 594364 290691 594365
rect 290703 594353 290737 594977
rect 290749 594965 290750 594966
rect 291348 594965 291349 594966
rect 290748 594964 290749 594965
rect 291349 594964 291350 594965
rect 290748 594365 290749 594366
rect 291349 594365 291350 594366
rect 290749 594364 290750 594365
rect 291348 594364 291349 594365
rect 291361 594353 291395 594977
rect 291407 594965 291408 594966
rect 292006 594965 292007 594966
rect 291406 594964 291407 594965
rect 292007 594964 292008 594965
rect 291406 594365 291407 594366
rect 292007 594365 292008 594366
rect 291407 594364 291408 594365
rect 292006 594364 292007 594365
rect 292019 594353 292053 594977
rect 292133 594353 292167 594977
rect 292830 594966 293252 594977
rect 292830 594943 293600 594966
rect 292830 594890 293252 594943
rect 288581 594319 292167 594353
rect 288615 594260 288649 594319
rect 288530 594250 288723 594260
rect 288615 594232 288649 594250
rect 288502 594222 288723 594232
rect 288615 593695 288649 594222
rect 288729 593695 288763 594319
rect 288775 594307 288776 594308
rect 289374 594307 289375 594308
rect 288774 594306 288775 594307
rect 289375 594306 289376 594307
rect 288774 593707 288775 593708
rect 289375 593707 289376 593708
rect 288775 593706 288776 593707
rect 289374 593706 289375 593707
rect 289387 593695 289421 594319
rect 289433 594307 289434 594308
rect 290032 594307 290033 594308
rect 289432 594306 289433 594307
rect 290033 594306 290034 594307
rect 289432 593707 289433 593708
rect 290033 593707 290034 593708
rect 289433 593706 289434 593707
rect 290032 593706 290033 593707
rect 290045 593695 290079 594319
rect 290091 594307 290092 594308
rect 290690 594307 290691 594308
rect 290090 594306 290091 594307
rect 290691 594306 290692 594307
rect 290090 593707 290091 593708
rect 290691 593707 290692 593708
rect 290091 593706 290092 593707
rect 290690 593706 290691 593707
rect 290703 593695 290737 594319
rect 290749 594307 290750 594308
rect 291348 594307 291349 594308
rect 290748 594306 290749 594307
rect 291349 594306 291350 594307
rect 290748 593707 290749 593708
rect 291349 593707 291350 593708
rect 290749 593706 290750 593707
rect 291348 593706 291349 593707
rect 291361 593695 291395 594319
rect 291407 594307 291408 594308
rect 292006 594307 292007 594308
rect 291406 594306 291407 594307
rect 292007 594306 292008 594307
rect 291406 593707 291407 593708
rect 292007 593707 292008 593708
rect 291407 593706 291408 593707
rect 292006 593706 292007 593707
rect 292019 593695 292053 594319
rect 292133 593695 292167 594319
rect 288581 593661 292167 593695
rect 286332 591748 286356 593150
rect 288615 593037 288649 593661
rect 288729 593037 288763 593661
rect 288775 593649 288776 593650
rect 289374 593649 289375 593650
rect 288774 593648 288775 593649
rect 289375 593648 289376 593649
rect 288774 593049 288775 593050
rect 289375 593049 289376 593050
rect 288775 593048 288776 593049
rect 289374 593048 289375 593049
rect 289387 593037 289421 593661
rect 289433 593649 289434 593650
rect 290032 593649 290033 593650
rect 289432 593648 289433 593649
rect 290033 593648 290034 593649
rect 289432 593049 289433 593050
rect 290033 593049 290034 593050
rect 289433 593048 289434 593049
rect 290032 593048 290033 593049
rect 290045 593037 290079 593661
rect 290091 593649 290092 593650
rect 290690 593649 290691 593650
rect 290090 593648 290091 593649
rect 290691 593648 290692 593649
rect 290090 593049 290091 593050
rect 290691 593049 290692 593050
rect 290091 593048 290092 593049
rect 290690 593048 290691 593049
rect 290703 593037 290737 593661
rect 290749 593649 290750 593650
rect 291348 593649 291349 593650
rect 290748 593648 290749 593649
rect 291349 593648 291350 593649
rect 290748 593049 290749 593050
rect 291349 593049 291350 593050
rect 290749 593048 290750 593049
rect 291348 593048 291349 593049
rect 291361 593037 291395 593661
rect 291407 593649 291408 593650
rect 292006 593649 292007 593650
rect 291406 593648 291407 593649
rect 292007 593648 292008 593649
rect 291406 593049 291407 593050
rect 292007 593049 292008 593050
rect 291407 593048 291408 593049
rect 292006 593048 292007 593049
rect 292019 593037 292053 593661
rect 292133 593037 292167 593661
rect 288581 593003 292167 593037
rect 287574 592462 287576 592868
rect 287602 592462 287632 592840
rect 287921 592650 287955 592704
rect 287921 592618 287954 592650
rect 287887 592197 287900 592618
rect 287921 592265 287955 592618
rect 287986 592616 288376 592650
rect 287986 592265 288020 592616
rect 288023 592391 288054 592616
rect 288200 592548 288247 592595
rect 288162 592514 288247 592548
rect 288342 592484 288376 592616
rect 288088 592466 288104 592467
rect 288088 592379 288134 592466
rect 288217 592455 288262 592466
rect 288268 592462 288562 592484
rect 288342 592456 288376 592462
rect 288145 592391 288146 592392
rect 288216 592391 288217 592392
rect 288146 592390 288147 592391
rect 288215 592390 288216 592391
rect 288228 592379 288262 592455
rect 288268 592434 288534 592456
rect 288342 592379 288376 592434
rect 288615 592379 288649 593003
rect 288729 592379 288763 593003
rect 288775 592991 288776 592992
rect 289374 592991 289375 592992
rect 288774 592990 288775 592991
rect 289375 592990 289376 592991
rect 288774 592391 288775 592392
rect 289375 592391 289376 592392
rect 288775 592390 288776 592391
rect 289374 592390 289375 592391
rect 289387 592379 289421 593003
rect 289433 592991 289434 592992
rect 290032 592991 290033 592992
rect 289432 592990 289433 592991
rect 290033 592990 290034 592991
rect 289432 592391 289433 592392
rect 290033 592391 290034 592392
rect 289433 592390 289434 592391
rect 290032 592390 290033 592391
rect 290045 592379 290079 593003
rect 290091 592991 290092 592992
rect 290690 592991 290691 592992
rect 290090 592990 290091 592991
rect 290691 592990 290692 592991
rect 290090 592391 290091 592392
rect 290691 592391 290692 592392
rect 290091 592390 290092 592391
rect 290690 592390 290691 592391
rect 290703 592379 290737 593003
rect 290749 592991 290750 592992
rect 291348 592991 291349 592992
rect 290748 592990 290749 592991
rect 291349 592990 291350 592991
rect 290748 592391 290749 592392
rect 291349 592391 291350 592392
rect 290749 592390 290750 592391
rect 291348 592390 291349 592391
rect 291361 592379 291395 593003
rect 291407 592991 291408 592992
rect 292006 592991 292007 592992
rect 291406 592990 291407 592991
rect 292007 592990 292008 592991
rect 291406 592391 291407 592392
rect 292007 592391 292008 592392
rect 291407 592390 291408 592391
rect 292006 592390 292007 592391
rect 292019 592379 292053 593003
rect 292133 592379 292167 593003
rect 288088 592376 288376 592379
rect 288100 592345 288376 592376
rect 288581 592345 292167 592379
rect 288100 592319 288134 592345
rect 288228 592319 288262 592345
rect 288088 592267 288146 592319
rect 288216 592267 288274 592319
rect 288342 592265 288376 592345
rect 288615 592265 288649 592345
rect 288729 592265 288763 592345
rect 289387 592265 289421 592345
rect 290045 592265 290079 592345
rect 290703 592265 290737 592345
rect 291361 592265 291395 592345
rect 292019 592265 292053 592345
rect 292133 592265 292167 592345
rect 293650 592265 296323 595749
rect 297636 592604 298008 593308
rect 287921 592231 287954 592265
rect 287986 592231 296323 592265
rect 287986 592195 288020 592231
rect 288146 592197 288216 592220
rect 287644 592132 287764 592152
rect 287950 592134 288190 592195
rect 288342 592180 288376 592231
rect 288615 592195 288649 592231
rect 287950 592132 288240 592134
rect 287638 592104 287792 592124
rect 287950 592106 288190 592132
rect 287950 592104 288268 592106
rect 287950 592048 288190 592104
rect 288579 592048 288666 592195
rect 286284 591494 286324 591506
rect 286278 591482 286324 591494
rect 246156 591272 246160 591362
rect 246184 591288 246188 591334
rect 287092 591064 287104 591346
rect 287126 591098 287138 591320
rect 287618 591272 287632 591626
rect 288615 591381 288649 592048
rect 292133 591568 292167 592231
rect 293650 592195 296323 592231
rect 295098 592184 295172 592195
rect 298098 592048 298338 592686
rect 291526 591319 292167 591568
rect 291526 591249 292146 591319
rect 292162 591285 292167 591319
rect 292196 591285 292221 591554
rect 292196 591260 292201 591285
rect 287660 590988 287736 590990
rect 287660 590986 287732 590988
rect 210406 590534 210440 590973
rect 210498 590972 211046 590973
rect 211096 590918 211756 590973
rect 211064 590534 211098 590568
rect 211722 590534 211756 590918
rect 211836 590534 211870 590973
rect 287632 590960 287764 590962
rect 287632 590958 287760 590960
rect 219831 590716 219848 590772
rect 287624 590743 287658 590748
rect 287752 590743 287786 590748
rect 287590 590709 287692 590714
rect 287718 590709 287820 590714
rect 287890 590712 287900 590766
rect 210356 590500 215776 590534
rect 287908 590528 287936 590748
rect 287944 590564 287954 590712
rect 288130 590564 296106 590598
rect 210356 590434 210390 590500
rect 210356 588824 210394 590434
rect 210406 590396 210440 590500
rect 211064 590454 211098 590500
rect 210492 590434 211490 590454
rect 211064 590420 211098 590434
rect 211490 590420 211710 590431
rect 211722 590420 211756 590500
rect 211836 590420 211870 590500
rect 210526 590400 211870 590420
rect 210406 590358 210492 590396
rect 210542 590386 211870 590400
rect 211051 590374 211052 590375
rect 211052 590373 211053 590374
rect 210406 589740 210440 590358
rect 210442 589774 210452 590358
rect 210458 589790 210492 590358
rect 210458 589774 210474 589790
rect 211052 589774 211053 589775
rect 211051 589773 211052 589774
rect 211064 589762 211098 590386
rect 211110 590374 211111 590375
rect 211709 590374 211710 590375
rect 211109 590373 211110 590374
rect 211710 590373 211711 590374
rect 211109 589774 211110 589775
rect 211710 589774 211711 589775
rect 211110 589773 211111 589774
rect 211709 589773 211710 589774
rect 211722 589762 211756 590386
rect 211836 589762 211870 590386
rect 215084 590380 215140 590390
rect 216834 590338 217938 590362
rect 215084 590324 215140 590334
rect 216806 590310 217966 590334
rect 218670 590084 218704 590438
rect 215452 590050 223704 590084
rect 212254 589864 212716 590032
rect 212730 589864 213192 590032
rect 212092 589854 213192 589864
rect 210406 589738 210446 589740
rect 210406 589712 210492 589738
rect 210542 589728 211870 589762
rect 211051 589716 211052 589717
rect 211052 589715 211053 589716
rect 210406 589666 210498 589712
rect 210406 589650 210492 589666
rect 210406 589202 210440 589650
rect 210442 589202 210452 589650
rect 210458 589202 210492 589650
rect 210986 589636 211028 589650
rect 210406 589132 210492 589202
rect 210406 589120 210474 589132
rect 210406 589116 210452 589120
rect 210458 589116 210474 589120
rect 211052 589116 211053 589117
rect 210406 589092 210446 589116
rect 211051 589115 211052 589116
rect 211064 589104 211098 589728
rect 211110 589716 211111 589717
rect 211709 589716 211710 589717
rect 211109 589715 211110 589716
rect 211710 589715 211711 589716
rect 211136 589636 211190 589650
rect 211638 589636 211716 589650
rect 211109 589116 211110 589117
rect 211710 589116 211711 589117
rect 211110 589115 211111 589116
rect 211709 589115 211710 589116
rect 211722 589104 211756 589728
rect 211836 589104 211870 589728
rect 212254 589394 212716 589854
rect 212730 589394 213192 589854
rect 215452 589894 215486 590050
rect 218530 589970 218633 589982
rect 215638 589967 218633 589970
rect 215516 589908 215588 589946
rect 215638 589936 218618 589967
rect 218530 589924 218618 589936
rect 215452 589854 215548 589894
rect 215452 589762 215486 589854
rect 215542 589826 215548 589838
rect 215554 589774 215588 589908
rect 215594 589854 218562 589894
rect 215594 589826 218562 589838
rect 218568 589790 218602 589924
rect 218608 589854 218634 589894
rect 218608 589826 218662 589838
rect 215538 589766 215626 589774
rect 215516 589762 215626 589766
rect 218518 589762 218529 589773
rect 215418 589728 218529 589762
rect 212308 589310 212658 589344
rect 212308 589222 212342 589310
rect 212518 589282 212528 589284
rect 212500 589242 212538 589280
rect 211932 589202 212416 589222
rect 212466 589208 212538 589242
rect 211932 589196 212106 589202
rect 212308 589166 212342 589202
rect 212416 589169 212444 589170
rect 212411 589166 212456 589169
rect 212106 589146 212456 589166
rect 212499 589158 212544 589169
rect 212308 589104 212342 589146
rect 212422 589104 212456 589146
rect 212467 589116 212468 589117
rect 212498 589116 212499 589117
rect 212468 589115 212469 589116
rect 212497 589115 212498 589116
rect 212510 589104 212544 589158
rect 212624 589104 212658 589310
rect 212784 589310 213134 589344
rect 212666 589202 212740 589222
rect 212666 589146 212740 589166
rect 212784 589104 212818 589310
rect 212976 589242 213014 589280
rect 212838 589202 212892 589222
rect 212942 589208 213014 589242
rect 212892 589169 212920 589170
rect 212887 589166 212932 589169
rect 212838 589146 212932 589166
rect 212975 589158 213020 589169
rect 212898 589104 212932 589146
rect 212943 589116 212944 589117
rect 212974 589116 212975 589117
rect 212944 589115 212945 589116
rect 212973 589115 212974 589116
rect 212980 589110 213020 589158
rect 212986 589104 213020 589110
rect 213100 589104 213134 589310
rect 215452 589104 215486 589728
rect 215538 589716 215626 589728
rect 215554 589340 215588 589716
rect 218530 589700 218602 589738
rect 218568 589324 218602 589700
rect 218530 589312 218618 589324
rect 215516 589250 215588 589288
rect 215638 589278 218618 589312
rect 218530 589266 218618 589278
rect 215554 589116 215588 589250
rect 215598 589202 218562 589242
rect 215654 589146 218562 589186
rect 218568 589132 218602 589266
rect 218608 589202 218628 589242
rect 218670 589186 218704 590050
rect 287134 589566 287454 590008
rect 288462 589310 289822 589324
rect 218608 589146 218704 589186
rect 215538 589108 215626 589116
rect 215516 589104 215626 589108
rect 218518 589104 218529 589115
rect 210406 589082 210440 589092
rect 210406 589080 210446 589082
rect 210406 588986 210492 589080
rect 210542 589070 218529 589104
rect 211051 589058 211052 589059
rect 211052 589057 211053 589058
rect 210406 588843 210440 588986
rect 210442 588843 210452 588986
rect 210406 588828 210452 588843
rect 210406 588824 210440 588828
rect 210356 588756 210412 588824
rect 210458 588790 210492 588986
rect 211064 588840 211098 589070
rect 211110 589058 211111 589059
rect 211709 589058 211710 589059
rect 211109 589057 211110 589058
rect 211710 589057 211711 589058
rect 211722 588840 211756 589070
rect 210529 588828 210530 588829
rect 210530 588827 210531 588828
rect 211036 588790 211074 588828
rect 211694 588790 211732 588828
rect 210458 588756 211074 588790
rect 211126 588756 211732 588790
rect 210356 588688 210390 588756
rect 210458 588688 210492 588756
rect 211836 588688 211870 589070
rect 212308 588830 212342 589070
rect 212422 588982 212456 589070
rect 212468 589058 212469 589059
rect 212497 589058 212498 589059
rect 212467 589057 212468 589058
rect 212498 589057 212499 589058
rect 212510 588982 212544 589070
rect 212500 588932 212538 588970
rect 212466 588898 212538 588932
rect 212624 588830 212658 589070
rect 212308 588796 212658 588830
rect 212784 588830 212818 589070
rect 212898 588982 212932 589070
rect 212986 589064 213020 589070
rect 212944 589058 212945 589059
rect 212973 589058 212974 589059
rect 212943 589057 212944 589058
rect 212974 589057 212975 589058
rect 212980 588986 213020 589064
rect 212986 588982 213020 588986
rect 212976 588932 213014 588970
rect 212942 588898 213014 588932
rect 213100 588830 213134 589070
rect 212784 588796 213134 588830
rect 203247 588631 206703 588665
rect 208414 588654 211870 588688
rect 201724 588410 201736 588618
rect 201758 588444 201770 588618
rect 202142 588442 202532 588476
rect 202142 587944 202176 588442
rect 202271 588363 202403 588410
rect 202302 588351 202403 588363
rect 202318 588340 202403 588351
rect 202245 588281 202290 588292
rect 202373 588281 202418 588292
rect 202256 588105 202290 588281
rect 202384 588105 202418 588281
rect 202356 588046 202403 588093
rect 202318 588012 202403 588046
rect 202498 587944 202532 588442
rect 203992 588318 205344 588342
rect 202142 587910 202532 587944
rect 201342 587764 201750 587773
rect 201392 587754 201750 587764
rect 201794 587750 201994 587773
rect 201766 587739 202022 587745
rect 201308 587730 202022 587739
rect 201358 587722 202022 587730
rect 201358 587720 201784 587722
rect 202124 587240 202546 587860
rect 202690 587746 202950 587773
rect 202690 587718 202950 587745
rect 197616 587098 201646 587115
rect 201774 587098 202514 587115
rect 203150 587098 203962 587115
rect 205314 587098 205672 587115
rect 197644 587042 201702 587087
rect 201746 587081 202010 587087
rect 201742 587064 202548 587081
rect 203094 587042 203962 587087
rect 205314 587042 205644 587087
rect 205793 587029 205827 588631
rect 210356 587078 210390 588654
rect 215452 588584 215486 589070
rect 215538 589058 215626 589070
rect 215554 588682 215588 589058
rect 218530 589042 218602 589080
rect 218568 588666 218602 589042
rect 218530 588654 218618 588666
rect 215516 588592 215588 588630
rect 215638 588620 218618 588654
rect 218530 588608 218618 588620
rect 215452 588538 215548 588584
rect 215452 588446 215486 588538
rect 215542 588510 215548 588528
rect 215554 588458 215588 588592
rect 215594 588538 218562 588584
rect 215594 588510 218562 588528
rect 215598 588482 218562 588510
rect 218568 588474 218602 588608
rect 218608 588538 218640 588584
rect 218670 588528 218704 589146
rect 218608 588482 218704 588528
rect 215538 588450 215626 588458
rect 215516 588446 215626 588450
rect 218518 588446 218529 588457
rect 215418 588412 218529 588446
rect 210832 588370 211604 588384
rect 215452 587920 215486 588412
rect 215538 588400 215626 588412
rect 215554 588024 215588 588400
rect 218530 588384 218602 588422
rect 218568 588008 218602 588384
rect 218530 587996 218618 588008
rect 215516 587934 215588 587972
rect 215638 587962 218618 587996
rect 218530 587950 218618 587962
rect 215452 587880 215548 587920
rect 211548 587848 211604 587850
rect 211548 587748 211718 587794
rect 215452 587788 215486 587880
rect 215530 587824 215548 587864
rect 215554 587800 215588 587934
rect 215594 587880 218562 587920
rect 215594 587824 218562 587864
rect 218568 587816 218602 587950
rect 218608 587880 218644 587920
rect 218670 587864 218704 588482
rect 288328 588044 289842 588058
rect 288062 588006 288086 588028
rect 288040 587982 288086 588006
rect 296150 588006 296174 588028
rect 296150 587982 296196 588006
rect 218608 587824 218704 587864
rect 215538 587792 215626 587800
rect 215516 587788 215626 587792
rect 218518 587788 218529 587799
rect 215418 587754 218529 587788
rect 211548 587720 211718 587740
rect 215452 587130 215486 587754
rect 215538 587742 215626 587754
rect 215554 587366 215588 587742
rect 218530 587726 218602 587764
rect 218568 587350 218602 587726
rect 218530 587338 218618 587350
rect 215516 587276 215588 587314
rect 215638 587304 218618 587338
rect 218530 587292 218618 587304
rect 215508 587228 215548 587240
rect 215536 587172 215548 587212
rect 215554 587142 215588 587276
rect 215594 587228 218562 587240
rect 215594 587172 218562 587212
rect 218568 587158 218602 587292
rect 218608 587228 218640 587240
rect 218670 587212 218704 587824
rect 218608 587172 218704 587212
rect 215538 587134 215626 587142
rect 215516 587130 215626 587134
rect 218518 587130 218529 587141
rect 215418 587096 218529 587130
rect 215452 587016 215486 587096
rect 215523 587084 215626 587096
rect 218670 587016 218704 587172
rect 210452 586982 218704 587016
rect 215452 586628 215486 586982
rect 282962 586830 284142 587202
rect 219924 586730 219980 586742
rect 219924 586674 219980 586686
rect 288740 586554 288760 586612
rect 288768 586554 288788 586606
rect 214518 586478 214522 586512
rect 214552 586504 214556 586530
rect 215060 586308 215082 586314
rect 215060 586304 215078 586308
rect 215060 586248 215102 586258
rect 215157 586197 215210 586451
rect 288684 586314 289322 586554
rect 215411 586104 215464 586197
rect 216174 586148 216848 586161
rect 286412 586158 287292 586206
rect 215543 586127 216848 586148
rect 215447 585946 215481 586065
rect 215558 585985 216178 586127
rect 216228 586093 216762 586112
rect 286356 586102 287236 586150
rect 216262 586078 216760 586093
rect 215549 585946 216178 585985
rect 215447 585860 216178 585946
rect 200924 585500 200940 585530
rect 200890 585466 200906 585496
rect 215447 585463 215481 585860
rect 215549 585708 216178 585860
rect 216228 586053 216794 586059
rect 216228 586047 216262 586053
rect 216760 586047 216794 586053
rect 216228 586044 216794 586047
rect 216228 585972 216262 586044
rect 216385 586032 216637 586036
rect 216373 586013 216649 586032
rect 216599 585998 216610 586001
rect 216407 585983 216615 585998
rect 216283 585972 216364 585983
rect 216407 585979 216692 585983
rect 216228 585930 216268 585972
rect 216276 585936 216364 585972
rect 216423 585964 216610 585979
rect 216611 585936 216692 585979
rect 216276 585930 216296 585936
rect 216228 585756 216262 585930
rect 216330 585898 216364 585936
rect 216658 585898 216692 585936
rect 216599 585870 216610 585881
rect 216423 585836 216610 585870
rect 216760 585756 216794 586044
rect 288740 585982 288742 586158
rect 288768 586010 288770 586130
rect 289160 586042 289194 586114
rect 289160 586038 289190 586042
rect 289216 586014 289222 586142
rect 289216 586010 289218 586014
rect 216228 585722 216794 585756
rect 215549 585654 215583 585708
rect 215549 585463 216178 585654
rect 216228 585602 216794 585636
rect 216228 585463 216262 585602
rect 216599 585522 216610 585533
rect 216423 585497 216610 585522
rect 216407 585488 216615 585497
rect 216276 585463 216278 585482
rect 216760 585463 216794 585602
rect 289207 585486 289622 585517
rect 285654 585481 289622 585486
rect 294278 585486 294699 585517
rect 294278 585481 299638 585486
rect 210429 585430 218699 585463
rect 280583 585447 284419 585481
rect 285654 585452 299638 585481
rect 289207 585447 294699 585452
rect 210367 585429 218699 585430
rect 210367 585395 210402 585396
rect 215447 585349 215481 585429
rect 215549 585417 216178 585429
rect 215558 585387 216178 585417
rect 216228 585389 216262 585429
rect 216276 585395 216278 585429
rect 216330 585406 216364 585429
rect 216658 585423 216692 585429
rect 216650 585414 216702 585423
rect 216652 585410 216698 585414
rect 216658 585406 216692 585410
rect 216412 585401 216610 585405
rect 216423 585389 216599 585394
rect 216622 585389 216730 585395
rect 216760 585389 216794 585429
rect 216228 585387 216794 585389
rect 215558 585383 218542 585387
rect 215558 585361 218554 585383
rect 215502 585355 218554 585361
rect 215502 585349 216178 585355
rect 216228 585349 216262 585355
rect 216760 585349 216794 585355
rect 197670 585266 205646 585300
rect 210401 585210 210402 585337
rect 215413 585334 218520 585349
rect 215413 585321 218597 585334
rect 215413 585315 218515 585321
rect 210435 585210 210436 585303
rect 198916 584014 201882 584952
rect 202428 584686 204078 584956
rect 204514 584686 205868 584954
rect 208792 584778 208800 584804
rect 202428 584664 205868 584686
rect 194378 583716 194660 583740
rect 180080 583652 184048 583686
rect 190056 583681 195616 583686
rect 185289 583652 195616 583681
rect 180080 583584 183342 583652
rect 185289 583647 191601 583652
rect 183464 583590 183492 583616
rect 183634 583600 183645 583611
rect 183657 583600 183668 583611
rect 183634 583584 183668 583600
rect 180080 583550 183668 583584
rect 180080 583511 183342 583550
rect 183350 583511 183372 583516
rect 179220 580156 179228 580210
rect 179718 580192 179954 580446
rect 179714 580156 179954 580192
rect 180080 580156 183372 583511
rect 179039 579692 179068 579711
rect 177791 579620 177825 579668
rect 177791 579600 177836 579620
rect 177872 579600 178254 579668
rect 178255 579652 178313 579668
rect 178267 579620 178301 579652
rect 178267 579600 178312 579620
rect 178394 579600 178422 579662
rect 178449 579620 178483 579668
rect 178449 579600 178494 579620
rect 178518 579600 178730 579668
rect 178913 579652 178971 579668
rect 179008 579668 179068 579692
rect 179008 579666 179073 579668
rect 178956 579637 178971 579652
rect 178842 579612 178856 579618
rect 178842 579606 178919 579612
rect 178925 579600 178959 579634
rect 179039 579612 179073 579666
rect 179116 579618 179120 579662
rect 178965 579606 179120 579612
rect 179039 579600 179073 579606
rect 177609 579566 179132 579600
rect 179274 579590 179282 580156
rect 179714 580122 183372 580156
rect 179714 580054 179954 580122
rect 179964 580054 180011 580101
rect 179714 580020 180011 580054
rect 179714 579773 179954 580020
rect 179981 579961 180026 579972
rect 179992 579785 180026 579961
rect 179714 579747 180011 579773
rect 179714 579734 179954 579747
rect 179714 579716 179968 579734
rect 179714 579700 179964 579716
rect 180080 579700 183372 580122
rect 179714 579666 183372 579700
rect 177609 579088 177654 579566
rect 177686 579182 177714 579566
rect 177742 579182 177770 579566
rect 177791 579088 177836 579566
rect 177872 579232 178254 579566
rect 178267 579088 178312 579566
rect 178394 579182 178422 579566
rect 178449 579088 178494 579566
rect 178518 579456 178816 579566
rect 178518 579232 178730 579456
rect 176293 578528 176327 579088
rect 176475 578528 176509 579088
rect 176293 576713 176338 578528
rect 176354 576713 176382 577994
rect 176410 576713 176438 577994
rect 176475 576713 176520 578528
rect 176951 577604 176985 579088
rect 173005 576679 176593 576713
rect 173005 576611 173556 576679
rect 173748 576664 175230 576679
rect 175521 576664 175555 576679
rect 175635 576664 175680 576679
rect 175696 576664 175724 576679
rect 175752 576664 175780 576679
rect 175817 576664 175862 576679
rect 173748 576658 176238 576664
rect 176293 576658 176338 576679
rect 176354 576658 176382 576679
rect 176410 576658 176438 576679
rect 173748 576611 176464 576658
rect 173005 576609 175806 576611
rect 175817 576609 176464 576611
rect 173005 576577 176464 576609
rect 176475 576600 176520 576679
rect 169968 575399 169979 575410
rect 169991 575399 170002 575410
rect 173005 575372 173556 576577
rect 173748 576562 175874 576577
rect 176062 576562 176109 576577
rect 173748 576528 176109 576562
rect 173748 576112 175230 576528
rect 173694 576036 175230 576112
rect 173748 575550 175230 576036
rect 173748 575532 175280 575550
rect 173614 575498 175280 575532
rect 175521 575498 175555 576528
rect 175635 575510 175680 576528
rect 175776 576518 175862 576528
rect 175787 575510 175862 576518
rect 176079 576469 176124 576480
rect 175787 575498 175832 575510
rect 176090 575498 176124 576469
rect 173614 575451 175874 575498
rect 176078 575451 176137 575498
rect 176204 575451 176238 576577
rect 176293 575510 176327 576577
rect 176354 576256 176382 576571
rect 176346 575457 176382 576256
rect 176410 576529 176438 576571
rect 176475 576529 176509 576600
rect 176410 576518 176509 576529
rect 176410 576200 176438 576518
rect 176402 575498 176438 576200
rect 176445 575510 176509 576518
rect 176445 575498 176490 575510
rect 176402 575457 176491 575498
rect 176433 575451 176491 575457
rect 176559 575451 176593 576679
rect 176951 576600 176996 577604
rect 176951 575510 176985 576600
rect 177016 575457 177044 577994
rect 177072 575457 177100 577994
rect 177133 577604 177167 579088
rect 177609 577604 177643 579088
rect 177133 576600 177178 577604
rect 177609 576600 177654 577604
rect 177133 575510 177167 576600
rect 177609 575528 177643 576600
rect 177686 575528 177714 577994
rect 177742 575528 177770 577994
rect 177791 577604 177825 579088
rect 178267 577604 178301 579088
rect 177791 576600 177836 577604
rect 178267 576754 178312 577604
rect 178394 576754 178422 577994
rect 178449 577604 178483 579088
rect 178449 576754 178494 577604
rect 178563 576754 178597 579232
rect 179039 576754 179073 579566
rect 179260 579530 179264 579540
rect 179314 579400 179334 579636
rect 179342 579372 179362 579664
rect 179714 579658 179954 579666
rect 179410 579638 179530 579640
rect 179714 579638 180006 579658
rect 180080 579646 183372 579666
rect 180016 579638 183372 579646
rect 179714 579630 179954 579638
rect 179714 579624 180012 579630
rect 179382 579610 179558 579612
rect 179714 579598 180044 579624
rect 180080 579620 183372 579638
rect 183384 579620 183406 583550
rect 180080 579598 183383 579620
rect 179714 579564 183383 579598
rect 179714 579554 179954 579564
rect 180080 579540 183383 579564
rect 179736 579528 183383 579540
rect 180116 579408 180150 579528
rect 180258 579458 180270 579528
rect 180286 579486 180298 579528
rect 179434 579360 179510 579362
rect 179926 579360 179968 579382
rect 179406 579332 179538 579334
rect 179416 579110 179526 579130
rect 179454 579072 179488 579092
rect 180088 579052 180150 579408
rect 180260 579402 180270 579458
rect 180288 579430 180298 579486
rect 180324 579356 180362 579382
rect 180116 577974 180150 579052
rect 180592 577974 180626 579528
rect 180706 579088 180751 579528
rect 180782 579182 180810 579356
rect 180838 579182 180866 579356
rect 180888 579088 180933 579528
rect 180950 579212 181352 579528
rect 181140 579208 181352 579212
rect 181364 579088 181409 579528
rect 181434 579182 181462 579528
rect 181490 579182 181518 579528
rect 181546 579088 181591 579528
rect 181616 579212 182000 579528
rect 181616 579208 181828 579212
rect 182022 579088 182067 579528
rect 180706 577974 180740 579088
rect 180782 577974 180810 577994
rect 179280 577952 180848 577974
rect 179280 577948 180810 577952
rect 178076 576718 179109 576754
rect 180116 576718 180150 577948
rect 180592 576718 180626 577948
rect 180706 577604 180740 577948
rect 180706 576718 180751 577604
rect 180782 576718 180810 577948
rect 180888 577604 180922 579088
rect 181364 577604 181398 579088
rect 180888 576718 180933 577604
rect 181364 576718 181409 577604
rect 181434 576718 181462 577994
rect 181490 576718 181518 577994
rect 181546 577604 181580 579088
rect 182022 577604 182056 579088
rect 181546 576718 181591 577604
rect 178076 576684 181664 576718
rect 177791 575528 177825 576600
rect 178076 575528 179109 576684
rect 177478 575492 179109 575528
rect 179542 575492 179576 575526
rect 180116 575492 180150 576684
rect 180592 576654 180626 576684
rect 180706 576654 180751 576684
rect 180782 576654 180810 576684
rect 180888 576654 180933 576684
rect 181364 576654 181409 576684
rect 181434 576654 181462 576684
rect 181490 576654 181518 576684
rect 180166 576576 180184 576622
rect 180194 576548 180212 576650
rect 180226 576616 180868 576654
rect 180884 576616 181526 576654
rect 180230 576582 180868 576616
rect 180888 576582 181526 576616
rect 181546 576600 181591 576684
rect 180230 576544 180276 576582
rect 180230 576532 180264 576544
rect 180200 575508 180264 576532
rect 180200 575492 180234 575508
rect 180592 575492 180626 576582
rect 180706 575508 180740 576582
rect 180782 575492 180810 576576
rect 180888 576543 180922 576582
rect 180847 576532 180922 576543
rect 180858 575512 180922 576532
rect 180846 575508 180922 575512
rect 181364 575508 181398 576582
rect 181434 575952 181462 576576
rect 181490 576543 181518 576576
rect 181546 576543 181580 576600
rect 181490 575952 181580 576543
rect 181440 575540 181462 575952
rect 181468 575508 181580 575952
rect 180846 575492 180904 575508
rect 181468 575492 181562 575508
rect 181630 575492 181664 576684
rect 182022 576600 182067 577604
rect 182022 575508 182056 576600
rect 182092 575492 182120 579528
rect 182148 575524 182176 579528
rect 182204 579088 182249 579528
rect 182264 579212 182668 579528
rect 182456 579206 182668 579212
rect 182680 579088 182725 579528
rect 182204 577604 182238 579088
rect 182680 577604 182714 579088
rect 182204 576600 182249 577604
rect 182680 576600 182725 577604
rect 182204 575508 182238 576600
rect 182680 575508 182714 576600
rect 182756 575492 182784 579528
rect 182812 575492 182840 579528
rect 182862 579088 182907 579528
rect 182932 579206 183312 579528
rect 183100 579194 183312 579206
rect 183338 579088 183383 579528
rect 182862 577604 182896 579088
rect 183338 577604 183372 579088
rect 183384 579052 183406 579088
rect 182862 576600 182907 577604
rect 183338 576600 183383 577604
rect 182862 575524 182896 576600
rect 183338 575524 183372 576600
rect 182862 575508 182868 575524
rect 177478 575480 182840 575492
rect 183464 575480 183492 583544
rect 183509 583500 183565 583511
rect 183520 579052 183565 583500
rect 183520 577604 183554 579052
rect 183520 576600 183565 577604
rect 183520 575524 183554 576600
rect 177478 575474 182834 575480
rect 183634 575474 183668 583550
rect 185193 576970 185227 583585
rect 188013 583579 188047 583617
rect 188711 583595 188722 583606
rect 188734 583595 188745 583606
rect 188711 583579 188745 583595
rect 188013 583545 188745 583579
rect 187946 579964 187973 583502
rect 187980 579998 188007 583536
rect 185157 576814 185244 576970
rect 185288 576814 185362 576880
rect 185124 576738 185362 576814
rect 184034 576718 184042 576734
rect 184012 576700 184042 576718
rect 185157 576716 185244 576738
rect 184052 576700 184180 576716
rect 184528 576700 184768 576716
rect 185004 576700 185244 576716
rect 185288 576714 185362 576738
rect 184012 576664 184180 576700
rect 185193 576680 185227 576700
rect 185288 576680 185368 576714
rect 184184 576664 184382 576680
rect 184660 576664 184858 576680
rect 185136 576664 185430 576680
rect 184030 576630 186386 576664
rect 184030 576481 184180 576630
rect 185193 576612 185227 576630
rect 185288 576616 185362 576630
rect 185274 576612 185362 576616
rect 184214 576600 184352 576612
rect 184690 576600 184828 576612
rect 185193 576600 185362 576612
rect 184248 576566 184318 576578
rect 184264 576562 184302 576566
rect 184444 576562 184478 576600
rect 184242 576535 184478 576562
rect 184226 576528 184478 576535
rect 184366 576522 184398 576525
rect 184404 576522 184478 576528
rect 184202 576497 184236 576501
rect 184330 576497 184364 576501
rect 184190 576481 184198 576497
rect 184202 576494 184248 576497
rect 184211 576485 184248 576494
rect 184030 576469 184198 576481
rect 184202 576481 184248 576485
rect 184318 576481 184376 576497
rect 184202 576469 184236 576481
rect 184030 576309 184236 576469
rect 184330 576309 184364 576481
rect 184030 576286 184214 576309
rect 184030 576154 184220 576286
rect 184222 576182 184248 576258
rect 184302 576250 184349 576297
rect 184264 576216 184349 576250
rect 184222 576162 184342 576182
rect 184030 576148 184370 576154
rect 184404 576148 184416 576154
rect 184444 576148 184478 576522
rect 184030 576114 184478 576148
rect 184564 576562 184598 576600
rect 184724 576566 184794 576578
rect 184740 576562 184778 576566
rect 184920 576562 184954 576600
rect 184564 576528 184954 576562
rect 184564 576148 184598 576528
rect 184678 576497 184712 576501
rect 184806 576497 184840 576501
rect 184666 576481 184724 576497
rect 184794 576481 184852 576497
rect 184678 576309 184712 576481
rect 184806 576309 184840 576481
rect 184778 576250 184825 576297
rect 184740 576216 184825 576250
rect 184920 576148 184954 576528
rect 184564 576114 184954 576148
rect 185040 576148 185074 576600
rect 185193 576578 185227 576600
rect 185246 576584 185262 576588
rect 185246 576580 185266 576584
rect 185274 576580 185362 576600
rect 185193 576566 185270 576578
rect 185193 576562 185254 576566
rect 185288 576562 185362 576580
rect 185396 576609 185430 576630
rect 185959 576609 186005 576630
rect 185396 576562 185443 576609
rect 185931 576578 185954 576580
rect 185959 576578 186012 576609
rect 185931 576568 186012 576578
rect 185953 576562 186012 576568
rect 186210 576562 186257 576609
rect 185193 576535 186257 576562
rect 185120 576528 186257 576535
rect 185154 576497 185188 576501
rect 185193 576497 185227 576528
rect 185288 576501 185362 576528
rect 185282 576497 185362 576501
rect 185142 576481 185227 576497
rect 185270 576481 185362 576497
rect 185154 576309 185188 576481
rect 185159 576293 185188 576309
rect 185193 576250 185227 576481
rect 185282 576309 185362 576481
rect 185288 576297 185362 576309
rect 185254 576250 185362 576297
rect 185193 576226 185362 576250
rect 185193 576216 185301 576226
rect 185193 576148 185227 576216
rect 185307 576182 185341 576226
rect 185307 576148 185368 576182
rect 185396 576148 185430 576528
rect 185953 576522 186011 576528
rect 185040 576114 185430 576148
rect 185931 576481 186011 576522
rect 185931 576142 185954 576481
rect 185959 576142 186005 576481
rect 186227 576469 186272 576480
rect 184030 576064 184198 576114
rect 184404 576096 184416 576114
rect 184404 576064 184418 576096
rect 185193 576064 185227 576114
rect 185307 576064 185341 576114
rect 177478 575458 183968 575474
rect 177478 575451 179109 575458
rect 173614 575440 179109 575451
rect 170064 575358 173556 575372
rect 173710 575362 173716 575440
rect 173748 575417 179109 575440
rect 145826 574974 145846 575340
rect 146196 575324 154195 575358
rect 155296 575338 173556 575358
rect 155296 575324 172892 575338
rect 146348 575164 147830 575324
rect 146408 574064 146442 575164
rect 146482 574064 146516 575164
rect 146596 574064 146641 575164
rect 147066 574064 147111 575164
rect 147180 574974 147214 575164
rect 147180 574864 147232 574974
rect 147180 574064 147214 574864
rect 147254 574064 147288 575164
rect 148530 574974 148542 575324
rect 143626 574059 149932 574064
rect 138693 574030 149932 574059
rect 138693 574025 144999 574030
rect 137432 569712 137440 569766
rect 138555 569748 138642 570002
rect 137450 569110 137578 569748
rect 137588 569329 137596 569529
rect 137926 569214 138166 569748
rect 138402 569712 138642 569748
rect 138705 569712 138739 574025
rect 139363 574004 139397 574025
rect 140021 574004 140055 574025
rect 140679 574004 140713 574025
rect 141337 574004 141371 574025
rect 139335 573957 139397 574004
rect 139993 573957 140055 574004
rect 140651 573957 140713 574004
rect 141309 573957 141371 574004
rect 141411 574004 141445 574025
rect 141525 574022 141570 574025
rect 141995 574022 142040 574025
rect 141525 574004 141559 574022
rect 141995 574004 142029 574022
rect 141411 573957 141458 574004
rect 141525 573957 141572 574004
rect 141995 573957 142042 574004
rect 142109 573957 142143 574025
rect 142183 574004 142217 574025
rect 142155 573957 142217 574004
rect 142807 574004 142822 574025
rect 142835 574004 142878 574025
rect 143499 574004 143533 574025
rect 142807 573991 142878 574004
rect 143471 573991 143533 574004
rect 142807 573957 142881 573991
rect 142891 573957 142909 573963
rect 143471 573957 143548 573991
rect 143549 573957 143576 573963
rect 143626 573962 144999 574025
rect 145092 574000 145126 574030
rect 145750 574000 145784 574030
rect 146408 574000 146442 574030
rect 146482 574000 146516 574030
rect 146596 574000 146641 574030
rect 147066 574000 147111 574030
rect 147180 574000 147214 574030
rect 147254 574000 147288 574030
rect 147912 574000 147946 574030
rect 148570 574000 148604 574030
rect 149228 574000 149262 574030
rect 149886 574000 149920 574030
rect 145064 573996 145126 574000
rect 145722 573996 145784 574000
rect 145064 573968 145132 573996
rect 145722 573968 145790 573996
rect 145058 573962 145132 573968
rect 145142 573962 145160 573968
rect 145716 573962 145790 573968
rect 145800 573962 145818 573968
rect 146196 573962 149920 574000
rect 143626 573957 145132 573962
rect 138751 573923 139397 573957
rect 139409 573923 140055 573957
rect 140067 573923 140713 573957
rect 140725 573923 141371 573957
rect 141383 573923 142217 573957
rect 142229 573923 142881 573957
rect 142887 573928 145132 573957
rect 145138 573928 145790 573962
rect 145796 573928 146448 573962
rect 142887 573923 144999 573928
rect 138402 569678 138828 569712
rect 137620 569194 137740 569214
rect 137926 569194 138216 569214
rect 138402 569196 138642 569678
rect 138672 569644 138688 569648
rect 138644 569616 138660 569620
rect 138644 569570 138664 569616
rect 138644 569568 138660 569570
rect 138672 569542 138692 569644
rect 138693 569576 138699 569657
rect 138672 569540 138688 569542
rect 138705 569517 138739 569678
rect 138680 569341 138739 569517
rect 138686 569258 138690 569284
rect 138693 569248 138699 569329
rect 138402 569194 138672 569196
rect 137926 569186 138166 569194
rect 137614 569166 137768 569186
rect 137926 569166 138244 569186
rect 138266 569168 138290 569186
rect 138402 569180 138642 569194
rect 138705 569180 138739 569341
rect 138794 569180 138828 569678
rect 138294 569168 138318 569174
rect 137926 569110 138166 569166
rect 138402 569146 138828 569180
rect 138402 569110 138642 569146
rect 137508 568964 137542 569110
rect 138591 569096 138625 569110
rect 138705 569096 138739 569146
rect 137504 568608 137542 568964
rect 137584 568912 137774 568914
rect 137612 568884 137658 568886
rect 137700 568884 137746 568886
rect 137120 568506 137428 568544
rect 133674 568472 137428 568506
rect 133678 568466 133696 568472
rect 133628 568404 133662 568438
rect 133990 568404 134024 568472
rect 134092 568456 134150 568472
rect 134104 568408 134138 568456
rect 134104 568404 134149 568408
rect 134180 568404 134208 568466
rect 134286 568408 134320 568472
rect 134750 568456 134808 568472
rect 134762 568408 134796 568456
rect 134286 568404 134331 568408
rect 134762 568404 134807 568408
rect 134832 568404 134860 568466
rect 134888 568404 134916 568466
rect 134944 568408 134978 568472
rect 135408 568456 135466 568472
rect 135420 568408 135454 568456
rect 134944 568404 134989 568408
rect 135420 568404 135465 568408
rect 135490 568404 135518 568466
rect 135546 568404 135574 568466
rect 135602 568408 135636 568472
rect 136066 568456 136124 568472
rect 136078 568408 136112 568456
rect 135602 568404 135647 568408
rect 136078 568404 136123 568408
rect 136154 568404 136182 568466
rect 136210 568404 136238 568466
rect 136260 568408 136294 568472
rect 136724 568456 136782 568472
rect 136736 568408 136770 568456
rect 136260 568404 136305 568408
rect 136736 568404 136781 568408
rect 136862 568404 136890 568466
rect 136918 568408 136952 568472
rect 136918 568404 136963 568408
rect 137032 568404 137066 568472
rect 137360 568466 137378 568472
rect 137388 568438 137428 568472
rect 137394 568404 137428 568438
rect 133610 568370 137462 568404
rect 133990 565852 134024 568370
rect 134104 567308 134149 568370
rect 134180 568002 134208 568370
rect 134286 567308 134331 568370
rect 134656 567560 134660 567880
rect 134694 567560 134698 567880
rect 134762 567308 134807 568370
rect 134832 568002 134860 568370
rect 134888 568002 134916 568370
rect 134944 567308 134989 568370
rect 135420 567308 135465 568370
rect 135490 568002 135518 568370
rect 135546 568002 135574 568370
rect 135602 567308 135647 568370
rect 136078 567496 136123 568370
rect 136154 568002 136182 568370
rect 136210 568002 136238 568370
rect 136260 567496 136305 568370
rect 134104 565902 134138 567308
rect 134180 565902 134208 566814
rect 134286 565902 134320 567308
rect 134762 565902 134796 567308
rect 134832 565918 134860 566814
rect 134888 565918 134916 566814
rect 134944 565902 134978 567308
rect 135420 565902 135454 567308
rect 135490 565858 135518 566814
rect 135546 565902 135574 566814
rect 135602 565902 135636 567308
rect 136078 565902 136112 567496
rect 136154 565858 136182 566814
rect 136210 565858 136238 566814
rect 136260 565902 136294 567496
rect 136736 567470 136781 568370
rect 136862 568002 136890 568370
rect 136918 567470 136963 568370
rect 136736 565902 136770 567470
rect 136806 566618 136834 566814
rect 136862 565858 136890 566814
rect 136918 565902 136952 567470
rect 137032 565852 137066 568370
rect 137432 567058 137440 567112
rect 137508 567094 137542 568608
rect 138555 568483 138842 569096
rect 139363 568530 139397 573923
rect 140021 568530 140055 573923
rect 140679 568530 140713 573923
rect 141337 568530 141371 573923
rect 139335 568517 139397 568530
rect 139993 568517 140055 568530
rect 140651 568517 140713 568530
rect 141309 568517 141371 568530
rect 139335 568489 139403 568517
rect 139993 568489 140061 568517
rect 140651 568489 140719 568517
rect 141309 568489 141377 568517
rect 139329 568483 139403 568489
rect 139413 568483 139431 568489
rect 139987 568483 140061 568489
rect 140071 568483 140089 568489
rect 140645 568483 140719 568489
rect 140729 568483 140747 568489
rect 141303 568483 141377 568489
rect 141387 568483 141405 568489
rect 141411 568483 141445 573923
rect 141525 568530 141559 573923
rect 141744 572712 141956 572720
rect 141588 572272 141956 572712
rect 141588 572264 141800 572272
rect 141744 570058 141956 570066
rect 141588 569618 141956 570058
rect 141588 569610 141800 569618
rect 141995 568530 142029 573923
rect 142109 573570 142143 573923
rect 142109 572218 142146 573570
rect 141513 568483 141572 568530
rect 141995 568483 142042 568530
rect 142109 568483 142143 572218
rect 142183 568530 142217 573923
rect 142807 573917 142825 573923
rect 142807 573782 142822 573917
rect 142835 573889 142881 573923
rect 142891 573917 142909 573923
rect 143499 573889 143548 573923
rect 143549 573917 143576 573923
rect 142835 573726 142878 573889
rect 142841 573188 142875 573726
rect 142820 573154 143210 573188
rect 142820 572656 142854 573154
rect 143034 573086 143081 573133
rect 142996 573052 143081 573086
rect 142923 572993 142968 573004
rect 143051 572993 143096 573004
rect 142934 572822 142968 572993
rect 142900 572817 142968 572822
rect 143062 572817 143096 572993
rect 142900 572814 142962 572817
rect 142928 572805 142962 572814
rect 142872 572749 142881 572805
rect 142956 572749 142962 572766
rect 143034 572758 143081 572805
rect 142996 572724 143081 572758
rect 143054 572720 143060 572724
rect 143066 572684 143072 572720
rect 143176 572656 143210 573154
rect 142232 572620 142236 572632
rect 142820 572622 143210 572656
rect 142244 572592 142248 572620
rect 142806 571952 143228 572572
rect 143499 571956 143533 573889
rect 143434 571870 143533 571956
rect 143499 571006 143533 571870
rect 143576 573378 143578 573576
rect 143576 572804 143594 573378
rect 143576 571810 143578 572804
rect 143626 572678 144999 573923
rect 145058 573922 145076 573928
rect 145086 573894 145132 573928
rect 145142 573922 145160 573928
rect 145716 573922 145734 573928
rect 145744 573894 145790 573928
rect 145800 573922 145818 573928
rect 146374 573922 146392 573928
rect 146402 573894 146448 573928
rect 146458 573928 147294 573962
rect 146458 573922 146476 573928
rect 143626 572422 145008 572678
rect 145022 572450 145064 572650
rect 143626 571006 144999 572422
rect 142826 570980 144999 571006
rect 142820 570500 143210 570534
rect 142820 570002 142854 570500
rect 143034 570432 143081 570479
rect 142996 570398 143081 570432
rect 142923 570339 142968 570350
rect 143051 570339 143096 570350
rect 142934 570163 142968 570339
rect 143062 570163 143096 570339
rect 142900 570123 142908 570160
rect 142928 570151 142936 570160
rect 143034 570104 143081 570151
rect 142996 570070 143081 570104
rect 143054 570066 143060 570070
rect 143066 570030 143072 570066
rect 143176 570002 143210 570500
rect 143384 570008 143410 570150
rect 143412 570008 143438 570150
rect 142820 569968 143210 570002
rect 142806 569298 143228 569918
rect 143384 569704 143410 569808
rect 143412 569704 143438 569808
rect 143499 569302 143533 570980
rect 143576 570150 143594 570724
rect 143626 570024 144999 570980
rect 143626 569768 145008 570024
rect 145050 569996 145064 570248
rect 145022 569966 145064 569996
rect 145092 569966 145126 573894
rect 145750 573224 145784 573894
rect 145604 572686 146066 573224
rect 145604 572620 146214 572686
rect 145604 572586 146276 572620
rect 145726 572536 145818 572586
rect 146002 572544 146276 572586
rect 146002 572536 146214 572544
rect 145662 572502 146214 572536
rect 145662 572022 145696 572502
rect 145726 572472 145856 572502
rect 145726 572462 145892 572472
rect 145750 572350 145784 572462
rect 145804 572414 145892 572462
rect 145804 572400 145818 572414
rect 145820 572400 145892 572414
rect 145854 572392 145876 572396
rect 145796 572350 145810 572361
rect 145750 572174 145810 572350
rect 145830 572192 145846 572390
rect 145882 572364 145904 572396
rect 145858 572361 145874 572362
rect 145853 572350 145898 572361
rect 145858 572174 145898 572350
rect 145978 572238 146214 572502
rect 146374 572462 146378 572662
rect 146402 572434 146406 572690
rect 146408 572386 146442 573894
rect 145750 572160 145784 572174
rect 145858 572164 145874 572174
rect 145854 572160 145892 572162
rect 145750 572046 145790 572160
rect 145804 572074 145818 572132
rect 145854 572124 145898 572160
rect 145820 572090 145898 572124
rect 145854 572074 145870 572090
rect 145882 572046 145898 572090
rect 145750 572022 145784 572046
rect 145978 572022 146012 572238
rect 145662 571988 146012 572022
rect 145750 570570 145784 571988
rect 146374 571810 146398 572358
rect 146402 571782 146442 572386
rect 145854 571008 145856 571208
rect 145882 570980 145884 571236
rect 145604 570032 146066 570570
rect 145604 569966 146214 570032
rect 146344 570008 146370 570150
rect 146372 570008 146398 570150
rect 145022 569834 145182 569966
rect 145604 569932 146276 569966
rect 146002 569890 146276 569932
rect 146002 569882 146214 569890
rect 145662 569848 146214 569882
rect 145022 569796 145064 569834
rect 142820 569258 142894 569298
rect 142841 568530 142875 569258
rect 143434 569216 143533 569302
rect 142155 568517 142217 568530
rect 142155 568489 142223 568517
rect 142813 568489 142875 568530
rect 143384 568489 143410 569156
rect 143412 568489 143438 569156
rect 143499 568530 143533 569216
rect 143576 569156 143578 569704
rect 142149 568483 142223 568489
rect 142233 568483 142251 568489
rect 142807 568483 142875 568489
rect 143471 568483 143533 568530
rect 143626 568506 144999 569768
rect 145050 568846 145064 569796
rect 145074 569246 145148 569834
rect 145662 569368 145696 569848
rect 145750 569742 145784 569848
rect 145854 569780 145892 569818
rect 145804 569746 145818 569780
rect 145820 569746 145892 569780
rect 145750 569710 145790 569742
rect 145800 569738 145818 569742
rect 145854 569738 145876 569742
rect 145882 569710 145904 569742
rect 145750 569696 145784 569710
rect 145796 569696 145810 569707
rect 145853 569696 145898 569707
rect 145750 569520 145810 569696
rect 145864 569520 145898 569696
rect 145978 569584 146214 569848
rect 146344 569704 146370 569808
rect 146372 569704 146398 569808
rect 145750 569368 145784 569520
rect 145854 569506 145894 569508
rect 145854 569470 145898 569506
rect 145804 569436 145818 569470
rect 145820 569436 145898 569470
rect 145854 569420 145870 569436
rect 145854 569408 145866 569420
rect 145882 569392 145898 569436
rect 145882 569380 145894 569392
rect 145978 569368 146012 569584
rect 145662 569334 146012 569368
rect 145092 568544 145126 569246
rect 145750 568544 145784 569334
rect 146374 569156 146396 569374
rect 146344 568782 146370 569156
rect 146372 568810 146398 569156
rect 145064 568540 145126 568544
rect 145064 568512 145132 568540
rect 145058 568506 145132 568512
rect 145142 568506 145160 568512
rect 145722 568506 145784 568544
rect 145854 568512 145856 568554
rect 145882 568512 145884 568582
rect 146408 568544 146442 571782
rect 146478 568810 146480 570212
rect 146380 568540 146442 568544
rect 146380 568512 146448 568540
rect 146374 568506 146448 568512
rect 146458 568506 146476 568512
rect 146482 568506 146516 573928
rect 146596 573782 146641 573928
rect 147066 573782 147111 573928
rect 146596 569928 146630 573782
rect 147066 572908 147100 573782
rect 147180 573314 147214 573928
rect 147220 573922 147238 573928
rect 147248 573894 147294 573928
rect 147304 573928 147952 573962
rect 147304 573922 147322 573928
rect 147878 573922 147896 573928
rect 147906 573894 147952 573928
rect 147962 573928 148610 573962
rect 147962 573922 147980 573928
rect 148536 573922 148554 573928
rect 148564 573894 148610 573928
rect 148620 573928 149268 573962
rect 148620 573922 148638 573928
rect 149194 573922 149212 573928
rect 149222 573894 149268 573928
rect 149278 573928 149920 573962
rect 149278 573922 149296 573928
rect 149852 573922 149870 573928
rect 149880 573894 149920 573928
rect 147042 572692 147134 572908
rect 146840 572674 147134 572692
rect 146646 572450 147134 572674
rect 146646 572244 147052 572450
rect 146646 572226 146858 572244
rect 146840 570020 147052 570038
rect 146646 569928 147052 570020
rect 146580 569590 147052 569928
rect 146580 569572 146858 569590
rect 146580 569274 146654 569572
rect 146596 568544 146630 569274
rect 147066 568544 147100 572450
rect 147180 572210 147232 573314
rect 146584 568506 146642 568544
rect 147066 568506 147104 568544
rect 147180 568506 147214 572210
rect 147254 568544 147288 573894
rect 147912 573182 147946 573894
rect 147302 569722 147326 569804
rect 147598 569110 148060 569748
rect 148074 569110 148536 569748
rect 147912 569060 147946 569110
rect 147652 569026 148002 569060
rect 147652 568546 147686 569026
rect 147844 568958 147882 568996
rect 147810 568924 147882 568958
rect 147842 568916 147864 568920
rect 147755 568874 147800 568885
rect 147820 568882 147828 568912
rect 147870 568888 147892 568920
rect 147848 568885 147856 568886
rect 147878 568885 147888 568888
rect 147843 568874 147888 568885
rect 147766 568698 147800 568874
rect 147854 568698 147888 568874
rect 147878 568686 147888 568698
rect 147844 568682 147888 568686
rect 147844 568648 147882 568682
rect 147810 568614 147882 568648
rect 147912 568546 147946 569026
rect 147968 568546 148002 569026
rect 147652 568544 148002 568546
rect 148128 569026 148478 569060
rect 148128 568546 148162 569026
rect 148320 568958 148358 568996
rect 148286 568924 148358 568958
rect 148231 568874 148276 568885
rect 148319 568874 148364 568885
rect 148242 568698 148276 568874
rect 148330 568698 148364 568874
rect 148320 568648 148358 568686
rect 148286 568614 148358 568648
rect 148444 568546 148478 569026
rect 148128 568544 148478 568546
rect 148570 568544 148604 573894
rect 149228 568544 149262 573894
rect 149886 568544 149920 573894
rect 147226 568512 148482 568544
rect 148542 568540 148604 568544
rect 149200 568540 149262 568544
rect 148542 568512 148610 568540
rect 149200 568512 149268 568540
rect 149858 568512 149920 568544
rect 147220 568506 148482 568512
rect 148536 568506 148610 568512
rect 148620 568506 148638 568512
rect 149194 568506 149268 568512
rect 149278 568506 149296 568512
rect 149852 568506 149920 568512
rect 143626 568483 145132 568506
rect 138555 568476 139403 568483
rect 138591 567348 138625 568476
rect 138727 568415 138745 568476
rect 138755 568449 139403 568476
rect 139409 568449 140061 568483
rect 140067 568449 140719 568483
rect 140725 568449 141377 568483
rect 141383 568449 142223 568483
rect 142229 568449 142875 568483
rect 142887 568449 143533 568483
rect 143545 568472 145132 568483
rect 145138 568472 145784 568506
rect 145796 568472 146448 568506
rect 146454 568472 147288 568506
rect 147316 568472 147952 568506
rect 143545 568449 144999 568472
rect 145058 568466 145076 568472
rect 138755 568443 138773 568449
rect 139329 568443 139347 568449
rect 139357 568415 139403 568449
rect 139413 568443 139431 568449
rect 139987 568443 140005 568449
rect 140015 568415 140061 568449
rect 140071 568443 140089 568449
rect 140645 568443 140663 568449
rect 138705 568381 138739 568415
rect 139363 568381 139397 568415
rect 140021 568381 140055 568415
rect 140142 568381 140164 568438
rect 140673 568415 140719 568449
rect 140729 568443 140747 568449
rect 141303 568443 141321 568449
rect 141331 568415 141377 568449
rect 141387 568443 141405 568449
rect 140679 568381 140713 568415
rect 141337 568381 141371 568415
rect 141411 568381 141445 568449
rect 141513 568433 141571 568449
rect 141525 568381 141559 568433
rect 141995 568381 142029 568449
rect 142109 568381 142143 568449
rect 142149 568443 142167 568449
rect 142177 568415 142223 568449
rect 142233 568443 142251 568449
rect 142807 568443 142825 568449
rect 142835 568415 142875 568449
rect 142183 568381 142217 568415
rect 142841 568381 142875 568415
rect 143384 568381 143410 568443
rect 143412 568381 143438 568443
rect 143499 568381 143533 568449
rect 143626 568404 144999 568449
rect 145086 568438 145132 568472
rect 145142 568466 145160 568472
rect 145092 568404 145126 568438
rect 145750 568404 145784 568472
rect 146374 568466 146392 568472
rect 145854 568404 145856 568466
rect 145882 568404 145884 568466
rect 146402 568438 146448 568472
rect 146458 568466 146476 568472
rect 146408 568404 146442 568438
rect 146482 568404 146516 568472
rect 146584 568456 146642 568472
rect 146596 568408 146630 568456
rect 147066 568408 147100 568472
rect 146596 568404 146641 568408
rect 147066 568404 147111 568408
rect 147180 568404 147214 568472
rect 147220 568466 147238 568472
rect 147248 568438 147288 568472
rect 147254 568404 147288 568438
rect 147324 568404 147326 568472
rect 147874 568404 147886 568472
rect 147912 568438 147952 568472
rect 147962 568472 148610 568506
rect 148616 568472 149268 568506
rect 149274 568472 149920 568506
rect 147962 568466 147980 568472
rect 148536 568466 148554 568472
rect 148564 568438 148610 568472
rect 148620 568466 148638 568472
rect 149194 568466 149212 568472
rect 149222 568438 149268 568472
rect 149278 568466 149296 568472
rect 149852 568466 149870 568472
rect 149880 568438 149920 568472
rect 147912 568404 147946 568438
rect 148570 568404 148604 568438
rect 149228 568404 149262 568438
rect 149354 568404 149360 568438
rect 149886 568404 149920 568438
rect 143626 568381 149954 568404
rect 138687 568370 149954 568381
rect 138687 568347 144999 568370
rect 145854 568354 145856 568370
rect 138555 567094 138642 567348
rect 137450 566456 137578 567094
rect 137588 566675 137596 566875
rect 137926 566560 138166 567094
rect 138402 567058 138642 567094
rect 138705 567058 138766 567092
rect 138402 567024 138828 567058
rect 137620 566540 137740 566560
rect 137926 566540 138216 566560
rect 138402 566542 138642 567024
rect 138693 566922 138699 567003
rect 138705 566863 138739 567024
rect 138680 566687 138739 566863
rect 138686 566604 138690 566630
rect 138693 566594 138699 566675
rect 138705 566560 138739 566687
rect 138402 566540 138672 566542
rect 137926 566532 138166 566540
rect 137614 566512 137768 566532
rect 137926 566512 138244 566532
rect 138266 566514 138290 566532
rect 138402 566526 138642 566540
rect 138705 566526 138766 566560
rect 138794 566526 138828 567024
rect 138294 566514 138318 566520
rect 137926 566456 138166 566512
rect 138402 566492 138828 566526
rect 138402 566456 138642 566492
rect 137508 566310 137542 566456
rect 138591 566442 138625 566456
rect 137504 565954 137542 566310
rect 137584 566258 137774 566260
rect 137612 566230 137658 566232
rect 137700 566230 137746 566232
rect 133990 565818 137366 565852
rect 133990 565802 134024 565818
rect 135490 565806 135518 565812
rect 133990 565791 134001 565802
rect 134013 565791 134024 565802
rect 136154 565800 136182 565812
rect 136210 565806 136238 565812
rect 136862 565800 136890 565812
rect 137032 565802 137066 565818
rect 137508 565812 137542 565954
rect 138555 565822 138842 566442
rect 140021 565888 140055 568347
rect 140142 568004 140164 568347
rect 140306 568158 140696 568192
rect 140306 567660 140340 568158
rect 140520 568090 140567 568137
rect 140482 568056 140567 568090
rect 140662 568130 140696 568158
rect 140409 567997 140454 568008
rect 140537 567997 140582 568008
rect 140420 567821 140454 567997
rect 140548 567821 140582 567997
rect 140520 567762 140567 567809
rect 140482 567728 140567 567762
rect 140662 567722 140730 568130
rect 140662 567660 140696 567722
rect 140306 567626 140696 567660
rect 140288 567066 140710 567576
rect 140288 566956 140712 567066
rect 140645 566814 140678 566956
rect 140679 566780 140712 566956
rect 141411 565829 141445 568347
rect 141525 565888 141559 568347
rect 141995 565888 142029 568347
rect 142109 565829 142143 568347
rect 143384 568002 143410 568347
rect 143412 568002 143438 568347
rect 142820 566928 142894 567258
rect 142744 566698 142748 566814
rect 142820 566774 143026 566928
rect 142820 566604 142894 566774
rect 143384 565835 143410 566814
rect 143412 566754 143466 566814
rect 143412 565835 143438 566754
rect 143499 565888 143533 568347
rect 137032 565791 137043 565802
rect 137055 565791 137066 565802
rect 131961 565768 131972 565779
rect 131984 565768 131995 565779
rect 128539 565693 132375 565727
rect 133610 565716 137446 565750
rect 140016 565727 140986 565828
rect 141411 565795 142143 565829
rect 141411 565779 141445 565795
rect 141411 565768 141422 565779
rect 141434 565768 141445 565779
rect 142109 565779 142143 565795
rect 143384 565782 143410 565789
rect 142109 565768 142120 565779
rect 142132 565768 142143 565779
rect 143412 565754 143438 565789
rect 143626 565750 144999 568347
rect 145882 568326 145884 568370
rect 145050 566192 145064 566814
rect 145854 566754 145866 566814
rect 145882 566698 145922 566814
rect 146344 566128 146370 566814
rect 146372 566156 146398 566814
rect 146478 566156 146480 566814
rect 146482 565852 146516 568370
rect 146596 567308 146641 568370
rect 147066 567308 147111 568370
rect 146596 565902 146630 567308
rect 147066 565902 147100 567308
rect 147180 565852 147214 568370
rect 147254 565920 147288 568370
rect 147912 568356 147924 568370
rect 149228 568284 149262 568370
rect 149170 568202 149262 568284
rect 147302 567068 147326 567150
rect 147598 566456 148060 567094
rect 148074 566456 148536 567094
rect 148702 566628 148714 566814
rect 147912 566406 147940 566440
rect 147652 566372 148002 566406
rect 147254 565902 147302 565920
rect 147288 565898 147302 565902
rect 147652 565892 147686 566372
rect 147844 566304 147882 566342
rect 147810 566270 147882 566304
rect 147842 566262 147864 566266
rect 147755 566220 147800 566231
rect 147820 566228 147828 566258
rect 147870 566234 147892 566266
rect 147912 566258 147922 566270
rect 147848 566231 147856 566232
rect 147878 566231 147888 566234
rect 147843 566220 147888 566231
rect 147766 566044 147800 566220
rect 147854 566044 147888 566220
rect 147878 566032 147888 566044
rect 147844 566028 147888 566032
rect 147844 565994 147882 566028
rect 147912 566006 147926 566258
rect 147912 565994 147922 566006
rect 147810 565960 147882 565994
rect 147934 565926 147946 566372
rect 147912 565902 147946 565926
rect 147934 565898 147946 565902
rect 147968 565892 148002 566372
rect 147250 565858 147266 565886
rect 146482 565818 147214 565852
rect 147222 565852 147238 565858
rect 147222 565830 147242 565852
rect 147234 565818 147242 565830
rect 146482 565802 146516 565818
rect 146482 565791 146493 565802
rect 146505 565791 146516 565802
rect 147180 565802 147214 565818
rect 147180 565791 147191 565802
rect 147203 565791 147214 565802
rect 147268 565784 147276 565886
rect 147652 565858 148002 565892
rect 148128 566372 148478 566406
rect 148128 565892 148162 566372
rect 148320 566304 148358 566342
rect 148286 566270 148358 566304
rect 148231 566220 148276 566231
rect 148319 566220 148364 566231
rect 148242 566044 148276 566220
rect 148330 566044 148364 566220
rect 148320 565994 148358 566032
rect 148286 565960 148358 565994
rect 148444 565892 148478 566372
rect 149228 565902 149262 568202
rect 149354 568004 149360 568370
rect 149466 567590 149928 568228
rect 149952 567774 149954 567818
rect 149520 567506 149870 567540
rect 149520 567026 149554 567506
rect 149712 567472 149750 567476
rect 149704 567470 149762 567472
rect 149712 567438 149750 567470
rect 149678 567404 149750 567438
rect 149623 567354 149668 567365
rect 149711 567354 149756 567365
rect 149634 567178 149668 567354
rect 149722 567178 149756 567354
rect 149712 567128 149750 567166
rect 149678 567094 149750 567128
rect 149836 567032 149870 567506
rect 149886 567066 149904 567470
rect 149924 567456 149926 567564
rect 149952 567456 149954 567564
rect 149836 567026 149874 567032
rect 149520 566992 149874 567026
rect 149852 566814 149874 566992
rect 149886 566780 149908 567066
rect 148128 565858 148478 565892
rect 147316 565826 147884 565852
rect 147316 565818 147886 565826
rect 147934 565784 147950 565858
rect 147962 565812 147978 565858
rect 150000 565812 150034 575324
rect 150571 575288 154195 575324
rect 150607 569712 150641 575288
rect 153353 574059 153387 575288
rect 150709 574025 154057 574059
rect 150721 574004 150755 574025
rect 151379 574004 151413 574025
rect 152037 574004 152071 574025
rect 152695 574004 152729 574025
rect 153353 574004 153387 574025
rect 154011 574004 154045 574025
rect 150721 573957 154045 574004
rect 150721 573889 150761 573957
rect 150771 573923 151419 573957
rect 150771 573917 150789 573923
rect 151345 573917 151363 573923
rect 151373 573889 151419 573923
rect 151429 573923 152077 573957
rect 151429 573917 151447 573923
rect 152003 573917 152021 573923
rect 152031 573889 152077 573923
rect 152087 573923 152735 573957
rect 152087 573917 152105 573923
rect 152661 573917 152679 573923
rect 152689 573889 152735 573923
rect 152745 573923 153393 573957
rect 152745 573917 152763 573923
rect 153319 573917 153337 573923
rect 153347 573889 153393 573923
rect 153403 573923 154045 573957
rect 153403 573917 153421 573923
rect 153977 573917 153995 573923
rect 154005 573889 154045 573923
rect 150683 569722 150684 569804
rect 150721 569712 150755 573889
rect 150550 569678 150844 569712
rect 150607 569610 150641 569678
rect 150614 569567 150641 569610
rect 150709 569576 150715 569657
rect 150573 569325 150602 569533
rect 150607 569291 150641 569567
rect 150721 569517 150755 569678
rect 150696 569341 150755 569517
rect 150614 569248 150641 569291
rect 150702 569258 150706 569284
rect 150709 569248 150715 569329
rect 150607 569214 150641 569248
rect 150588 569194 150688 569214
rect 150607 569186 150641 569194
rect 150582 569180 150688 569186
rect 150721 569180 150755 569341
rect 150810 569180 150844 569678
rect 150550 569146 150844 569180
rect 150930 569678 151320 569712
rect 150930 569180 150964 569678
rect 151144 569610 151191 569657
rect 151106 569576 151191 569610
rect 151033 569517 151078 569528
rect 151161 569517 151206 569528
rect 151044 569341 151078 569517
rect 151172 569341 151206 569517
rect 151144 569282 151191 569329
rect 151106 569248 151191 569282
rect 151286 569180 151320 569678
rect 150930 569146 151320 569180
rect 150602 569134 150641 569146
rect 150607 569096 150641 569134
rect 150721 569096 150755 569146
rect 150571 568530 150858 569096
rect 150912 568530 151334 569096
rect 151379 568530 151413 573889
rect 151468 569168 151478 569518
rect 151496 569168 151506 569546
rect 151468 568694 151478 568982
rect 151496 568666 151506 568982
rect 152037 568530 152071 573889
rect 152695 568530 152729 573889
rect 153353 568530 153387 573889
rect 154011 568530 154045 573889
rect 150571 568483 151334 568530
rect 151351 568517 151413 568530
rect 152009 568517 152071 568530
rect 152667 568517 152729 568530
rect 153325 568517 153387 568530
rect 151351 568489 151419 568517
rect 152009 568489 152077 568517
rect 152667 568489 152735 568517
rect 153325 568489 153393 568517
rect 153983 568489 154045 568530
rect 151345 568483 151419 568489
rect 151429 568483 151447 568489
rect 152003 568483 152077 568489
rect 152087 568483 152105 568489
rect 152661 568483 152735 568489
rect 152745 568483 152763 568489
rect 153319 568483 153393 568489
rect 153403 568483 153421 568489
rect 153977 568483 154045 568489
rect 150571 568476 151419 568483
rect 150042 567174 150050 567276
rect 150070 567150 150078 567248
rect 150607 567058 150641 568476
rect 150683 568394 150706 568476
rect 150721 568415 150770 568476
rect 150771 568449 151419 568476
rect 151425 568449 152077 568483
rect 152083 568449 152735 568483
rect 152741 568449 153393 568483
rect 153399 568449 154045 568483
rect 150771 568443 150798 568449
rect 151345 568443 151363 568449
rect 151373 568415 151419 568449
rect 151429 568443 151447 568449
rect 152003 568443 152021 568449
rect 152031 568415 152077 568449
rect 152087 568443 152105 568449
rect 152661 568443 152679 568449
rect 152689 568415 152735 568449
rect 152745 568443 152763 568449
rect 153319 568443 153337 568449
rect 153347 568415 153393 568449
rect 153403 568443 153421 568449
rect 153977 568443 153995 568449
rect 154005 568415 154045 568449
rect 150721 568381 150755 568415
rect 151379 568381 151413 568415
rect 152037 568381 152071 568415
rect 152695 568381 152729 568415
rect 153353 568381 153387 568415
rect 154011 568381 154045 568415
rect 150703 568347 154057 568381
rect 154063 568347 154079 568381
rect 150683 567068 150684 567150
rect 150721 567092 150722 567188
rect 150721 567058 150782 567092
rect 150550 567024 150844 567058
rect 150607 566956 150641 567024
rect 150614 566913 150641 566956
rect 150709 566922 150715 567003
rect 150573 566671 150602 566879
rect 150607 566637 150641 566913
rect 150721 566863 150755 567024
rect 150696 566687 150755 566863
rect 150614 566636 150641 566637
rect 150588 566618 150688 566636
rect 150614 566594 150641 566618
rect 150702 566604 150706 566630
rect 150709 566594 150715 566675
rect 150607 566560 150641 566594
rect 150721 566560 150755 566687
rect 150588 566540 150688 566560
rect 150607 566532 150641 566540
rect 150582 566526 150688 566532
rect 150721 566526 150782 566560
rect 150810 566526 150844 567024
rect 150550 566492 150844 566526
rect 150930 567024 151320 567058
rect 150930 566526 150964 567024
rect 151144 566956 151191 567003
rect 151106 566922 151191 566956
rect 151033 566863 151078 566874
rect 151161 566863 151206 566874
rect 151044 566687 151078 566863
rect 151172 566687 151206 566863
rect 151144 566628 151191 566675
rect 151106 566594 151191 566628
rect 151286 566526 151320 567024
rect 150930 566492 151320 566526
rect 151468 566514 151478 566814
rect 151496 566628 151534 566814
rect 151496 566514 151506 566628
rect 150602 566480 150641 566492
rect 150607 566442 150641 566480
rect 150571 565822 150858 566442
rect 150912 565822 151334 566442
rect 151468 566040 151478 566328
rect 151496 566012 151506 566328
rect 150743 565761 150770 565822
rect 150771 565789 150798 565822
rect 154125 565789 154159 575288
rect 155678 565812 155712 575324
rect 157842 574846 157862 575042
rect 158424 574064 158458 575324
rect 155780 574030 159128 574064
rect 155792 574000 155826 574030
rect 156450 574000 156484 574030
rect 157108 574000 157142 574030
rect 157766 574000 157800 574030
rect 158424 574000 158458 574030
rect 159082 574000 159116 574030
rect 155792 573962 159116 574000
rect 155792 568540 155826 573962
rect 155854 573928 156490 573962
rect 156416 573922 156434 573928
rect 156444 573894 156490 573928
rect 156500 573928 157148 573962
rect 156500 573922 156518 573928
rect 157074 573922 157092 573928
rect 157102 573894 157148 573928
rect 157158 573928 157806 573962
rect 157158 573922 157176 573928
rect 157732 573922 157750 573928
rect 157760 573894 157806 573928
rect 157816 573928 158464 573962
rect 157816 573922 157834 573928
rect 158390 573922 158408 573928
rect 158418 573894 158464 573928
rect 158474 573928 159116 573962
rect 158474 573922 158492 573928
rect 159048 573922 159066 573928
rect 159076 573894 159116 573928
rect 155858 569706 155864 569962
rect 155886 569734 155892 569934
rect 155858 569306 155864 569562
rect 155886 569334 155892 569534
rect 156450 568544 156484 573894
rect 157108 568544 157142 573894
rect 157766 568544 157800 573894
rect 158424 568544 158458 573894
rect 159082 568544 159116 573894
rect 156422 568540 156484 568544
rect 157080 568540 157142 568544
rect 157738 568540 157800 568544
rect 158396 568540 158458 568544
rect 155792 568438 155832 568540
rect 156422 568512 156490 568540
rect 157080 568512 157148 568540
rect 157738 568512 157806 568540
rect 158396 568512 158464 568540
rect 159054 568512 159116 568544
rect 155842 568506 155860 568512
rect 156416 568506 156490 568512
rect 156500 568506 156518 568512
rect 157074 568506 157148 568512
rect 157158 568506 157176 568512
rect 157732 568506 157806 568512
rect 157816 568506 157834 568512
rect 158390 568506 158464 568512
rect 158474 568506 158492 568512
rect 159048 568506 159116 568512
rect 155838 568472 156490 568506
rect 156496 568472 157148 568506
rect 157154 568472 157806 568506
rect 157812 568472 158464 568506
rect 158470 568472 159116 568506
rect 155842 568466 155860 568472
rect 156416 568466 156434 568472
rect 156444 568438 156490 568472
rect 156500 568466 156518 568472
rect 157074 568466 157092 568472
rect 157102 568438 157148 568472
rect 157158 568466 157176 568472
rect 157732 568466 157750 568472
rect 157760 568438 157806 568472
rect 157816 568466 157834 568472
rect 158390 568466 158408 568472
rect 158418 568438 158464 568472
rect 158474 568466 158492 568472
rect 159048 568466 159066 568472
rect 159076 568438 159116 568472
rect 155792 568404 155826 568438
rect 156450 568404 156484 568438
rect 157108 568404 157142 568438
rect 157766 568404 157800 568438
rect 158424 568404 158458 568438
rect 159082 568404 159116 568438
rect 155774 568370 159150 568404
rect 156450 565902 156484 568370
rect 159196 565812 159230 575324
rect 164861 575288 168485 575324
rect 173005 575302 173556 575338
rect 173748 575349 175230 575417
rect 175521 575349 175555 575417
rect 175787 575349 175832 575417
rect 176078 575401 176136 575417
rect 176090 575349 176124 575401
rect 176204 575349 176238 575417
rect 176433 575411 176491 575417
rect 176346 575388 176382 575411
rect 176402 575401 176491 575411
rect 176346 575349 176362 575388
rect 176402 575349 176438 575401
rect 176476 575386 176491 575401
rect 176445 575349 176479 575383
rect 176559 575349 176593 575417
rect 177016 575404 177044 575411
rect 177072 575404 177100 575411
rect 177478 575390 179109 575417
rect 179542 575406 179580 575428
rect 179530 575390 179588 575406
rect 180116 575390 180150 575458
rect 180292 575440 183968 575458
rect 184030 575444 184492 576064
rect 184546 575444 184968 576064
rect 185022 575451 185444 576064
rect 185965 575942 185999 576142
rect 185931 575498 185954 575942
rect 185959 575498 186005 575942
rect 186238 575498 186272 576469
rect 185931 575470 185984 575498
rect 185937 575451 185984 575470
rect 186226 575451 186284 575498
rect 185022 575444 185984 575451
rect 180296 575434 180332 575440
rect 180200 575406 180238 575428
rect 180592 575406 180626 575440
rect 180780 575434 180984 575440
rect 181432 575434 181468 575440
rect 180780 575428 180810 575434
rect 180838 575428 180984 575434
rect 180846 575424 180904 575428
rect 181504 575424 182716 575440
rect 182800 575434 182834 575440
rect 180858 575406 180896 575424
rect 181516 575406 181562 575424
rect 181630 575406 181664 575424
rect 182336 575416 182698 575424
rect 182756 575422 182784 575434
rect 182800 575428 182840 575434
rect 182800 575424 182834 575428
rect 182800 575413 182811 575424
rect 182823 575413 182834 575424
rect 183464 575422 183492 575434
rect 183634 575424 183668 575440
rect 183634 575413 183645 575424
rect 183657 575413 183668 575424
rect 180188 575396 182658 575406
rect 180188 575390 182670 575396
rect 177478 575372 181562 575390
rect 181630 575372 181664 575390
rect 182092 575388 182670 575390
rect 182092 575372 182336 575388
rect 182800 575372 182834 575396
rect 184030 575372 184198 575444
rect 177478 575356 184198 575372
rect 177478 575349 179109 575356
rect 173748 575315 179109 575349
rect 179530 575318 179588 575356
rect 180116 575338 184198 575356
rect 185193 575349 185227 575444
rect 185369 575417 185984 575444
rect 186027 575417 186284 575451
rect 186226 575401 186284 575417
rect 186269 575386 186284 575401
rect 186238 575349 186272 575383
rect 186352 575349 186386 576630
rect 187927 575528 187985 575546
rect 188013 575528 188047 583545
rect 188116 583486 188172 583497
rect 188586 583486 188642 583497
rect 188127 579998 188172 583486
rect 188597 579998 188642 583486
rect 188711 583192 188745 583545
rect 190123 583511 190150 583613
rect 190151 583539 190178 583585
rect 188711 581840 188748 583192
rect 188127 577604 188161 579998
rect 188346 579680 188558 579688
rect 188190 579240 188558 579680
rect 188190 579232 188402 579240
rect 188597 577604 188631 579998
rect 188127 576600 188172 577604
rect 188597 576600 188642 577604
rect 188127 575528 188161 576600
rect 188597 575528 188631 576600
rect 188711 575528 188745 581840
rect 188785 575546 188819 583486
rect 190178 582414 190180 583198
rect 190228 582414 191601 583647
rect 191664 583615 191702 583622
rect 191652 583550 191702 583615
rect 192122 583615 192160 583622
rect 192122 583600 192168 583615
rect 192110 583584 192168 583600
rect 191756 583550 192168 583584
rect 191652 583512 191698 583550
rect 192110 583512 192168 583550
rect 188920 582380 191601 582414
rect 188846 581840 188870 582038
rect 188846 581114 188852 581362
rect 188920 580128 188954 582380
rect 189443 582300 189477 582380
rect 190101 582300 190135 582380
rect 190178 582306 190180 582380
rect 190228 582300 191601 582380
rect 188975 582238 189056 582285
rect 189115 582266 191601 582300
rect 189430 582254 189431 582255
rect 189431 582253 189432 582254
rect 189022 580270 189056 582238
rect 189443 580346 189477 582266
rect 189489 582254 189490 582255
rect 190088 582254 190089 582255
rect 189488 582253 189489 582254
rect 190089 582253 190090 582254
rect 190101 580346 190135 582266
rect 190147 582254 190148 582255
rect 190146 582253 190147 582254
rect 190178 581982 190180 582260
rect 189443 580255 189488 580346
rect 190101 580255 190146 580346
rect 189431 580254 189432 580255
rect 189443 580254 189489 580255
rect 190089 580254 190090 580255
rect 190101 580254 190147 580255
rect 189430 580253 189431 580254
rect 189424 580242 189431 580253
rect 189443 580242 189477 580254
rect 189489 580253 189490 580254
rect 190088 580253 190089 580254
rect 189489 580242 190089 580253
rect 190101 580242 190135 580254
rect 190147 580253 190148 580254
rect 190178 580253 190196 580346
rect 190147 580242 190196 580253
rect 190228 580242 191601 582266
rect 191658 583500 191698 583512
rect 191710 583500 191728 583511
rect 191658 580920 191728 583500
rect 191642 580852 191728 580920
rect 191642 580646 191739 580852
rect 192122 580800 192156 583512
rect 192236 582652 192270 583652
rect 193084 583584 193118 583631
rect 193782 583600 193793 583611
rect 193805 583600 193816 583611
rect 193782 583584 193816 583600
rect 193084 583550 193816 583584
rect 192236 582542 192404 582652
rect 192236 582516 192420 582542
rect 192236 580800 192270 582516
rect 192328 582084 192420 582516
rect 193084 582508 193118 583550
rect 193187 583500 193232 583511
rect 193657 583500 193702 583511
rect 193198 582952 193232 583500
rect 193668 582952 193702 583500
rect 193198 582508 193243 582952
rect 193668 582530 193713 582952
rect 193782 582936 193816 583550
rect 194344 583236 194378 583652
rect 194486 583628 194552 583648
rect 194472 583618 194552 583628
rect 194472 583610 194578 583618
rect 194472 583606 194556 583610
rect 194472 583600 194486 583606
rect 194518 583600 194552 583606
rect 194560 583598 194594 583600
rect 194424 583590 194486 583598
rect 194424 583584 194498 583590
rect 194444 583582 194502 583584
rect 194452 583580 194502 583582
rect 194452 583578 194498 583580
rect 194464 583576 194492 583578
rect 194504 583576 194534 583598
rect 194560 583584 194614 583598
rect 194546 583582 194606 583584
rect 194546 583576 194576 583582
rect 194446 583564 194524 583576
rect 194545 583564 194592 583576
rect 194446 583550 194520 583564
rect 194446 583512 194502 583550
rect 194514 583512 194526 583516
rect 194546 583512 194592 583564
rect 194458 583388 194498 583512
rect 194424 583348 194430 583378
rect 194452 583376 194458 583378
rect 194480 583376 194498 583388
rect 194504 583500 194534 583512
rect 194546 583500 194580 583512
rect 194504 583388 194580 583500
rect 194504 583376 194548 583388
rect 194480 583372 194492 583376
rect 194504 583372 194552 583376
rect 194504 583354 194570 583372
rect 194502 583304 194570 583354
rect 194502 583288 194552 583304
rect 194660 583236 194694 583652
rect 195824 583500 195870 583512
rect 195830 583488 195870 583500
rect 194344 583202 194694 583236
rect 193644 582508 193736 582530
rect 193782 582508 193834 582936
rect 192848 581570 195814 582508
rect 196360 582476 196672 582512
rect 197209 582476 197243 583585
rect 197448 583250 200797 583717
rect 202428 583686 204078 584664
rect 204514 583686 205868 584664
rect 208708 584526 208726 584748
rect 208736 584725 208800 584748
rect 208742 584722 208800 584725
rect 210026 584725 210098 584746
rect 210026 584722 210092 584725
rect 210026 584550 210048 584722
rect 202280 583652 205868 583686
rect 202280 583326 202314 583652
rect 202428 583584 204078 583652
rect 204340 583584 204378 583622
rect 204514 583584 205868 583652
rect 202428 583550 204378 583584
rect 204430 583550 205868 583584
rect 202428 583518 204078 583550
rect 204514 583516 205868 583550
rect 205657 583512 205658 583513
rect 205730 583512 205752 583516
rect 205658 583511 205659 583512
rect 202383 583500 202428 583511
rect 203041 583500 203086 583511
rect 203699 583500 203744 583511
rect 204357 583500 204402 583511
rect 205015 583500 205060 583511
rect 202394 583326 202428 583500
rect 202439 583338 202440 583339
rect 203040 583338 203041 583339
rect 202440 583337 202441 583338
rect 203039 583337 203040 583338
rect 203052 583326 203086 583500
rect 203097 583338 203098 583339
rect 203698 583338 203699 583339
rect 203098 583337 203099 583338
rect 203697 583337 203698 583338
rect 203710 583326 203744 583500
rect 203755 583338 203756 583339
rect 204356 583338 204357 583339
rect 203756 583337 203757 583338
rect 204355 583337 204356 583338
rect 204368 583326 204402 583500
rect 204413 583338 204414 583339
rect 205014 583338 205015 583339
rect 204414 583337 204415 583338
rect 205013 583337 205014 583338
rect 205026 583326 205060 583500
rect 205672 583354 205752 583512
rect 205071 583338 205072 583339
rect 205672 583338 205730 583354
rect 205072 583337 205073 583338
rect 205646 583332 205657 583337
rect 205646 583326 205658 583332
rect 202246 583298 205662 583326
rect 205678 583302 205696 583338
rect 205715 583323 205730 583338
rect 205678 583298 205730 583302
rect 202246 583292 205730 583298
rect 202280 583250 202314 583292
rect 202394 583250 202428 583292
rect 202440 583280 202441 583281
rect 203039 583280 203040 583281
rect 202439 583279 202440 583280
rect 203040 583279 203041 583280
rect 197448 582679 202780 583250
rect 203052 582952 203086 583292
rect 203098 583280 203099 583281
rect 203697 583280 203698 583281
rect 203097 583279 203098 583280
rect 203698 583279 203699 583280
rect 203710 582952 203744 583292
rect 203756 583280 203757 583281
rect 204355 583280 204356 583281
rect 203755 583279 203756 583280
rect 204356 583279 204357 583280
rect 202974 582746 203008 582752
rect 203008 582696 203030 582746
rect 203052 582681 203097 582952
rect 203144 582746 203226 582752
rect 203040 582680 203041 582681
rect 203052 582680 203098 582681
rect 203039 582679 203040 582680
rect 197448 582678 203040 582679
rect 203052 582678 203086 582680
rect 203098 582679 203099 582680
rect 203150 582679 203170 582696
rect 203178 582679 203226 582746
rect 203710 582681 203755 582952
rect 203698 582680 203699 582681
rect 203710 582680 203756 582681
rect 204356 582680 204357 582681
rect 203697 582679 203698 582680
rect 203098 582678 203698 582679
rect 197448 582668 203698 582678
rect 203710 582668 203744 582680
rect 203756 582679 203757 582680
rect 204355 582679 204356 582680
rect 203756 582668 204334 582679
rect 204368 582668 204402 583292
rect 204414 583280 204415 583281
rect 205013 583280 205014 583281
rect 204413 583279 204414 583280
rect 205014 583279 205015 583280
rect 204413 582680 204414 582681
rect 205014 582680 205015 582681
rect 204414 582679 204415 582680
rect 205013 582679 205014 582680
rect 205026 582668 205060 583292
rect 205650 583286 205658 583292
rect 205072 583280 205073 583281
rect 205071 583279 205072 583280
rect 205662 583264 205730 583292
rect 205672 582696 205752 583264
rect 205071 582680 205072 582681
rect 205672 582680 205730 582696
rect 205072 582679 205073 582680
rect 205646 582668 205657 582679
rect 197448 582640 205662 582668
rect 205684 582644 205696 582680
rect 205715 582665 205730 582680
rect 205680 582640 205730 582644
rect 197448 582634 205730 582640
rect 197448 582512 202780 582634
rect 202982 582628 203150 582634
rect 202982 582542 203170 582628
rect 203178 582542 203226 582628
rect 203697 582622 203698 582623
rect 203710 582622 203744 582634
rect 203756 582622 203757 582623
rect 204355 582622 204356 582623
rect 203698 582621 203699 582622
rect 203710 582621 203756 582622
rect 204356 582621 204357 582622
rect 202982 582512 203150 582542
rect 203710 582512 203755 582621
rect 197323 582476 197357 582510
rect 197448 582476 204174 582512
rect 196360 582442 204174 582476
rect 193084 580800 193118 581570
rect 193198 580800 193232 581570
rect 193668 580800 193702 581570
rect 193782 580800 193816 581570
rect 195838 580806 195870 582244
rect 195894 580806 195898 582188
rect 196360 581144 196672 582442
rect 197209 582374 197243 582442
rect 197448 582421 204174 582442
rect 197112 581992 197122 582316
rect 197209 582315 197210 582347
rect 197214 582315 197243 582374
rect 197162 582288 197208 582293
rect 197209 582288 197243 582315
rect 197311 582340 204174 582421
rect 197311 582293 197369 582340
rect 197140 582281 197243 582288
rect 197140 582278 197202 582281
rect 197140 582020 197178 582278
rect 197162 581848 197178 582020
rect 197204 582020 197243 582281
rect 197162 581305 197202 581848
rect 197204 581305 197208 582020
rect 197162 581293 197208 581305
rect 197175 581289 197202 581293
rect 197209 581255 197243 582020
rect 197323 581848 197368 582293
rect 197448 582010 204174 582340
rect 204284 582094 204328 582114
rect 204328 582058 204340 582094
rect 204356 582022 204357 582023
rect 204355 582021 204356 582022
rect 204368 582010 204402 582634
rect 204414 582622 204415 582623
rect 205013 582622 205014 582623
rect 204413 582621 204414 582622
rect 205014 582621 205015 582622
rect 204413 582022 204414 582023
rect 205014 582022 205015 582023
rect 204414 582021 204415 582022
rect 205013 582021 205014 582022
rect 205026 582010 205060 582634
rect 205072 582622 205073 582623
rect 205071 582621 205072 582622
rect 205662 582606 205730 582634
rect 205672 582038 205752 582606
rect 205071 582022 205072 582023
rect 205672 582022 205730 582038
rect 205072 582021 205073 582022
rect 205646 582010 205657 582021
rect 197448 581976 205662 582010
rect 197448 581896 204174 581976
rect 204328 581896 204340 581922
rect 204368 581896 204402 581976
rect 205026 581896 205060 581976
rect 205684 581942 205696 582022
rect 205715 582007 205730 582022
rect 197448 581862 205730 581896
rect 197323 581293 197357 581848
rect 197448 581826 204174 581862
rect 197826 581788 197871 581826
rect 197826 581460 197860 581788
rect 197940 581658 197974 581826
rect 197981 581658 198021 581826
rect 198026 581812 198094 581826
rect 198026 581658 198077 581812
rect 198482 581658 198516 581826
rect 198596 581658 198630 581826
rect 198639 581658 198673 581826
rect 198794 581808 199016 581826
rect 199192 581790 199208 581826
rect 199254 581658 199288 581826
rect 199297 581658 199337 581826
rect 199348 581658 199365 581826
rect 199906 581790 199946 581826
rect 199912 581658 199946 581790
rect 199955 581658 199984 581826
rect 200026 581658 200060 581826
rect 200586 581666 200654 581826
rect 200688 581666 200713 581826
rect 200727 581666 200761 581826
rect 202244 581674 204174 581826
rect 204328 581814 204340 581862
rect 197918 581460 198910 581658
rect 197590 581293 198910 581460
rect 197214 581246 197243 581255
rect 197311 581246 197370 581293
rect 197448 581291 198910 581293
rect 197448 581246 199016 581291
rect 197214 581244 199016 581246
rect 199108 581244 200100 581658
rect 197214 581212 200100 581244
rect 197209 581144 197243 581212
rect 197311 581196 197369 581212
rect 197590 581210 200100 581212
rect 197311 581181 197326 581196
rect 197323 581144 197357 581178
rect 197590 581144 198924 581210
rect 196360 581142 198924 581144
rect 198946 581142 198984 581202
rect 199038 581154 199062 581200
rect 199052 581142 199062 581154
rect 199108 581142 200100 581210
rect 196360 581110 200100 581142
rect 196360 581074 196672 581110
rect 191664 580628 191739 580646
rect 191638 580400 191784 580628
rect 191664 580390 191739 580400
rect 191604 580360 191610 580390
rect 191632 580388 191739 580390
rect 191766 580388 191790 580390
rect 191642 580330 191739 580388
rect 191794 580360 191818 580390
rect 189115 580208 191601 580242
rect 191630 580216 191636 580258
rect 191658 580256 191739 580330
rect 191658 580244 191664 580256
rect 191694 580244 191739 580256
rect 191826 580244 194134 580800
rect 189443 580156 189477 580208
rect 189422 580128 189812 580156
rect 190101 580128 190135 580208
rect 190178 580128 190196 580202
rect 190228 580128 191601 580208
rect 191690 580206 194134 580244
rect 191694 580172 194134 580206
rect 191694 580156 191740 580172
rect 188920 580104 191601 580128
rect 191826 580104 194134 580172
rect 188920 580094 194134 580104
rect 189422 579624 189456 580094
rect 189636 580054 189683 580094
rect 189598 580020 189683 580054
rect 189525 579961 189570 579972
rect 189653 579961 189698 579972
rect 189536 579785 189570 579961
rect 189664 579785 189698 579961
rect 189636 579726 189683 579773
rect 189598 579692 189683 579726
rect 189656 579688 189662 579692
rect 189668 579652 189674 579688
rect 189778 579624 189812 580094
rect 189984 579936 189992 579966
rect 189956 579908 189992 579910
rect 189422 579590 189812 579624
rect 189408 578920 189830 579540
rect 190101 578924 190135 580094
rect 190178 579772 190196 580094
rect 190228 580070 194134 580094
rect 190206 579936 190222 579966
rect 190228 579910 191601 580070
rect 191688 580002 191692 580058
rect 190206 579908 191601 579910
rect 190178 579764 190194 579772
rect 190228 579646 191601 579908
rect 190228 579390 191610 579646
rect 191624 579418 191666 579618
rect 190036 578838 190135 578924
rect 189986 577974 190012 578778
rect 190014 577974 190040 578778
rect 190101 577974 190135 578838
rect 190178 578778 190180 579326
rect 190228 577974 191601 579390
rect 191826 579362 194134 580070
rect 194404 580736 196672 580806
rect 194404 579438 196676 580736
rect 194404 579368 196672 579438
rect 191936 579212 192148 579362
rect 192264 579178 192298 579362
rect 192322 579178 192332 579362
rect 192352 579332 192392 579362
rect 192402 579360 192420 579362
rect 192456 579360 192478 579362
rect 192484 579332 192506 579362
rect 192352 579318 192386 579332
rect 192398 579318 192423 579329
rect 192455 579318 192511 579329
rect 192352 579178 192423 579318
rect 192466 579178 192511 579318
rect 192580 579206 192816 579362
rect 192580 579178 192614 579206
rect 189428 577948 191601 577974
rect 189422 576550 189496 576880
rect 189422 576396 189628 576550
rect 189422 576226 189496 576396
rect 188773 575528 188831 575546
rect 189431 575528 189489 575546
rect 189986 575528 190012 577948
rect 190014 575528 190040 577948
rect 190101 575546 190135 577948
rect 190089 575528 190147 575546
rect 190228 575528 191601 577948
rect 191886 579144 192806 579178
rect 191886 577864 191920 579144
rect 192264 579076 192298 579144
rect 192322 579114 192332 579144
rect 192352 579142 192423 579144
rect 192466 579142 192511 579144
rect 192352 579130 192386 579142
rect 192392 579130 192406 579138
rect 192472 579130 192484 579138
rect 192352 579128 192494 579130
rect 192352 579114 192500 579128
rect 192580 579114 192614 579144
rect 192322 579076 192668 579114
rect 192062 579042 192668 579076
rect 191989 578992 192034 579003
rect 192000 578016 192034 578992
rect 192264 578990 192298 579042
rect 192322 579024 192332 579042
rect 192340 579024 192398 579042
rect 192322 579004 192398 579024
rect 192322 578996 192397 579004
rect 192326 578990 192397 578996
rect 192580 578990 192614 579042
rect 192647 578992 192703 579003
rect 192264 578956 192614 578990
rect 192352 578004 192397 578956
rect 192658 578016 192703 578992
rect 192322 577966 192668 578004
rect 192062 577932 192668 577966
rect 192340 577916 192398 577932
rect 192352 577864 192386 577916
rect 192772 577864 192806 579144
rect 192976 578778 193000 579326
rect 192888 578650 192898 578756
rect 192984 578652 192994 578756
rect 193004 577926 193028 579354
rect 193084 579178 193118 579362
rect 193198 579178 193243 579362
rect 193248 579212 193654 579362
rect 193248 579194 193460 579212
rect 193668 579178 193702 579362
rect 193782 579178 193816 579362
rect 197209 579234 197243 581110
rect 197590 581108 200100 581110
rect 197590 581038 198924 581108
rect 197918 580984 198924 581038
rect 197590 580630 198924 580984
rect 198946 580690 198984 581108
rect 199052 581096 199062 581108
rect 197590 580562 198910 580630
rect 197918 580238 198910 580562
rect 199108 580238 200100 581108
rect 197327 579234 197357 580221
rect 200418 580187 201410 581666
rect 201586 581642 204174 581674
rect 204368 581642 204402 581676
rect 205026 581642 205060 581676
rect 205684 581642 205718 581676
rect 205798 581642 205832 583516
rect 208744 581758 208782 584526
rect 208800 581814 208810 584526
rect 210297 581875 210496 585210
rect 215447 584691 215481 585315
rect 215533 585303 216178 585315
rect 215549 585232 216178 585303
rect 216228 585309 216284 585315
rect 216228 585280 216262 585309
rect 216760 585280 216794 585315
rect 218516 585287 218597 585321
rect 216228 585246 216794 585280
rect 215549 584759 215583 585232
rect 215926 584784 216056 584800
rect 216256 584784 217384 584800
rect 215954 584756 216056 584772
rect 216256 584756 217356 584772
rect 216778 584737 217356 584756
rect 218563 584743 218597 585287
rect 216778 584731 218242 584737
rect 218516 584731 218613 584743
rect 218665 584731 218699 585429
rect 215642 584725 223618 584731
rect 215413 584657 215481 584691
rect 215502 584703 215583 584704
rect 215502 584691 215617 584703
rect 215626 584697 223618 584725
rect 215502 584685 215583 584691
rect 215592 584685 218520 584691
rect 215502 584676 218520 584685
rect 215502 584663 218597 584676
rect 215502 584657 218515 584663
rect 215447 584033 215481 584657
rect 215533 584645 215630 584657
rect 215549 584101 215583 584645
rect 216056 584628 216256 584638
rect 218516 584629 218597 584663
rect 216028 584600 216284 584610
rect 218563 584085 218597 584629
rect 218516 584073 218613 584085
rect 215642 584067 218613 584073
rect 215413 583999 215481 584033
rect 215502 584045 215583 584046
rect 215626 584045 218613 584067
rect 215502 584033 215617 584045
rect 215626 584039 218554 584045
rect 215502 584027 215583 584033
rect 215592 584027 218520 584033
rect 215502 584018 218520 584027
rect 215502 584005 218597 584018
rect 215502 583999 218515 584005
rect 215447 583375 215481 583999
rect 215533 583987 215630 583999
rect 215549 583443 215583 583987
rect 218516 583971 218597 584005
rect 216864 583950 218216 583968
rect 216836 583922 218244 583940
rect 215904 583462 217362 583480
rect 215932 583434 217334 583452
rect 218563 583427 218597 583971
rect 218516 583415 218613 583427
rect 215642 583409 218613 583415
rect 215413 583341 215481 583375
rect 215502 583387 215583 583388
rect 215626 583387 218613 583409
rect 215502 583375 215617 583387
rect 215626 583381 218554 583387
rect 215502 583369 215583 583375
rect 215592 583369 218520 583375
rect 215502 583360 218520 583369
rect 215502 583347 218597 583360
rect 215502 583341 218515 583347
rect 215447 582643 215481 583341
rect 215533 583329 215630 583341
rect 215549 582785 215583 583329
rect 218516 583313 218597 583347
rect 218563 582769 218597 583313
rect 218516 582757 218613 582769
rect 215642 582751 218613 582757
rect 215626 582729 218613 582751
rect 215626 582723 218554 582729
rect 215592 582689 218520 582717
rect 215604 582685 218504 582689
rect 218563 582655 218597 582677
rect 218665 582643 218699 584697
rect 278928 583681 278962 584824
rect 280487 583681 280521 585385
rect 280963 585379 280997 585417
rect 284005 585395 284016 585406
rect 284028 585395 284039 585406
rect 284005 585379 284039 585395
rect 280663 585345 284339 585379
rect 280963 583681 280997 585345
rect 281066 585286 281122 585297
rect 281248 585286 281304 585297
rect 281724 585286 281780 585297
rect 281906 585286 281962 585297
rect 282382 585286 282427 585297
rect 282564 585286 282609 585297
rect 283040 585286 283085 585297
rect 283222 585286 283267 585297
rect 283698 585286 283743 585297
rect 283880 585286 283925 585297
rect 281077 585030 281798 585286
rect 281077 583681 281122 585030
rect 281138 583681 281166 584962
rect 281259 583681 281304 585030
rect 281735 583681 281780 585030
rect 281796 583681 281824 584962
rect 281852 583681 281880 584962
rect 281917 583681 281962 585286
rect 278619 583647 282171 583681
rect 223643 582735 223650 582808
rect 223677 582769 223684 582842
rect 215447 582609 223717 582643
rect 218665 582007 218699 582609
rect 266686 582380 266720 583112
rect 267458 582474 267492 582508
rect 268116 582474 268150 582508
rect 269288 582476 269298 582530
rect 269404 582476 269412 582510
rect 270036 582476 270070 582510
rect 270694 582476 270728 582510
rect 271352 582476 271386 582510
rect 271466 582476 271500 583118
rect 267238 582440 268816 582474
rect 266686 581938 266730 582380
rect 218080 581914 218338 581926
rect 266696 581658 266730 581938
rect 267238 581876 267272 582440
rect 267374 582304 267398 582406
rect 267458 582388 267505 582419
rect 267402 582372 267426 582378
rect 267446 582372 267505 582388
rect 267982 582372 268029 582419
rect 267402 582338 268029 582372
rect 267402 582332 267426 582338
rect 267446 582291 267504 582338
rect 268032 582304 268050 582406
rect 268116 582388 268163 582419
rect 268060 582372 268078 582378
rect 268104 582372 268163 582388
rect 268640 582372 268687 582419
rect 268782 582412 268816 582440
rect 268748 582378 268816 582412
rect 269342 582420 269352 582476
rect 269366 582442 272798 582476
rect 269366 582420 269376 582442
rect 268060 582338 268687 582372
rect 268060 582336 268078 582338
rect 268104 582336 268162 582338
rect 268060 582332 268162 582336
rect 268104 582308 268162 582332
rect 268080 582304 268162 582308
rect 267341 582279 267386 582290
rect 267352 582025 267386 582279
rect 267458 582037 267492 582291
rect 267999 582279 268044 582290
rect 268010 582025 268044 582279
rect 268052 582110 268074 582286
rect 268080 582082 268102 582304
rect 268104 582291 268162 582304
rect 268116 582037 268150 582291
rect 268657 582279 268702 582290
rect 268668 582025 268702 582279
rect 268782 582071 268842 582378
rect 268774 582037 268842 582071
rect 267340 581978 267399 582025
rect 267430 581984 267477 582025
rect 267422 581978 267477 581984
rect 267998 581978 268057 582025
rect 268088 581984 268135 582025
rect 268076 581978 268135 581984
rect 268656 581978 268714 582025
rect 267340 581944 267477 581978
rect 267520 581944 268135 581978
rect 268178 581944 268714 581978
rect 268748 581944 268762 581978
rect 267340 581928 267398 581944
rect 267422 581938 267442 581944
rect 267340 581913 267355 581928
rect 267450 581910 267470 581944
rect 267998 581928 268056 581944
rect 268076 581938 268100 581944
rect 268104 581910 268128 581944
rect 268656 581928 268714 581944
rect 268699 581913 268714 581928
rect 268782 581876 268816 582037
rect 269342 581882 269376 582420
rect 269378 582027 269410 582420
rect 270036 582390 270083 582421
rect 270024 582374 270083 582390
rect 270086 582374 270133 582421
rect 270694 582390 270741 582421
rect 270682 582374 270741 582390
rect 270744 582374 270791 582421
rect 271352 582390 271398 582421
rect 271340 582374 271398 582390
rect 271466 582374 271500 582442
rect 269518 582340 270133 582374
rect 270176 582340 270791 582374
rect 270834 582340 271398 582374
rect 271402 582340 271420 582374
rect 269422 582292 269446 582321
rect 270024 582293 270082 582340
rect 270682 582334 270756 582340
rect 270682 582314 270740 582334
rect 270682 582306 270766 582314
rect 270682 582293 270740 582306
rect 271340 582304 271398 582340
rect 271466 582315 271472 582347
rect 271476 582315 271500 582374
rect 271340 582293 271420 582304
rect 269450 582292 269474 582293
rect 269422 582281 269490 582292
rect 269422 582038 269446 582281
rect 269450 582031 269490 582281
rect 270036 582074 270076 582293
rect 270103 582288 270148 582292
rect 270086 582281 270148 582288
rect 270086 582102 270104 582281
rect 270036 582043 270070 582074
rect 270114 582031 270148 582281
rect 270694 582043 270728 582293
rect 270761 582281 270806 582292
rect 270772 582031 270806 582281
rect 271352 582054 271392 582293
rect 271396 582082 271420 582293
rect 271352 582043 271386 582054
rect 269444 581984 269503 582031
rect 270008 581984 270055 582031
rect 270102 581984 270161 582031
rect 270666 581984 270713 582031
rect 270760 581984 270819 582031
rect 271324 581984 271371 582031
rect 269444 581950 270055 581984
rect 270098 581950 270713 581984
rect 270756 581950 271371 581984
rect 269444 581934 269502 581950
rect 270102 581934 270160 581950
rect 270760 581934 270818 581950
rect 269444 581919 269459 581934
rect 271430 581882 271438 581916
rect 271466 581882 271500 582315
rect 266782 581842 268826 581876
rect 269342 581848 271500 581882
rect 267238 581738 267272 581842
rect 267132 581718 267794 581738
rect 267174 581698 267740 581718
rect 267238 581694 267272 581698
rect 267202 581670 267740 581694
rect 267238 581658 267272 581670
rect 268782 581658 268816 581842
rect 269342 581666 269376 581848
rect 201586 581608 206238 581642
rect 201586 581540 204174 581608
rect 204184 581540 204222 581578
rect 204368 581556 204406 581578
rect 204356 581540 204414 581556
rect 204842 581540 204880 581578
rect 205026 581556 205064 581578
rect 205014 581540 205072 581556
rect 205500 581540 205538 581578
rect 205684 581571 205722 581578
rect 205684 581556 205730 581571
rect 205672 581540 205730 581556
rect 201586 581506 204222 581540
rect 204274 581506 204880 581540
rect 204932 581506 205538 581540
rect 205590 581506 205730 581540
rect 201586 580223 204174 581506
rect 204201 581456 204246 581467
rect 204212 580223 204246 581456
rect 204250 580223 204284 581500
rect 204306 580223 204340 581500
rect 204356 581468 204414 581506
rect 204368 580223 204402 581468
rect 204859 581456 204904 581467
rect 204870 580223 204904 581456
rect 204908 580223 204948 581500
rect 204964 580223 205004 581500
rect 205014 581468 205072 581506
rect 205026 580223 205060 581468
rect 205517 581456 205562 581467
rect 205528 580223 205562 581456
rect 205628 580223 205656 581500
rect 205672 581468 205730 581506
rect 205684 580223 205718 581468
rect 201586 580187 205763 580223
rect 197361 580153 205763 580187
rect 197361 579234 197395 580153
rect 197912 580073 197969 580084
rect 197981 580073 198015 580153
rect 198605 580106 198610 580108
rect 198633 580106 198638 580136
rect 198027 580078 198627 580084
rect 198639 580078 198673 580153
rect 199297 580134 199337 580153
rect 199263 580084 199282 580106
rect 198685 580078 198912 580084
rect 198027 580073 198926 580078
rect 199110 580073 199285 580084
rect 199291 580079 199337 580134
rect 199344 580084 199365 580138
rect 199297 580073 199331 580079
rect 199343 580073 199943 580084
rect 199955 580073 199989 580153
rect 200418 580094 201410 580153
rect 201438 580122 205763 580153
rect 201438 580094 201472 580122
rect 200001 580073 200110 580084
rect 200418 580073 201506 580094
rect 201586 580088 205763 580122
rect 201580 580086 205763 580088
rect 201567 580073 205763 580086
rect 197416 580011 197497 580058
rect 197556 580039 205763 580073
rect 197968 580027 197969 580028
rect 197981 580027 198015 580039
rect 198027 580027 198028 580028
rect 197969 580026 197970 580027
rect 197981 580026 198027 580027
rect 197463 579443 197497 580011
rect 197981 579428 198026 580026
rect 198224 580018 198926 580039
rect 199297 580033 199331 580039
rect 198088 579958 198098 579984
rect 198060 579930 198098 579956
rect 198224 579806 198582 580018
rect 198605 579956 198610 579998
rect 198633 579956 198638 579998
rect 198639 579428 198684 580018
rect 199263 579998 199282 580033
rect 199284 580027 199285 580028
rect 199291 580027 199337 580033
rect 199344 580028 199365 580033
rect 199343 580027 199365 580028
rect 199942 580027 199943 580028
rect 199955 580027 199989 580039
rect 200001 580027 200002 580028
rect 199285 580026 199286 580027
rect 199291 580026 199343 580027
rect 199291 579970 199342 580026
rect 199297 579428 199342 579970
rect 199344 579956 199365 580027
rect 199943 580026 199944 580027
rect 199955 580026 200001 580027
rect 199955 579428 200000 580026
rect 200418 579854 201410 580039
rect 201438 579854 201472 580039
rect 201586 579972 205763 580039
rect 201541 579961 205763 579972
rect 201552 579854 205763 579961
rect 200418 579654 205763 579854
rect 200418 579646 201734 579654
rect 197969 579427 197970 579428
rect 197981 579427 198027 579428
rect 198627 579427 198628 579428
rect 198639 579427 198685 579428
rect 199285 579427 199286 579428
rect 199297 579427 199343 579428
rect 199943 579427 199944 579428
rect 199955 579427 200001 579428
rect 200586 579427 200658 579646
rect 200700 579508 200761 579646
rect 200776 579518 201046 579646
rect 201286 579642 201734 579646
rect 200700 579504 200768 579508
rect 197968 579426 197969 579427
rect 197912 579415 197969 579426
rect 197981 579415 198015 579427
rect 198027 579426 198028 579427
rect 198626 579426 198627 579427
rect 198027 579415 198627 579426
rect 198639 579415 198673 579427
rect 198685 579426 198686 579427
rect 199284 579426 199285 579427
rect 198685 579415 198912 579426
rect 199110 579415 199285 579426
rect 199297 579415 199331 579427
rect 199343 579426 199344 579427
rect 199942 579426 199943 579427
rect 199343 579415 199943 579426
rect 199955 579415 199989 579427
rect 200001 579426 200002 579427
rect 200586 579426 200654 579427
rect 200001 579415 200110 579426
rect 200404 579415 200654 579426
rect 200700 579426 200761 579504
rect 201358 579428 201403 579642
rect 201404 579556 201416 579642
rect 201438 579624 201472 579642
rect 201794 579624 201828 579654
rect 202016 579640 202061 579654
rect 202244 579640 205763 579654
rect 201438 579590 201828 579624
rect 201346 579427 201347 579428
rect 201358 579427 201404 579428
rect 201345 579426 201346 579427
rect 200700 579415 201346 579426
rect 201358 579415 201392 579427
rect 201404 579426 201405 579427
rect 201424 579426 201846 579540
rect 201920 579462 205763 579640
rect 201946 579436 202010 579449
rect 201920 579426 201946 579436
rect 201976 579430 202010 579436
rect 202016 579430 202106 579462
rect 202016 579428 202061 579430
rect 202004 579427 202005 579428
rect 202016 579427 202062 579428
rect 202003 579426 202004 579427
rect 201404 579415 201416 579426
rect 201424 579421 202004 579426
rect 202016 579421 202056 579427
rect 202062 579426 202063 579427
rect 202244 579426 205763 579462
rect 202062 579421 205763 579426
rect 201424 579415 202010 579421
rect 202016 579415 202050 579421
rect 202056 579415 205763 579421
rect 197416 579353 197497 579400
rect 197556 579381 205763 579415
rect 197968 579369 197969 579370
rect 197981 579369 198015 579381
rect 198027 579369 198028 579370
rect 198626 579369 198627 579370
rect 198639 579369 198673 579381
rect 198685 579369 198686 579370
rect 199284 579369 199285 579370
rect 199297 579369 199331 579381
rect 199343 579369 199344 579370
rect 199942 579369 199943 579370
rect 199955 579369 199989 579381
rect 200001 579369 200002 579370
rect 200586 579369 200654 579381
rect 197969 579368 197970 579369
rect 197981 579368 198027 579369
rect 198627 579368 198628 579369
rect 198639 579368 198685 579369
rect 199285 579368 199286 579369
rect 199297 579368 199343 579369
rect 199943 579368 199944 579369
rect 199955 579368 200001 579369
rect 197463 579234 197497 579353
rect 197981 579234 198026 579368
rect 198542 579298 198546 579348
rect 198570 579298 198574 579320
rect 198639 579234 198684 579368
rect 199297 579234 199342 579368
rect 199955 579234 200000 579368
rect 193856 579178 193890 579212
rect 194514 579186 194548 579220
rect 195172 579186 195206 579220
rect 195830 579194 195864 579228
rect 193076 579144 193996 579178
rect 193042 579082 193044 579116
rect 191886 577830 192806 577864
rect 193076 577864 193118 579144
rect 193198 579092 193243 579144
rect 193668 579114 193702 579144
rect 193198 579004 193244 579092
rect 193668 579076 193706 579114
rect 193782 579076 193816 579144
rect 193856 579138 193890 579144
rect 193850 579114 193890 579138
rect 193820 579076 193890 579114
rect 193252 579042 193890 579076
rect 193198 579003 193243 579004
rect 193179 578992 193243 579003
rect 193190 578016 193243 578992
rect 193198 578004 193243 578016
rect 193668 578004 193702 579042
rect 193782 578338 193816 579042
rect 193822 579036 193832 579042
rect 193850 579008 193890 579042
rect 193848 579004 193890 579008
rect 193842 579003 193890 579004
rect 193837 578992 193890 579003
rect 193842 578980 193890 578992
rect 193782 578028 193838 578338
rect 193848 578028 193890 578980
rect 193198 577916 193244 578004
rect 193668 577966 193706 578004
rect 193782 577966 193816 578028
rect 193842 578004 193890 578028
rect 193820 577966 193890 578004
rect 193252 577932 193890 577966
rect 193198 577864 193243 577916
rect 193668 577868 193702 577932
rect 193668 577864 193713 577868
rect 193782 577864 193816 577932
rect 193822 577926 193832 577932
rect 193850 577870 193890 577932
rect 193856 577864 193890 577870
rect 193962 577864 193996 579144
rect 193076 577830 193996 577864
rect 194386 579152 195306 579186
rect 191652 576638 191666 577216
rect 191652 576582 191692 576638
rect 192352 576584 192386 577830
rect 192484 576584 192524 576632
rect 192946 576584 192972 577208
rect 192974 576584 193000 577180
rect 193080 576584 193082 577180
rect 193084 576584 193118 577830
rect 193198 576584 193243 577830
rect 193668 576584 193713 577830
rect 193782 576584 193816 577830
rect 194386 577272 194420 579152
rect 194514 579100 194548 579152
rect 195130 579118 195168 579122
rect 194424 578750 194430 579036
rect 194514 579012 194560 579100
rect 195130 579084 195170 579118
rect 194562 579050 195170 579084
rect 195138 579044 195142 579050
rect 195166 579016 195170 579050
rect 194452 578778 194458 579008
rect 194489 579000 194502 579011
rect 194514 579000 194548 579012
rect 195147 579000 195160 579011
rect 195172 579000 195206 579152
rect 194500 577424 194548 579000
rect 195158 577424 195206 579000
rect 194514 577412 194548 577424
rect 194514 577324 194560 577412
rect 195130 577408 195168 577412
rect 195130 577374 195170 577408
rect 194562 577340 195170 577374
rect 195138 577334 195142 577340
rect 194514 577272 194548 577324
rect 195166 577306 195170 577340
rect 195172 577272 195206 577424
rect 195272 577272 195306 579152
rect 194386 577238 195306 577272
rect 195554 579160 196474 579194
rect 195554 577280 195588 579160
rect 195830 579108 195868 579130
rect 195818 579092 195876 579108
rect 196298 579092 196336 579130
rect 195730 579058 196336 579092
rect 195698 579019 195752 579052
rect 195657 579008 195752 579019
rect 195668 577432 195752 579008
rect 195698 577388 195752 577432
rect 195754 577388 195780 579052
rect 195818 579020 195876 579058
rect 195830 577420 195864 579020
rect 196315 579008 196360 579019
rect 196326 577432 196360 579008
rect 195818 577382 195876 577420
rect 196298 577382 196336 577420
rect 195730 577348 196336 577382
rect 195818 577332 195876 577348
rect 195830 577280 195864 577332
rect 196440 577280 196474 579160
rect 196488 577286 196508 579228
rect 197173 578757 200302 579234
rect 200586 578769 200658 579369
rect 200586 578768 200654 578769
rect 200404 578757 200654 578768
rect 200700 578768 200761 579381
rect 201345 579369 201346 579370
rect 201358 579369 201392 579381
rect 201404 579369 201405 579370
rect 201346 579368 201347 579369
rect 201358 579368 201404 579369
rect 201358 578770 201403 579368
rect 201424 578920 201846 579381
rect 201920 579375 202010 579381
rect 202016 579375 202050 579381
rect 202056 579375 202106 579381
rect 202003 579369 202004 579370
rect 202016 579369 202056 579375
rect 202062 579369 202063 579370
rect 202004 579368 202005 579369
rect 202016 579368 202062 579369
rect 202016 579326 202061 579368
rect 202016 579319 202106 579326
rect 202016 578924 202061 579319
rect 202016 578838 202088 578924
rect 201456 578778 201576 578791
rect 201988 578778 202010 578791
rect 202016 578770 202061 578838
rect 201346 578769 201347 578770
rect 201358 578769 201404 578770
rect 202004 578769 202005 578770
rect 202016 578769 202062 578770
rect 201345 578768 201346 578769
rect 200700 578757 201346 578768
rect 201358 578757 201392 578769
rect 201404 578768 201405 578769
rect 202003 578768 202004 578769
rect 201404 578757 201416 578768
rect 201576 578763 202004 578768
rect 201576 578757 202010 578763
rect 202016 578757 202050 578769
rect 202062 578768 202063 578769
rect 202244 578768 205763 579381
rect 202062 578757 205763 578768
rect 197173 578723 205763 578757
rect 197173 578110 200302 578723
rect 200586 578717 200694 578723
rect 200700 578717 200792 578723
rect 200586 578711 200654 578717
rect 200586 578698 200658 578711
rect 200700 578698 200761 578717
rect 201345 578711 201346 578712
rect 201358 578711 201392 578723
rect 201404 578711 201405 578712
rect 202003 578711 202004 578712
rect 202016 578711 202050 578723
rect 202062 578711 202063 578712
rect 201346 578710 201347 578711
rect 201358 578710 201404 578711
rect 202004 578710 202005 578711
rect 202016 578710 202062 578711
rect 200586 578689 200694 578698
rect 200700 578689 200764 578698
rect 200586 578636 200681 578689
rect 200586 578144 200658 578636
rect 200700 578305 200761 578689
rect 201358 578305 201403 578710
rect 202016 578305 202061 578710
rect 200727 578293 200761 578305
rect 202244 578293 205763 578723
rect 200715 578246 201377 578293
rect 201576 578246 205763 578293
rect 200727 578144 200761 578246
rect 200762 578212 201377 578246
rect 201420 578234 202035 578246
rect 202078 578234 205763 578246
rect 201420 578230 205763 578234
rect 205798 578230 205832 581608
rect 206180 579182 206182 579421
rect 206186 578280 206220 581456
rect 266674 581074 266766 581658
rect 267202 581262 267666 581658
rect 267202 581072 267680 581262
rect 267684 581210 267740 581228
rect 267794 581210 267846 581228
rect 215470 579422 215504 580994
rect 223648 580318 223650 580942
rect 223682 580330 223684 580930
rect 267642 580630 267680 581072
rect 267702 580690 267740 581202
rect 267794 581182 267818 581200
rect 267864 581072 268852 581658
rect 216252 579678 216604 579764
rect 216252 579660 217000 579678
rect 223648 579660 223650 580284
rect 223682 579672 223684 580272
rect 215776 579626 223632 579660
rect 269306 579646 270166 581666
rect 270342 579654 271334 581674
rect 271502 581444 272930 581678
rect 271502 581116 272952 581444
rect 216252 579604 217000 579626
rect 216252 579490 216604 579604
rect 214744 579388 218200 579422
rect 215470 579354 215504 579388
rect 215448 579320 215504 579354
rect 215572 579320 215606 579388
rect 216050 579320 216088 579358
rect 216708 579320 216746 579358
rect 217366 579320 217404 579358
rect 218024 579320 218062 579358
rect 215470 579286 216088 579320
rect 216140 579286 216746 579320
rect 216798 579286 217404 579320
rect 217456 579286 218062 579320
rect 215452 579244 215460 579248
rect 215470 579244 215504 579286
rect 215386 579182 215412 579244
rect 215452 579182 215504 579244
rect 212332 578494 212349 578526
rect 212332 578424 212350 578494
rect 201420 578212 206842 578230
rect 201956 578210 206842 578212
rect 202244 578206 206842 578210
rect 201426 578188 201682 578204
rect 201956 578196 206842 578206
rect 201454 578160 201654 578176
rect 201956 578154 205763 578196
rect 202244 578144 205763 578154
rect 200586 578128 205763 578144
rect 205798 578128 205832 578196
rect 200586 578110 206238 578128
rect 197173 578099 200601 578110
rect 200613 578099 200647 578110
rect 200727 578099 200761 578110
rect 197173 578065 200795 578099
rect 202244 578094 206238 578110
rect 197173 577441 200302 578065
rect 200600 578053 200601 578054
rect 200613 578053 200647 578065
rect 200601 578052 200602 578053
rect 200613 577626 200658 578053
rect 200601 577453 200602 577454
rect 200600 577452 200601 577453
rect 200613 577441 200647 577626
rect 200727 577441 200761 578065
rect 201454 577976 201654 577994
rect 201426 577948 201682 577966
rect 197173 577407 200761 577441
rect 195554 577246 196474 577280
rect 193866 576652 193890 576810
rect 193904 576690 193928 576772
rect 194200 576584 194662 576716
rect 194676 576584 195138 576716
rect 195738 576588 195752 577236
rect 195830 576588 195864 577246
rect 196790 576690 196810 576772
rect 196828 576652 196848 576810
rect 197173 576794 200302 577407
rect 200600 577395 200601 577396
rect 200601 577394 200602 577395
rect 200613 577028 200647 577407
rect 200601 576795 200602 576796
rect 200613 576795 200658 577028
rect 200600 576794 200601 576795
rect 197173 576783 200601 576794
rect 200613 576783 200647 576795
rect 200727 576783 200761 577407
rect 202244 576842 205763 578094
rect 197173 576749 200795 576783
rect 200797 576749 205763 576842
rect 205798 576749 205832 578094
rect 213772 577786 213830 577816
rect 213806 577752 213830 577782
rect 211274 577580 211656 577680
rect 210488 577208 211668 577580
rect 215470 577572 215504 579182
rect 215572 579030 215606 579286
rect 215644 579248 215645 579249
rect 215643 579247 215644 579248
rect 216067 579236 216112 579247
rect 216725 579236 216770 579247
rect 217383 579236 217428 579247
rect 218041 579236 218086 579247
rect 216066 579014 216067 579015
rect 216065 579013 216066 579014
rect 216078 579002 216112 579236
rect 216123 579014 216124 579015
rect 216724 579014 216725 579015
rect 216124 579013 216125 579014
rect 216723 579013 216724 579014
rect 216736 579002 216770 579236
rect 216781 579014 216782 579015
rect 217382 579014 217383 579015
rect 216782 579013 216783 579014
rect 217381 579013 217382 579014
rect 217394 579002 217428 579236
rect 217439 579014 217440 579015
rect 218040 579014 218041 579015
rect 217440 579013 217441 579014
rect 218039 579013 218040 579014
rect 218052 579002 218086 579236
rect 218166 579002 218200 579388
rect 222904 579086 222960 579098
rect 223648 579002 223650 579626
rect 223682 579014 223684 579614
rect 269482 579476 269496 579646
rect 269510 579504 269524 579646
rect 215534 578940 215606 578978
rect 215656 578968 218200 579002
rect 216065 578956 216066 578957
rect 216066 578955 216067 578956
rect 215572 578528 215606 578940
rect 216078 578528 216112 578968
rect 216124 578956 216125 578957
rect 216723 578956 216724 578957
rect 216123 578955 216124 578956
rect 216724 578955 216725 578956
rect 216736 578528 216770 578968
rect 216782 578956 216783 578957
rect 217381 578956 217382 578957
rect 216781 578955 216782 578956
rect 217382 578955 217383 578956
rect 217394 578528 217428 578968
rect 217440 578956 217441 578957
rect 218039 578956 218040 578957
rect 217439 578955 217440 578956
rect 218040 578955 218041 578956
rect 215572 578372 215644 578528
rect 216078 578357 216123 578528
rect 216736 578434 216781 578528
rect 217394 578434 217439 578528
rect 216286 578362 217466 578434
rect 216338 578357 217439 578362
rect 216066 578356 216067 578357
rect 216078 578356 216124 578357
rect 216338 578356 217440 578357
rect 218040 578356 218041 578357
rect 216065 578355 216066 578356
rect 215645 578344 216066 578355
rect 216078 578344 216112 578356
rect 216124 578355 216125 578356
rect 216338 578355 217428 578356
rect 216124 578344 217428 578355
rect 217440 578355 217441 578356
rect 218039 578355 218040 578356
rect 217440 578344 217984 578355
rect 218052 578344 218086 578968
rect 218166 578344 218200 578968
rect 222904 578906 222960 578926
rect 222904 578850 222960 578870
rect 223648 578344 223650 578968
rect 223682 578406 223684 578956
rect 223676 578384 223700 578406
rect 223676 578360 223722 578384
rect 223682 578356 223684 578360
rect 215534 578282 215644 578320
rect 215656 578310 223632 578344
rect 216065 578298 216066 578299
rect 216078 578298 216112 578310
rect 216124 578298 216125 578299
rect 216338 578298 217428 578310
rect 217440 578298 217441 578299
rect 218039 578298 218040 578299
rect 216066 578297 216067 578298
rect 216078 578297 216124 578298
rect 216338 578297 217440 578298
rect 218040 578297 218041 578298
rect 215572 577714 215644 578282
rect 216078 577699 216123 578297
rect 216338 578288 217439 578297
rect 216286 578062 217466 578288
rect 216736 577699 216781 578062
rect 217394 577699 217439 578062
rect 216066 577698 216067 577699
rect 216078 577698 216124 577699
rect 216724 577698 216725 577699
rect 216736 577698 216782 577699
rect 217382 577698 217383 577699
rect 217394 577698 217440 577699
rect 216065 577697 216066 577698
rect 215645 577686 216066 577697
rect 216078 577686 216112 577698
rect 216124 577697 216125 577698
rect 216723 577697 216724 577698
rect 216124 577686 216724 577697
rect 216736 577686 216770 577698
rect 216782 577697 216783 577698
rect 217381 577697 217382 577698
rect 216782 577686 217382 577697
rect 217394 577686 217428 577698
rect 217440 577697 217441 577698
rect 218018 577697 218042 577782
rect 217440 577686 218042 577697
rect 218052 577686 218086 578310
rect 218166 577686 218200 578310
rect 223648 577686 223650 578310
rect 223682 577698 223684 578298
rect 268840 578138 268866 579062
rect 268874 578138 268900 579028
rect 270772 578305 270806 579654
rect 271476 578212 271492 578246
rect 271502 578074 272930 581116
rect 278619 580588 278653 583647
rect 278814 583595 278860 583626
rect 278802 583579 278860 583595
rect 278795 583545 278860 583579
rect 278802 583498 278860 583545
rect 278722 583486 278767 583497
rect 278733 580737 278767 583486
rect 278814 580749 278848 583498
rect 278721 580690 278780 580737
rect 278786 580690 278833 580737
rect 278721 580656 278833 580690
rect 278721 580640 278779 580656
rect 278721 580625 278736 580640
rect 278733 580588 278767 580622
rect 278928 580588 278962 583647
rect 276256 580554 278962 580588
rect 215656 577652 218200 577686
rect 216078 577572 216112 577652
rect 216736 577572 216770 577652
rect 217394 577572 217428 577652
rect 218052 577572 218086 577652
rect 218166 577572 218200 577652
rect 215470 577538 223722 577572
rect 212284 577244 213276 577256
rect 213452 577238 214444 577256
rect 197173 576716 200302 576749
rect 197020 576669 200302 576716
rect 200613 576669 200647 576749
rect 200727 576669 200761 576749
rect 200797 576713 205868 576749
rect 200797 576679 207119 576713
rect 200797 576669 205868 576679
rect 197020 576635 205868 576669
rect 206348 576658 206546 576679
rect 206344 576649 206546 576658
rect 206824 576649 207022 576679
rect 191624 576382 191636 576582
rect 191652 576382 191664 576582
rect 191652 576326 191692 576382
rect 191652 576238 191666 576326
rect 191652 576182 191692 576238
rect 191624 575982 191636 576182
rect 191652 575982 191664 576182
rect 191758 576078 195138 576584
rect 195248 576136 195260 576456
rect 195270 576420 196672 576588
rect 196678 576420 196920 576588
rect 191758 576044 194724 576078
rect 191652 575926 191692 575982
rect 191652 575814 191666 575926
rect 191752 575854 194724 576044
rect 191724 575814 194724 575854
rect 191724 575798 191728 575814
rect 191758 575646 194724 575814
rect 194730 575994 195080 576028
rect 191688 575546 191692 575582
rect 187626 575492 191601 575528
rect 191682 575512 191740 575546
rect 192340 575512 192398 575546
rect 187626 575487 192982 575492
rect 187626 575481 191693 575487
rect 191729 575481 192351 575487
rect 192387 575481 192982 575487
rect 187626 575469 191682 575481
rect 191740 575469 192340 575481
rect 192398 575469 192982 575481
rect 187626 575458 191693 575469
rect 191729 575458 192351 575469
rect 192387 575458 192982 575469
rect 186618 575349 187588 575450
rect 187626 575448 191601 575458
rect 187626 575424 191682 575448
rect 191740 575424 192340 575448
rect 192398 575424 192864 575448
rect 192948 575424 192982 575458
rect 187626 575406 191601 575424
rect 192484 575416 192846 575424
rect 187626 575396 192806 575406
rect 187626 575390 192818 575396
rect 187626 575372 191601 575390
rect 192456 575388 192818 575390
rect 192806 575372 192818 575388
rect 192834 575372 192846 575416
rect 192948 575413 192959 575424
rect 192971 575413 192982 575424
rect 193084 575474 193118 575646
rect 193198 575524 193243 575646
rect 193668 575524 193713 575646
rect 193782 575474 193816 575646
rect 194254 575514 194288 575646
rect 194374 575616 194484 575646
rect 194514 575628 194528 575646
rect 194412 575582 194484 575616
rect 194514 575524 194542 575548
rect 194570 575514 194604 575646
rect 193852 575480 193868 575508
rect 194254 575480 194604 575514
rect 194730 575514 194764 575994
rect 194850 575926 194960 575964
rect 194888 575892 194960 575926
rect 194833 575842 194889 575853
rect 194921 575842 194977 575853
rect 194844 575666 194889 575842
rect 194932 575666 194977 575842
rect 194850 575616 194960 575654
rect 194888 575582 194960 575616
rect 195046 575514 195080 575994
rect 195248 575662 195260 575950
rect 195270 575684 196920 576420
rect 197020 576552 200302 576635
rect 200727 576552 200761 576635
rect 200797 576599 205868 576635
rect 206252 576646 206642 576649
rect 206252 576618 206286 576646
rect 206316 576618 206332 576630
rect 206218 576617 206332 576618
rect 206344 576617 206360 576646
rect 206218 576611 206320 576617
rect 202244 576584 203084 576588
rect 203627 576584 205868 576599
rect 202244 576552 205868 576584
rect 206252 576552 206286 576611
rect 206370 576594 206397 576627
rect 206508 576617 206530 576646
rect 206536 576617 206558 576630
rect 206608 576618 206642 576646
rect 206728 576646 207077 576649
rect 206728 576618 206762 576646
rect 206574 576611 206676 576618
rect 206694 576611 206796 576618
rect 206952 576617 206984 576630
rect 207008 576617 207012 576646
rect 206332 576571 206344 576584
rect 206412 576578 206439 576594
rect 206316 576552 206332 576571
rect 206344 576552 206360 576571
rect 206412 576552 206466 576578
rect 206471 576577 206504 576611
rect 206530 576571 206536 576584
rect 206508 576552 206530 576571
rect 206536 576552 206558 576571
rect 206608 576552 206642 576611
rect 206728 576577 207039 576611
rect 206728 576552 206762 576577
rect 206904 576552 206942 576577
rect 206984 576571 207008 576577
rect 206952 576552 206984 576571
rect 207008 576552 207012 576571
rect 207084 576552 207109 576584
rect 197020 576518 207032 576552
rect 197020 576078 200302 576518
rect 200613 576466 200659 576497
rect 200601 576450 200659 576466
rect 200330 576416 200659 576450
rect 200601 576369 200659 576416
rect 197173 576028 200302 576078
rect 197074 575994 200302 576028
rect 197074 575684 197108 575994
rect 197173 575694 200302 575994
rect 200613 575694 200647 576369
rect 197173 575684 200313 575694
rect 194730 575480 195080 575514
rect 195270 575650 200313 575684
rect 195270 575614 196920 575650
rect 193084 575440 193816 575474
rect 193824 575452 193840 575480
rect 193918 575448 194486 575474
rect 193918 575440 194488 575448
rect 193084 575424 193118 575440
rect 193084 575413 193095 575424
rect 193107 575413 193118 575424
rect 193782 575424 193816 575440
rect 193782 575413 193793 575424
rect 193805 575413 193816 575424
rect 194536 575406 194552 575480
rect 194564 575434 194580 575480
rect 192948 575372 192982 575396
rect 195270 575372 196854 575614
rect 197074 575576 197108 575650
rect 197173 575614 200313 575650
rect 187626 575364 196854 575372
rect 197173 575444 197460 575614
rect 197506 575498 197936 575614
rect 197981 575510 198026 575614
rect 198164 575498 198209 575614
rect 198639 575510 198684 575614
rect 198732 575498 198756 575614
rect 198760 575498 198812 575614
rect 198822 575498 198867 575614
rect 197494 575451 198868 575498
rect 187626 575349 196672 575364
rect 185193 575338 196672 575349
rect 180188 575318 180246 575338
rect 180846 575318 180904 575338
rect 173005 575288 173024 575302
rect 173121 575026 173144 575182
rect 172944 574982 173144 575026
rect 173149 574970 173172 575210
rect 173748 575164 175230 575315
rect 172916 574954 173172 574970
rect 173156 574404 173189 574448
rect 173190 574438 173223 574448
rect 173813 572996 173847 575164
rect 173874 574872 173898 574974
rect 173918 574332 173952 575164
rect 174032 574493 174077 575164
rect 174471 574481 174516 575164
rect 175129 574481 175174 575164
rect 175787 574481 175832 575315
rect 176090 574493 176124 575315
rect 174047 574434 175874 574481
rect 176062 574434 176109 574481
rect 174094 574400 176109 574434
rect 174459 574384 174517 574400
rect 175117 574384 175175 574400
rect 175775 574384 175833 574400
rect 174471 574332 174505 574366
rect 175129 574332 175163 574366
rect 175787 574332 175821 574366
rect 176204 574332 176238 575315
rect 173918 574298 176238 574332
rect 176559 574070 176593 575315
rect 177478 575279 179109 575315
rect 178112 574378 178146 575279
rect 178226 574518 178260 575279
rect 178884 574518 178918 575279
rect 179542 574518 179576 575318
rect 180200 574518 180245 575318
rect 180858 574518 180903 575318
rect 181468 574970 181488 575338
rect 181504 575318 181562 575338
rect 181258 574528 181262 574848
rect 181296 574528 181300 574848
rect 181516 574518 181561 575318
rect 178214 574480 178272 574518
rect 178872 574480 178930 574518
rect 179530 574480 179588 574518
rect 180114 574480 181562 574518
rect 178214 574446 181562 574480
rect 178214 574430 178272 574446
rect 178872 574430 178930 574446
rect 179530 574430 179588 574446
rect 180188 574430 180246 574446
rect 180846 574430 180904 574446
rect 181504 574430 181562 574446
rect 178214 574415 178229 574430
rect 181547 574415 181562 574430
rect 178226 574378 178260 574412
rect 178884 574378 178918 574412
rect 179542 574378 179576 574412
rect 180200 574378 180234 574412
rect 180858 574378 180892 574412
rect 181516 574378 181550 574412
rect 181630 574378 181664 575338
rect 182674 575313 182732 575318
rect 182800 574440 182834 575338
rect 184030 575302 184180 575338
rect 185193 575315 191601 575338
rect 192834 575322 192846 575338
rect 184066 574394 184100 575302
rect 184146 574546 184158 575302
rect 184180 574580 184192 575302
rect 184146 574443 184172 574546
rect 184180 574477 184206 574580
rect 186352 574394 186386 575315
rect 186618 575279 187588 575315
rect 187626 575279 191601 575315
rect 192822 575313 192880 575318
rect 191436 575182 191464 575279
rect 187062 575018 187134 575026
rect 187062 575016 187130 575018
rect 192948 574876 192982 575338
rect 195270 575302 196672 575338
rect 195734 575288 195896 575290
rect 197173 575279 197174 575444
rect 197345 575383 197372 575444
rect 197373 575411 197426 575444
rect 197392 575366 197426 575411
rect 197494 575417 198000 575451
rect 198043 575417 198658 575451
rect 197494 575404 197552 575417
rect 197494 575394 197572 575404
rect 198152 575394 198210 575417
rect 197456 575372 197572 575394
rect 198102 575388 198258 575394
rect 197494 575367 197552 575372
rect 198152 575367 198210 575388
rect 198663 575379 198670 575451
rect 198701 575417 198868 575451
rect 198810 575411 198868 575417
rect 198732 575376 198756 575411
rect 198760 575404 198868 575411
rect 198794 575394 198868 575404
rect 198794 575378 198888 575394
rect 198796 575370 198886 575378
rect 198810 575367 198868 575370
rect 197384 575354 197604 575366
rect 198102 575354 198258 575366
rect 198756 575355 198760 575366
rect 198766 575354 198916 575366
rect 197384 575350 198916 575354
rect 197384 575349 198914 575350
rect 198936 575349 198970 575614
rect 199496 575366 199530 575614
rect 199610 575498 199655 575614
rect 199955 575510 200000 575614
rect 200268 575498 200313 575614
rect 200613 575510 200658 575694
rect 199598 575451 200632 575498
rect 199598 575417 199974 575451
rect 200017 575417 200632 575451
rect 199598 575401 199656 575417
rect 200256 575401 200314 575417
rect 199598 575386 199613 575401
rect 199374 575349 199604 575366
rect 199610 575349 199644 575383
rect 199650 575349 199710 575366
rect 200206 575349 200262 575366
rect 200268 575349 200302 575383
rect 200308 575349 200360 575366
rect 200727 575349 200761 576518
rect 201490 576410 201644 576518
rect 202038 576514 205868 576518
rect 202244 576497 205868 576514
rect 206252 576497 206286 576518
rect 206409 576497 206455 576518
rect 206608 576497 206642 576518
rect 206728 576497 206762 576518
rect 206984 576515 207032 576518
rect 201942 576466 201953 576477
rect 201965 576466 201976 576477
rect 201942 576450 201976 576466
rect 202244 576450 206796 576497
rect 206842 576496 206889 576497
rect 206998 576496 207032 576515
rect 206831 576485 206889 576496
rect 206959 576485 207032 576496
rect 206842 576484 206889 576485
rect 206842 576450 206890 576484
rect 201942 576446 202214 576450
rect 202244 576446 206245 576450
rect 201942 576416 206245 576446
rect 201490 576396 201664 576410
rect 201632 576376 201664 576396
rect 201632 576358 201658 576376
rect 197305 575320 200761 575349
rect 197305 575315 198174 575320
rect 198188 575315 200761 575320
rect 197392 575280 197426 575315
rect 198226 575286 198794 575315
rect 198936 575280 198970 575315
rect 195772 575250 195858 575252
rect 196050 575186 196548 575214
rect 199496 575152 199530 575315
rect 200926 575152 200960 576357
rect 201560 576192 201658 576358
rect 201688 576353 201692 576410
rect 201560 576178 201638 576192
rect 201558 576008 201726 576178
rect 200966 575550 201586 575972
rect 201602 575534 201618 575992
rect 201942 575958 201976 576416
rect 202118 576412 205868 576416
rect 202244 576369 205868 576412
rect 202230 576365 205868 576369
rect 206252 576391 206286 576450
rect 206288 576416 206890 576450
rect 206252 576368 206294 576391
rect 202045 576353 202090 576364
rect 202231 576357 205868 576365
rect 206215 576357 206294 576368
rect 202056 575958 202090 576353
rect 201636 575924 202202 575958
rect 201636 575602 201670 575924
rect 201942 575844 201976 575924
rect 202056 575861 202090 575924
rect 202168 575865 202202 575924
rect 202242 575865 205868 576357
rect 202007 575844 202018 575855
rect 201691 575782 201772 575829
rect 201831 575810 202018 575844
rect 201738 575744 201772 575782
rect 201942 575716 201976 575810
rect 202019 575782 202100 575829
rect 202168 575818 205868 575865
rect 202102 575784 205868 575818
rect 202066 575728 202100 575782
rect 202007 575716 202018 575727
rect 202168 575716 202202 575784
rect 202230 575768 205868 575784
rect 202242 575716 205868 575768
rect 201831 575682 205868 575716
rect 202168 575602 202202 575682
rect 201636 575568 202202 575602
rect 202242 575646 205868 575682
rect 201504 575420 201512 575450
rect 201532 575420 201540 575422
rect 201660 575220 201676 575420
rect 201688 575192 201704 575448
rect 202242 575302 203084 575646
rect 203627 575322 205868 575646
rect 206226 576210 206294 576357
rect 206366 576369 206443 576416
rect 206366 576309 206400 576369
rect 206375 576293 206400 576309
rect 206409 576297 206443 576369
rect 206494 576309 206528 576416
rect 206409 576284 206455 576297
rect 206394 576250 206455 576284
rect 206466 576250 206513 576297
rect 206409 576216 206513 576250
rect 206226 576148 206286 576210
rect 206409 576200 206455 576216
rect 206409 576148 206443 576200
rect 206608 576148 206642 576416
rect 206226 576114 206642 576148
rect 206728 576148 206762 576416
rect 206842 576368 206876 576416
rect 206884 576368 206910 576373
rect 206842 576357 206918 576368
rect 206842 576309 206876 576357
rect 206850 576293 206876 576309
rect 206884 576284 206918 576357
rect 206970 576309 207032 576485
rect 206870 576250 206918 576284
rect 206942 576250 206989 576297
rect 206884 576216 206989 576250
rect 206884 576148 206918 576216
rect 206998 576148 207032 576309
rect 207084 576210 207135 576552
rect 207084 576148 207113 576210
rect 207181 576172 207215 576617
rect 207250 576586 207251 576749
rect 209820 576718 209854 577146
rect 209934 576718 209968 576752
rect 210592 576718 210626 576752
rect 210706 576718 210740 577146
rect 211010 576718 211044 577146
rect 211124 576718 211158 576752
rect 211782 576718 211816 576752
rect 211896 576718 211930 577146
rect 208830 576684 212190 576718
rect 209820 576588 209854 576684
rect 210586 576654 210588 576658
rect 209922 576588 210174 576654
rect 210188 576616 210638 576654
rect 210226 576588 210638 576616
rect 210706 576588 210740 576684
rect 211010 576588 211044 576684
rect 211112 576588 211490 576654
rect 211504 576616 211828 576654
rect 211542 576588 211828 576616
rect 211896 576588 211930 576684
rect 212320 576588 212340 576772
rect 213206 576588 213240 576606
rect 207504 576172 207505 576586
rect 208698 576172 209154 576586
rect 209608 576584 213240 576588
rect 209428 576576 209490 576584
rect 209556 576576 213240 576584
rect 207158 576148 209154 576172
rect 206728 576114 207113 576148
rect 206226 576064 206260 576114
rect 206409 576064 206443 576114
rect 206884 576064 206918 576114
rect 206998 576064 207032 576114
rect 206226 576012 206656 576064
rect 206710 576012 207132 576064
rect 206226 575866 207132 576012
rect 206226 575444 206656 575866
rect 206710 575444 207132 575866
rect 206226 575381 206271 575444
rect 206409 575369 206504 575444
rect 206884 575381 206929 575444
rect 205886 575322 206903 575369
rect 203627 575302 206245 575322
rect 202242 575152 202276 575302
rect 205454 575220 205488 575302
rect 205630 575288 206245 575302
rect 206288 575288 206903 575322
rect 205739 575272 205797 575288
rect 206397 575272 206455 575288
rect 206952 575220 206984 575230
rect 206998 575220 207032 575444
rect 205454 575186 207032 575220
rect 202278 575152 202310 575184
rect 197356 575148 199006 575152
rect 190736 574480 193018 574876
rect 193526 574710 194752 574744
rect 196318 574740 196332 574768
rect 187838 574446 193018 574480
rect 177610 574344 182738 574378
rect 173858 574034 176629 574070
rect 178112 574034 178146 574344
rect 178226 574034 178260 574068
rect 178884 574034 178918 574068
rect 179542 574034 179576 574068
rect 180200 574034 180234 574068
rect 180858 574034 180892 574068
rect 181516 574034 181550 574068
rect 181630 574034 181664 574344
rect 190736 574308 193018 574446
rect 186926 574056 186960 574068
rect 187084 574062 187118 574081
rect 194122 574070 194156 574651
rect 196318 574448 196332 574638
rect 196318 574440 196342 574448
rect 196306 574438 196342 574440
rect 196318 574406 196342 574438
rect 196280 574404 196342 574406
rect 196318 574374 196342 574404
rect 187242 574056 187276 574068
rect 190736 574034 193044 574070
rect 173858 574000 193044 574034
rect 173858 573348 176629 574000
rect 178112 573920 178146 574000
rect 178226 573920 178260 574000
rect 178884 573920 178918 574000
rect 179542 573920 179576 574000
rect 180200 573920 180234 574000
rect 180858 573920 180892 574000
rect 181516 573920 181550 574000
rect 181630 573920 181664 574000
rect 186926 573960 187276 573986
rect 184194 573938 184242 573954
rect 178112 573886 181664 573920
rect 178112 573462 178146 573886
rect 178226 573462 178260 573886
rect 178272 573874 178273 573875
rect 178871 573874 178872 573875
rect 178271 573873 178272 573874
rect 178872 573873 178873 573874
rect 178271 573474 178272 573475
rect 178872 573474 178873 573475
rect 178272 573473 178273 573474
rect 178871 573473 178872 573474
rect 178884 573462 178918 573886
rect 178930 573874 178931 573875
rect 179529 573874 179530 573875
rect 178929 573873 178930 573874
rect 179530 573873 179531 573874
rect 178929 573474 178930 573475
rect 179530 573474 179531 573475
rect 178930 573473 178931 573474
rect 179529 573473 179530 573474
rect 179542 573462 179576 573886
rect 179588 573874 179589 573875
rect 180187 573874 180188 573875
rect 179587 573873 179588 573874
rect 180188 573873 180189 573874
rect 179587 573474 179588 573475
rect 180188 573474 180189 573475
rect 179588 573473 179589 573474
rect 180187 573473 180188 573474
rect 180200 573462 180234 573886
rect 180246 573874 180247 573875
rect 180845 573874 180846 573875
rect 180245 573873 180246 573874
rect 180846 573873 180847 573874
rect 180245 573474 180246 573475
rect 180846 573474 180847 573475
rect 180246 573473 180247 573474
rect 180845 573473 180846 573474
rect 180858 573462 180892 573886
rect 180904 573874 180905 573875
rect 181503 573874 181504 573875
rect 180903 573873 180904 573874
rect 181504 573873 181505 573874
rect 180903 573474 180904 573475
rect 181504 573474 181505 573475
rect 180904 573473 180905 573474
rect 181503 573473 181504 573474
rect 181516 573462 181550 573886
rect 181630 573462 181664 573886
rect 184042 573905 184068 573932
rect 184194 573920 184208 573938
rect 184216 573920 184242 573932
rect 190736 573920 193044 574000
rect 184072 573905 184076 573908
rect 182158 573490 182742 573504
rect 178112 573428 181664 573462
rect 184042 573463 184076 573905
rect 184208 573905 184212 573908
rect 184216 573905 193044 573920
rect 184208 573886 193044 573905
rect 184106 573870 184140 573874
rect 184100 573790 184140 573870
rect 184106 573474 184140 573790
rect 184144 573474 184178 573874
rect 184208 573496 184242 573886
rect 184042 573440 184068 573463
rect 184072 573440 184076 573463
rect 184194 573463 184242 573496
rect 184194 573462 184212 573463
rect 184208 573440 184212 573462
rect 184216 573462 184242 573463
rect 183954 573428 184068 573440
rect 178112 573348 178146 573428
rect 178226 573348 178260 573428
rect 178884 573348 178918 573428
rect 179542 573348 179576 573428
rect 180200 573348 180234 573428
rect 180858 573348 180892 573428
rect 181516 573348 181550 573428
rect 181630 573348 181664 573428
rect 184042 573416 184068 573428
rect 184216 573428 184262 573462
rect 190736 573438 193044 573886
rect 193314 573444 194426 574070
rect 194746 573664 194774 573782
rect 184216 573416 184242 573428
rect 183988 573394 184042 573406
rect 173858 573314 194294 573348
rect 173858 573278 176629 573314
rect 178112 573182 178146 573314
rect 181630 573182 181664 573314
rect 197384 573274 197418 575020
rect 199460 574876 203084 575152
rect 203627 574882 205768 575152
rect 197860 573714 199262 573728
rect 199460 573438 203192 574876
rect 203462 574758 205768 574882
rect 203462 574430 205785 574758
rect 205792 574468 205823 574720
rect 203462 573444 205768 574430
rect 206409 574059 206443 574093
rect 206952 574059 206984 575186
rect 207008 574059 207012 575186
rect 207067 574059 207101 574093
rect 207181 574059 207215 576148
rect 207504 575148 207505 576148
rect 208698 575895 209154 576148
rect 209608 575920 213240 576576
rect 213632 576528 213642 577140
rect 216078 577100 216098 577134
rect 215612 577066 216160 577100
rect 215612 576784 215646 577066
rect 216092 577004 216112 577038
rect 215787 576986 215985 576997
rect 215992 576992 216006 577000
rect 215676 576942 215786 576980
rect 215798 576952 215985 576986
rect 215988 576980 216006 576992
rect 215986 576942 216096 576980
rect 215714 576908 215786 576942
rect 215787 576898 215985 576909
rect 215798 576864 215985 576898
rect 215988 576860 216006 576942
rect 216016 576908 216096 576942
rect 216016 576888 216034 576908
rect 216066 576892 216074 576908
rect 216020 576866 216034 576888
rect 216078 576870 216096 576908
rect 215992 576838 216006 576860
rect 216078 576784 216098 576818
rect 216114 576784 216118 576790
rect 216126 576784 216160 577066
rect 215612 576750 216160 576784
rect 216210 576749 216848 577154
rect 213775 576611 214444 576749
rect 214612 576611 217875 576749
rect 213775 576577 217875 576611
rect 209608 575918 213232 575920
rect 209608 575895 213240 575918
rect 208312 575859 208346 575893
rect 208698 575886 213240 575895
rect 213488 575912 213522 575918
rect 213775 575912 214444 576577
rect 214490 576536 214518 576577
rect 214462 576528 214490 576536
rect 214518 576528 214546 576536
rect 214612 576529 217875 576577
rect 214490 576480 214518 576528
rect 214572 576518 217875 576529
rect 218046 576528 218048 576630
rect 213488 575900 214444 575912
rect 214583 575908 217875 576518
rect 218166 575970 218200 577538
rect 218166 575908 218200 575913
rect 214583 575900 218200 575908
rect 213488 575895 218200 575900
rect 208698 575864 213232 575886
rect 213488 575878 218236 575895
rect 213775 575864 218236 575878
rect 208698 575859 218236 575864
rect 218520 575859 218554 576866
rect 219286 576754 219300 576779
rect 218846 576718 222108 576754
rect 228994 576718 230367 576749
rect 218846 576684 222814 576718
rect 228994 576713 235306 576718
rect 224055 576684 235306 576713
rect 218846 576616 222108 576684
rect 224055 576679 230367 576684
rect 222230 576622 222258 576648
rect 222400 576632 222411 576643
rect 222423 576632 222434 576643
rect 222400 576616 222434 576632
rect 218846 576582 222434 576616
rect 218846 576543 222108 576582
rect 222202 576576 222230 576582
rect 218846 575895 222149 576543
rect 222230 576528 222258 576576
rect 222275 576532 222331 576543
rect 218634 575859 218668 575893
rect 218846 575864 222225 575895
rect 222286 575864 222331 576532
rect 222400 575864 222434 576582
rect 222678 576576 222746 576584
rect 222762 575864 222796 575898
rect 222876 575864 222910 576622
rect 226779 576611 226813 576649
rect 227477 576627 227488 576638
rect 227500 576627 227511 576638
rect 227477 576611 227511 576627
rect 224123 576571 224190 576584
rect 224638 576571 224715 576584
rect 224781 576571 224848 576584
rect 225296 576571 225373 576584
rect 226779 576577 227511 576611
rect 226779 575900 226813 576577
rect 226882 576518 226927 576529
rect 227352 576518 227397 576529
rect 226893 575900 226927 576518
rect 223923 575864 227296 575900
rect 218846 575859 227296 575864
rect 208013 575850 227296 575859
rect 208013 575825 212322 575850
rect 208013 575218 208047 575825
rect 208489 575804 208523 575825
rect 208698 575804 212322 575825
rect 208142 575757 212322 575804
rect 208189 575723 212322 575757
rect 208300 575676 208358 575723
rect 208116 575664 208172 575675
rect 208127 575367 208172 575664
rect 208312 575379 208357 575676
rect 208489 575367 208523 575723
rect 208592 575664 208648 575675
rect 208698 575664 212322 575723
rect 213048 575830 227296 575850
rect 213048 575704 213232 575830
rect 213775 575825 222225 575830
rect 213560 575762 213594 575809
rect 213775 575804 217148 575825
rect 217215 575804 217260 575825
rect 217329 575804 217363 575825
rect 213775 575762 217737 575804
rect 213560 575757 217737 575762
rect 213560 575728 217560 575757
rect 213560 575704 213594 575728
rect 213775 575723 217560 575728
rect 217603 575723 217737 575757
rect 213775 575704 217148 575723
rect 213048 575668 217148 575704
rect 208603 575408 212322 575664
rect 208603 575367 208648 575408
rect 208698 575367 212322 575408
rect 208115 575320 212322 575367
rect 208115 575286 208331 575320
rect 208374 575286 212322 575320
rect 208115 575270 208173 575286
rect 208115 575255 208130 575270
rect 208244 575218 208252 575280
rect 208489 575218 208523 575286
rect 208603 575218 208648 575286
rect 208664 575218 208692 575280
rect 208698 575218 212322 575286
rect 207636 575184 212322 575218
rect 208013 574059 208047 575184
rect 208244 574059 208252 575184
rect 208489 574059 208523 575184
rect 208603 574059 208648 575184
rect 208664 574059 208692 575184
rect 208698 574100 212322 575184
rect 212374 575634 217148 575668
rect 212374 575340 212408 575634
rect 213048 575582 217148 575634
rect 213036 575566 217148 575582
rect 212550 575532 217148 575566
rect 213036 575485 217148 575532
rect 212477 575473 212522 575484
rect 212374 575126 212430 575340
rect 212452 575182 212458 575340
rect 212374 574336 212408 575126
rect 212426 574858 212430 575126
rect 212426 574658 212432 574858
rect 212426 574429 212430 574658
rect 212488 574497 212522 575473
rect 212628 574948 212820 575000
rect 213048 574948 217148 575485
rect 212604 574880 217148 574948
rect 213048 574485 217148 574880
rect 213036 574438 217148 574485
rect 212550 574404 217148 574438
rect 213036 574388 217148 574404
rect 213048 574336 217148 574388
rect 212374 574302 217148 574336
rect 212384 574100 212388 574302
rect 213048 574266 217148 574302
rect 213048 574100 213232 574266
rect 208698 574064 213232 574100
rect 213560 574064 213594 574266
rect 213674 574064 213719 574266
rect 213750 574064 217148 574266
rect 208698 574059 217148 574064
rect 217215 574059 217260 575723
rect 217329 574059 217363 575723
rect 217679 575676 217737 575723
rect 217530 575664 217586 575675
rect 217541 574059 217586 575664
rect 217620 574820 217626 575340
rect 217648 574848 217682 575340
rect 217658 574059 217682 574848
rect 217691 574059 217736 575676
rect 217805 574059 217839 575825
rect 218520 575757 218554 575825
rect 218637 575804 218671 575825
rect 218846 575804 222225 575825
rect 218622 575800 222225 575804
rect 222286 575800 222331 575830
rect 222400 575800 222434 575830
rect 218622 575797 222622 575800
rect 218603 575763 222622 575797
rect 218622 575757 222622 575763
rect 222636 575762 222808 575800
rect 218261 575728 222622 575757
rect 222674 575728 222808 575762
rect 218261 575723 222225 575728
rect 218199 574059 218233 574093
rect 218520 574059 218554 575723
rect 218622 575676 218702 575723
rect 218634 574059 218702 575676
rect 218740 575664 218796 575675
rect 218751 574059 218796 575664
rect 218846 574064 222225 575723
rect 222286 574064 222331 575728
rect 222400 574064 222434 575728
rect 222750 575690 222808 575728
rect 222601 575678 222657 575689
rect 222612 574064 222657 575678
rect 222714 575170 222734 575340
rect 222686 574820 222704 575114
rect 222714 574848 222760 575170
rect 222738 574064 222760 574848
rect 222762 574064 222807 575690
rect 222876 574064 222910 575830
rect 223708 575762 223742 575809
rect 223923 575762 227296 575830
rect 223708 575728 227296 575762
rect 223270 574064 223304 574098
rect 223708 574064 223742 575728
rect 223923 575689 227296 575728
rect 223811 575678 223856 575689
rect 223917 575678 227296 575689
rect 223822 575152 223856 575678
rect 223822 574064 223862 575152
rect 223888 574064 223890 575096
rect 223923 574064 227296 575678
rect 218846 574059 227296 574064
rect 195720 573240 199176 573274
rect 174471 572996 174505 573182
rect 175129 572996 175163 573182
rect 197384 573172 197418 573240
rect 197486 573172 197520 573182
rect 197684 573172 197722 573210
rect 198342 573172 198380 573210
rect 199000 573172 199038 573210
rect 197384 573138 197722 573172
rect 197774 573138 198380 573172
rect 198432 573138 199038 573172
rect 195732 573094 195778 573100
rect 195732 573088 195804 573094
rect 195738 573076 195804 573088
rect 173748 571420 175230 572996
rect 195772 572688 195804 573076
rect 195772 571584 195778 572688
rect 195828 572660 195832 573122
rect 197048 573088 197094 573100
rect 197048 573076 197088 573088
rect 196456 571640 196470 571886
rect 196484 571584 196526 571886
rect 197048 571840 197072 572748
rect 197384 571598 197418 573138
rect 197486 573056 197520 573138
rect 197678 573112 197780 573128
rect 198336 573122 198438 573128
rect 198306 573112 198464 573122
rect 198994 573112 199096 573128
rect 197558 573100 197559 573101
rect 197557 573099 197558 573100
rect 197706 573099 197752 573100
rect 198364 573099 198410 573100
rect 199022 573099 199068 573100
rect 197701 573088 197752 573099
rect 198359 573094 198410 573099
rect 197706 573084 197752 573088
rect 198334 573084 198436 573094
rect 199017 573088 199068 573099
rect 199022 573084 199068 573088
rect 197700 573040 197701 573041
rect 197699 573039 197700 573040
rect 197712 573028 197746 573084
rect 197757 573040 197758 573041
rect 198358 573040 198359 573041
rect 197758 573039 197759 573040
rect 198357 573039 198358 573040
rect 198370 573028 198404 573084
rect 198415 573040 198416 573041
rect 199016 573040 199017 573041
rect 198416 573039 198417 573040
rect 199015 573039 199016 573040
rect 199028 573028 199062 573084
rect 199142 573028 199176 573240
rect 197448 572966 197520 573004
rect 197570 572994 199176 573028
rect 197699 572982 197700 572983
rect 197700 572981 197701 572982
rect 197486 572398 197520 572966
rect 197700 572382 197701 572383
rect 197699 572381 197700 572382
rect 197712 572370 197746 572994
rect 197758 572982 197759 572983
rect 198357 572982 198358 572983
rect 197757 572981 197758 572982
rect 198358 572981 198359 572982
rect 197757 572382 197758 572383
rect 198358 572382 198359 572383
rect 197758 572381 197759 572382
rect 198357 572381 198358 572382
rect 198370 572370 198404 572994
rect 198416 572982 198417 572983
rect 199015 572982 199016 572983
rect 198415 572981 198416 572982
rect 199016 572981 199017 572982
rect 198415 572382 198416 572383
rect 199016 572382 199017 572383
rect 198416 572381 198417 572382
rect 199015 572381 199016 572382
rect 199028 572370 199062 572994
rect 199142 572370 199176 572994
rect 197448 572308 197520 572346
rect 197570 572336 199176 572370
rect 197699 572324 197700 572325
rect 197700 572323 197701 572324
rect 197486 571740 197520 572308
rect 197700 571724 197701 571725
rect 197699 571723 197700 571724
rect 197712 571712 197746 572336
rect 197758 572324 197759 572325
rect 198357 572324 198358 572325
rect 197757 572323 197758 572324
rect 198358 572323 198359 572324
rect 197757 571724 197758 571725
rect 198358 571724 198359 571725
rect 197758 571723 197759 571724
rect 198357 571723 198358 571724
rect 198370 571712 198404 572336
rect 198416 572324 198417 572325
rect 199015 572324 199016 572325
rect 198415 572323 198416 572324
rect 199016 572323 199017 572324
rect 198415 571724 198416 571725
rect 199016 571724 199017 571725
rect 198416 571723 198417 571724
rect 199015 571723 199016 571724
rect 199028 571712 199062 572336
rect 199142 571712 199176 572336
rect 199460 572150 203084 573438
rect 203627 573310 205768 573444
rect 206145 574030 227296 574059
rect 206145 574025 213232 574030
rect 206145 573310 206179 574025
rect 206320 573963 206332 574025
rect 206409 573973 206456 574004
rect 206397 573957 206456 573973
rect 206889 573957 206936 574004
rect 206952 573963 206984 574025
rect 207008 573976 207012 574025
rect 207008 573963 207040 573976
rect 207067 573973 207113 574004
rect 207055 573957 207113 573973
rect 206321 573923 206936 573957
rect 206979 573923 207113 573957
rect 206248 573864 206293 573875
rect 206259 573310 206293 573864
rect 206320 573310 206332 573917
rect 206397 573876 206455 573923
rect 206409 573310 206443 573876
rect 206906 573864 206951 573875
rect 206917 573310 206951 573864
rect 206952 573570 206984 573917
rect 207008 573626 207040 573917
rect 207055 573876 207113 573923
rect 206952 573310 207002 573570
rect 207008 573310 207058 573626
rect 207067 573310 207101 573876
rect 207181 573310 207215 574025
rect 208013 573310 208047 574025
rect 208188 574004 208196 574025
rect 208244 574019 208252 574025
rect 208244 574004 208273 574019
rect 208489 574004 208523 574025
rect 208603 574004 208648 574025
rect 208664 574004 208692 574025
rect 208698 574004 213232 574025
rect 208115 574000 213232 574004
rect 213308 574000 213344 574024
rect 213560 574000 213594 574030
rect 213674 574000 213719 574030
rect 213750 574025 222225 574030
rect 213750 574000 217148 574025
rect 208115 573968 217148 574000
rect 208115 573957 213316 573968
rect 213328 573964 217148 573968
rect 217215 574022 217260 574025
rect 217215 573964 217249 574022
rect 217329 573964 217363 574025
rect 217541 574022 217586 574025
rect 217541 573964 217575 574022
rect 217608 574018 217626 574019
rect 217658 573964 217682 574025
rect 217691 574022 217736 574025
rect 217691 573964 217725 574022
rect 217805 573964 217839 574025
rect 218199 574004 218233 574025
rect 217898 573964 217994 574004
rect 213328 573962 217994 573964
rect 218171 573991 218233 574004
rect 218171 573963 218239 573991
rect 208115 573923 208252 573957
rect 208295 573928 213316 573957
rect 213366 573957 217994 573962
rect 218165 573957 218239 573963
rect 218249 573957 218267 573963
rect 218520 573957 218554 574025
rect 218634 573957 218702 574025
rect 218751 574022 218796 574025
rect 218751 574004 218785 574022
rect 218846 574004 222225 574025
rect 218751 573973 218798 574004
rect 218739 573957 218798 573973
rect 218829 574000 222225 574004
rect 222286 574000 222331 574030
rect 222400 574000 222434 574030
rect 222612 574000 222657 574030
rect 222678 574010 222704 574024
rect 222738 574000 222760 574030
rect 222762 574000 222807 574030
rect 222876 574000 222910 574030
rect 223270 574000 223304 574030
rect 218829 573962 223650 574000
rect 223708 573962 223742 574030
rect 223822 573978 223862 574030
rect 223888 573996 223890 574030
rect 223923 574000 227296 574030
rect 223900 573996 227296 574000
rect 223888 573992 227296 573996
rect 223810 573968 223868 573978
rect 223900 573968 227296 573992
rect 223810 573962 227296 573968
rect 218829 573957 222657 573962
rect 213366 573930 218239 573957
rect 213366 573928 217575 573930
rect 208295 573923 213288 573928
rect 208115 573917 208217 573923
rect 208244 573917 208245 573923
rect 208115 573876 208196 573917
rect 208244 573876 208273 573917
rect 208127 573576 208196 573876
rect 208227 573875 208273 573876
rect 208222 573864 208278 573875
rect 208227 573576 208278 573864
rect 208127 573310 208172 573576
rect 208233 573310 208278 573576
rect 208489 573310 208523 573923
rect 208603 573310 208648 573923
rect 208698 573922 213288 573923
rect 208698 573890 213244 573922
rect 213308 573894 213316 573928
rect 208698 573888 213243 573890
rect 208698 573502 213232 573888
rect 213293 573878 213338 573889
rect 213304 573502 213338 573878
rect 213560 573502 213594 573928
rect 213674 573888 213719 573928
rect 213775 573923 217575 573928
rect 217587 573923 218239 573930
rect 218245 573928 222657 573957
rect 222674 573928 223310 573962
rect 218245 573923 222225 573928
rect 213674 573502 213708 573888
rect 213775 573862 217148 573923
rect 217160 573862 217207 573909
rect 213775 573828 217207 573862
rect 217215 573862 217249 573923
rect 217329 573862 217363 573923
rect 217541 573909 217575 573923
rect 217608 573917 217658 573923
rect 217541 573878 217588 573909
rect 217529 573862 217588 573878
rect 217658 573868 217664 573917
rect 217691 573909 217725 573923
rect 217608 573862 217658 573868
rect 217691 573862 217738 573909
rect 217805 573862 217839 573923
rect 217215 573828 217839 573862
rect 208698 573310 213748 573502
rect 203627 573262 213748 573310
rect 203444 573228 213748 573262
rect 203444 573028 203478 573228
rect 203627 573160 213748 573228
rect 203620 573126 213748 573160
rect 203524 573112 203626 573116
rect 203552 573087 203598 573088
rect 203547 573084 203598 573087
rect 203547 573076 203592 573084
rect 203558 573028 203592 573076
rect 203596 573034 203614 573084
rect 203627 573028 213748 573126
rect 203410 572994 213748 573028
rect 203444 572370 203478 572994
rect 203558 572370 203592 572994
rect 203596 572896 203614 572988
rect 203627 572564 213748 572994
rect 213775 572734 217148 573828
rect 217215 573780 217249 573828
rect 217177 573769 217249 573780
rect 217188 572793 217249 573769
rect 217160 572734 217207 572781
rect 213775 572700 217207 572734
rect 217215 572734 217249 572793
rect 217329 572734 217363 573828
rect 217529 573781 217587 573828
rect 217541 573048 217575 573781
rect 217524 572734 217594 573048
rect 217691 572781 217725 573828
rect 217805 573780 217839 573828
rect 217846 573780 217873 573785
rect 217805 573769 217880 573780
rect 217691 572734 217738 572781
rect 217805 572734 217839 573769
rect 217846 572793 217880 573769
rect 217846 572777 217873 572793
rect 217215 572700 217839 572734
rect 213775 572632 217148 572700
rect 217215 572652 217249 572700
rect 217215 572632 217260 572652
rect 217284 572632 217496 572700
rect 217524 572632 217594 572700
rect 217626 572694 217658 572700
rect 217658 572644 217682 572694
rect 217691 572652 217725 572700
rect 217626 572638 217658 572644
rect 217691 572632 217736 572652
rect 217805 572632 217839 572700
rect 217960 572632 217994 573923
rect 218165 573917 218183 573923
rect 218193 573889 218239 573923
rect 218249 573917 218267 573923
rect 218199 573188 218233 573889
rect 218520 573188 218554 573923
rect 218634 573280 218702 573923
rect 218739 573876 218797 573923
rect 218751 573378 218785 573876
rect 218751 573280 218796 573378
rect 218634 573198 218796 573280
rect 218634 573188 218702 573198
rect 218751 573188 218796 573198
rect 218846 573188 222225 573923
rect 213775 572598 217994 572632
rect 218040 573154 218430 573188
rect 218040 572656 218074 573154
rect 218182 573086 218199 573120
rect 218200 573086 218245 573102
rect 218254 573086 218301 573133
rect 218200 573052 218301 573086
rect 218200 573043 218245 573052
rect 218264 573044 218280 573052
rect 218148 573004 218162 573005
rect 218165 573004 218188 573009
rect 218143 572993 218188 573004
rect 218154 572817 218188 572993
rect 218148 572805 218162 572814
rect 218165 572801 218188 572817
rect 218199 573005 218245 573043
rect 218199 572805 218233 573005
rect 218271 572993 218316 573004
rect 218282 572817 218316 572993
rect 218199 572792 218245 572805
rect 218182 572767 218245 572792
rect 218182 572758 218199 572767
rect 218200 572766 218245 572767
rect 218254 572766 218301 572805
rect 218200 572724 218301 572766
rect 218200 572708 218245 572724
rect 218264 572684 218296 572724
rect 218292 572672 218296 572684
rect 218176 572670 218193 572672
rect 218239 572670 218296 572672
rect 218320 572656 218324 572791
rect 218396 572656 218430 573154
rect 218040 572622 218430 572656
rect 218516 573154 222225 573188
rect 218516 572656 218554 573154
rect 218634 573086 218702 573154
rect 218751 573133 218785 573154
rect 218730 573086 218785 573133
rect 218634 573052 218785 573086
rect 218634 573004 218702 573052
rect 218619 572993 218702 573004
rect 218630 572851 218702 572993
rect 218603 572817 218702 572851
rect 218634 572791 218702 572817
rect 218751 573009 218785 573052
rect 218751 572993 218796 573009
rect 218751 572817 218792 572993
rect 218751 572805 218796 572817
rect 218730 572801 218796 572805
rect 218637 572656 218671 572791
rect 218730 572779 218785 572801
rect 218730 572758 218798 572779
rect 218676 572732 218798 572758
rect 218846 572732 222225 573154
rect 218676 572724 222225 572732
rect 218680 572698 222225 572724
rect 218751 572692 218785 572698
rect 218751 572656 218791 572692
rect 218808 572656 218819 572692
rect 218846 572656 222225 572698
rect 218516 572622 222225 572656
rect 203596 572376 203598 572448
rect 203603 572382 203604 572383
rect 203604 572381 203605 572382
rect 203627 572370 213243 572564
rect 203410 572336 213243 572370
rect 200944 571940 200978 572150
rect 201058 572092 201092 572150
rect 201716 572092 201750 572150
rect 201688 572042 201726 572080
rect 201120 572008 201726 572042
rect 201830 571940 201864 572150
rect 200944 571906 201864 571940
rect 202134 571940 202168 572150
rect 202248 572092 202282 572150
rect 202906 572092 202940 572150
rect 202878 572042 202916 572080
rect 202310 572008 202916 572042
rect 203020 571940 203054 572150
rect 202134 571906 203054 571940
rect 202306 571796 202856 571798
rect 202334 571768 202828 571770
rect 203444 571712 203478 572336
rect 203558 571712 203592 572336
rect 203596 572244 203598 572330
rect 203604 572324 203605 572325
rect 203603 572323 203604 572324
rect 203627 572150 213243 572336
rect 213264 572226 213294 572564
rect 213264 572202 213266 572226
rect 213264 572192 213298 572202
rect 203596 571718 203598 571796
rect 203603 571724 203604 571725
rect 203604 571723 203605 571724
rect 203627 571712 212077 572150
rect 212084 571790 212110 572140
rect 212138 572120 212183 572150
rect 197570 571678 212077 571712
rect 197712 571598 197746 571678
rect 198370 571598 198404 571678
rect 199028 571598 199062 571678
rect 199142 571598 199176 571678
rect 203444 571598 203478 571678
rect 203558 571598 203592 571678
rect 203596 571598 203598 571672
rect 203627 571598 212077 571678
rect 197384 571564 212077 571598
rect 159784 569194 159904 569214
rect 160090 569196 160330 569748
rect 160090 569194 160380 569196
rect 159778 569166 159932 569186
rect 160090 569168 160330 569194
rect 160090 569166 160408 569168
rect 160090 569110 160330 569166
rect 173813 568542 173847 571420
rect 174471 568542 174505 571420
rect 175129 568542 175163 571420
rect 193212 570698 193236 571392
rect 193246 570698 193270 571358
rect 198286 571180 198304 571564
rect 198342 571180 198360 571512
rect 197526 571092 198074 571126
rect 197526 570810 197560 571092
rect 197712 571012 197746 571092
rect 197888 571012 197899 571023
rect 197590 570968 197662 571006
rect 197628 570934 197662 570968
rect 197712 570978 197899 571012
rect 197699 570966 197700 570967
rect 197700 570965 197701 570966
rect 197700 570936 197701 570937
rect 197699 570935 197700 570936
rect 197712 570924 197746 570978
rect 197900 570968 197972 571006
rect 197758 570966 197759 570967
rect 197757 570965 197758 570966
rect 197757 570936 197758 570937
rect 197758 570935 197759 570936
rect 197888 570924 197899 570935
rect 197938 570934 197972 570968
rect 197712 570890 197899 570924
rect 197712 570810 197746 570890
rect 198040 570810 198074 571092
rect 197526 570776 198074 570810
rect 198124 570718 198762 571180
rect 198286 570704 198304 570718
rect 198342 570704 198360 570718
rect 197526 570616 198074 570650
rect 197526 570334 197560 570616
rect 197712 570536 197746 570616
rect 197888 570536 197899 570547
rect 197590 570496 197662 570530
rect 197712 570502 197899 570536
rect 197590 570492 197670 570496
rect 197628 570458 197670 570492
rect 197699 570490 197700 570491
rect 197700 570489 197701 570490
rect 197700 570460 197701 570461
rect 197699 570459 197700 570460
rect 197644 570442 197670 570458
rect 197700 570440 197706 570454
rect 197712 570448 197746 570502
rect 197900 570492 197972 570530
rect 197758 570490 197759 570491
rect 197757 570489 197758 570490
rect 197757 570460 197758 570461
rect 197758 570459 197759 570460
rect 197752 570448 197806 570454
rect 197888 570448 197899 570459
rect 197938 570458 197972 570492
rect 197712 570414 197899 570448
rect 197712 570334 197746 570414
rect 198040 570334 198074 570616
rect 197526 570300 198074 570334
rect 198124 570242 198762 570704
rect 199022 570514 199024 571528
rect 199142 569822 199176 571564
rect 203444 571410 203478 571564
rect 203596 571488 203598 571564
rect 203627 571528 212077 571564
rect 203627 571278 204400 571528
rect 182218 569194 182338 569214
rect 182524 569196 182764 569748
rect 182524 569194 182814 569196
rect 182212 569166 182366 569186
rect 182524 569168 182764 569194
rect 182524 569166 182842 569168
rect 182524 569110 182764 569166
rect 203777 568542 203811 571278
rect 204401 569770 204406 571358
rect 204435 569770 204440 571392
rect 204576 571286 205568 571528
rect 205093 568542 205127 571286
rect 205736 569690 212077 571528
rect 212084 571316 212110 571604
rect 206145 568381 206179 569690
rect 206259 569258 206304 569690
rect 206259 568530 206293 569258
rect 206316 568776 206332 569690
rect 206247 568483 206306 568530
rect 206320 568489 206332 568776
rect 206409 569258 206454 569690
rect 206478 569618 206690 569690
rect 206917 569258 206962 569690
rect 206978 569306 206984 569566
rect 206409 568542 206443 569258
rect 206917 568530 206951 569258
rect 207034 568530 207040 569566
rect 207067 569258 207112 569690
rect 207067 568542 207101 569258
rect 206381 568483 206428 568530
rect 206905 568483 206964 568530
rect 207034 568489 207086 568530
rect 207039 568483 207086 568489
rect 206247 568449 206428 568483
rect 206471 568449 207086 568483
rect 206247 568433 206305 568449
rect 206320 568436 206332 568443
rect 206905 568433 206963 568449
rect 206247 568418 206262 568433
rect 207034 568381 207040 568443
rect 207181 568381 207215 569690
rect 207364 569658 207366 569670
rect 207376 569610 207378 569658
rect 203759 568347 207215 568381
rect 159784 566540 159904 566560
rect 160090 566542 160330 567094
rect 160090 566540 160380 566542
rect 159778 566512 159932 566532
rect 160090 566514 160330 566540
rect 160090 566512 160408 566514
rect 160090 566456 160330 566512
rect 206145 565789 206179 568347
rect 207575 567338 207609 569690
rect 208013 567527 208047 569690
rect 208127 569414 208172 569690
rect 208127 569258 208202 569414
rect 208127 567688 208161 569258
rect 208171 568058 208202 569258
rect 208167 568012 208202 568058
rect 208227 568002 208230 569442
rect 208167 567984 208230 568002
rect 208233 569258 208278 569690
rect 208233 567676 208267 569258
rect 208489 567676 208523 569690
rect 208603 569258 208648 569690
rect 208603 567688 208637 569258
rect 208698 568506 212077 569690
rect 212138 568556 212172 572120
rect 212206 571732 212668 572150
rect 212682 571732 213144 572150
rect 213198 572146 213243 572150
rect 213198 572136 213298 572146
rect 213198 572120 213243 572136
rect 213304 572120 213349 572564
rect 213354 572344 213376 572426
rect 213198 571864 213232 572120
rect 212252 571682 212286 571732
rect 212252 571648 212614 571682
rect 212252 571168 212298 571648
rect 212456 571580 212494 571618
rect 212422 571546 212494 571580
rect 212367 571496 212412 571507
rect 212455 571496 212500 571507
rect 212378 571320 212412 571496
rect 212466 571320 212500 571496
rect 212456 571270 212494 571308
rect 212422 571236 212494 571270
rect 212580 571168 212614 571648
rect 212646 571174 212648 571716
rect 213084 571682 213118 571732
rect 212740 571648 213118 571682
rect 212252 571134 212614 571168
rect 212740 571168 212774 571648
rect 212932 571580 212970 571618
rect 212898 571546 212970 571580
rect 212843 571496 212888 571507
rect 212931 571496 212976 571507
rect 212854 571320 212888 571496
rect 212942 571320 212976 571496
rect 212932 571270 212970 571308
rect 212898 571236 212970 571270
rect 213056 571168 213118 571648
rect 212740 571134 213118 571168
rect 212110 568506 212148 568544
rect 208698 568472 212148 568506
rect 208698 568404 212077 568472
rect 212252 568404 212286 571134
rect 213084 569748 213118 571134
rect 213198 571552 213238 571864
rect 213256 571750 213266 571808
rect 213254 571664 213266 571750
rect 213256 571608 213266 571664
rect 213198 571174 213232 571552
rect 213292 571534 213298 571560
rect 213236 571504 213238 571534
rect 213236 571478 213298 571504
rect 213304 571174 213338 572120
rect 213198 570956 213243 571174
rect 213304 571102 213349 571174
rect 213304 571016 213418 571102
rect 213304 570956 213349 571016
rect 213198 570900 213238 570956
rect 213198 569902 213232 570900
rect 213304 569902 213338 570956
rect 213198 569748 213243 569902
rect 213304 569748 213349 569902
rect 213560 569748 213594 572564
rect 213674 572120 213719 572564
rect 212670 569110 213132 569748
rect 213146 569110 213608 569748
rect 212724 569026 213074 569060
rect 212724 568546 212758 569026
rect 212916 568958 212954 568996
rect 212882 568924 212954 568958
rect 212827 568874 212872 568885
rect 212915 568874 212960 568885
rect 212838 568698 212872 568874
rect 212926 568698 212960 568874
rect 212916 568648 212954 568686
rect 212882 568614 212954 568648
rect 213040 568546 213074 569026
rect 212724 568512 213074 568546
rect 208698 568370 212286 568404
rect 208698 568334 212077 568370
rect 208785 567688 208830 568334
rect 208891 567676 208936 568334
rect 209261 567688 209306 568334
rect 209443 567688 209488 568334
rect 209549 567676 209594 568334
rect 208221 567629 208280 567676
rect 208489 567629 208536 567676
rect 208732 567629 209595 567676
rect 209663 567629 209697 568334
rect 209919 567688 209964 568334
rect 209984 568002 210012 568334
rect 210040 568002 210068 568334
rect 210101 567688 210146 568334
rect 210577 567688 210622 568334
rect 210654 568002 210682 568334
rect 210710 568002 210738 568334
rect 210759 567688 210804 568334
rect 211180 567629 212077 568334
rect 208189 567595 212077 567629
rect 208221 567579 208279 567595
rect 208233 567527 208267 567561
rect 208489 567527 208523 567595
rect 208879 567579 208937 567595
rect 209537 567579 209595 567595
rect 209549 567564 209595 567579
rect 208891 567527 208925 567561
rect 209549 567527 209583 567564
rect 209663 567527 209697 567595
rect 211180 567527 212077 567595
rect 208013 567493 212077 567527
rect 213084 567550 213118 569110
rect 213198 569060 213232 569110
rect 213304 569060 213338 569110
rect 213198 569026 213550 569060
rect 213198 568982 213243 569026
rect 213198 568964 213270 568982
rect 213198 568608 213234 568964
rect 213242 568882 213270 568964
rect 213304 568890 213338 569026
rect 213392 568958 213430 568996
rect 213342 568924 213430 568958
rect 213304 568874 213349 568890
rect 213391 568874 213436 568885
rect 213304 568698 213348 568874
rect 213402 568698 213436 568874
rect 213242 568608 213270 568688
rect 213198 568546 213270 568608
rect 213304 568682 213349 568698
rect 213304 568552 213338 568682
rect 213392 568648 213430 568686
rect 213342 568614 213430 568648
rect 213516 568552 213550 569026
rect 213304 568546 213349 568552
rect 213516 568546 213554 568552
rect 213198 568512 213554 568546
rect 213198 568334 213270 568512
rect 213198 567714 213232 568334
rect 213242 567986 213270 568334
rect 213304 568334 213349 568512
rect 213526 568334 213554 568512
rect 213198 567702 213238 567714
rect 213192 567690 213238 567702
rect 213304 567690 213338 568334
rect 213560 567690 213594 569110
rect 213674 567702 213708 572120
rect 213775 568858 217148 572598
rect 217215 572120 217260 572598
rect 217284 572592 217594 572598
rect 217284 572488 217586 572592
rect 217284 572264 217496 572488
rect 217215 569048 217249 572120
rect 217215 568858 217260 569048
rect 217329 568858 217363 572264
rect 217541 572120 217586 572488
rect 217658 572162 217682 572458
rect 217541 569048 217575 572120
rect 217541 568858 217586 569048
rect 217596 568858 217608 569076
rect 217658 569048 217664 572162
rect 217624 568858 217664 569048
rect 217691 572120 217736 572598
rect 217691 569048 217725 572120
rect 217691 568858 217736 569048
rect 217805 568858 217839 572598
rect 218520 572596 222225 572622
rect 218637 572572 218671 572596
rect 218751 572572 218796 572596
rect 218808 572572 218819 572596
rect 218846 572572 222225 572596
rect 218026 571952 218448 572572
rect 218502 571952 222225 572572
rect 218637 571006 218671 571952
rect 218713 571870 218740 571952
rect 218751 571810 218798 571952
rect 218846 571838 222225 571952
rect 222286 572084 222331 573928
rect 222286 571838 222320 572084
rect 222400 571838 222434 573928
rect 218751 571006 218785 571810
rect 218846 571390 222434 571838
rect 218846 571006 222225 571390
rect 218046 570980 222225 571006
rect 218637 570950 218671 570980
rect 218751 570950 218785 570980
rect 218846 570950 222225 570980
rect 217990 570924 222225 570950
rect 218130 569408 218193 569430
rect 218239 569408 218266 569430
rect 218158 569380 218193 569402
rect 218239 569380 218266 569402
rect 218178 568858 218252 569058
rect 213775 568824 217446 568858
rect 213775 568483 217148 568824
rect 217215 568790 217249 568824
rect 217198 568756 217249 568790
rect 217270 568756 217317 568803
rect 217215 568722 217317 568756
rect 217181 568674 217204 568679
rect 217159 568663 217204 568674
rect 217170 568483 217204 568663
rect 217215 568542 217249 568722
rect 217329 568674 217363 568824
rect 217287 568663 217363 568674
rect 217215 568526 217238 568542
rect 217298 568483 217363 568663
rect 217412 568530 217446 568824
rect 217532 568824 217922 568858
rect 217532 568530 217575 568824
rect 217596 568670 217608 568824
rect 217624 568679 217664 568824
rect 217691 568790 217725 568824
rect 217674 568756 217725 568790
rect 217746 568756 217793 568803
rect 217691 568722 217793 568756
rect 217624 568670 217680 568679
rect 217635 568663 217680 568670
rect 217646 568530 217680 568663
rect 217691 568542 217725 568722
rect 217805 568674 217839 568824
rect 217763 568663 217839 568674
rect 217691 568530 217714 568542
rect 217412 568483 217459 568530
rect 217529 568483 217587 568530
rect 217646 568526 217714 568530
rect 217646 568483 217710 568526
rect 217774 568487 217839 568663
rect 213775 568449 217710 568483
rect 213775 568381 217148 568449
rect 217270 568428 217317 568449
rect 217216 568394 217317 568428
rect 217329 568381 217363 568449
rect 217412 568381 217446 568449
rect 217529 568433 217587 568449
rect 217532 568381 217566 568433
rect 217658 568381 217664 568443
rect 217746 568428 217793 568475
rect 217692 568394 217793 568428
rect 217805 568381 217839 568487
rect 213775 568347 217839 568381
rect 213775 568326 217148 568347
rect 217412 568326 217446 568347
rect 213775 568311 217446 568326
rect 213856 567702 213890 568311
rect 213962 567690 213996 568311
rect 214332 567702 214366 568311
rect 214514 567702 214548 568311
rect 214620 567690 214654 568311
rect 213192 567658 213220 567690
rect 213292 567652 213350 567690
rect 213560 567652 213598 567690
rect 213950 567652 214008 567690
rect 214608 567652 214666 567690
rect 213260 567618 214666 567652
rect 213192 567556 213220 567612
rect 213292 567602 213350 567618
rect 213304 567550 213338 567584
rect 213560 567550 213594 567618
rect 213950 567602 214008 567618
rect 214608 567602 214666 567618
rect 214620 567587 214666 567602
rect 214734 567652 214768 568311
rect 214990 567702 215024 568311
rect 215060 568002 215088 568311
rect 215116 568002 215144 568311
rect 215172 567702 215206 568311
rect 215648 567702 215682 568311
rect 215724 568002 215752 568311
rect 215780 568002 215808 568311
rect 215830 567702 215864 568311
rect 216306 567702 216340 568311
rect 216376 568002 216404 568311
rect 216432 568002 216460 568311
rect 216488 567702 216522 568311
rect 216602 567652 216636 568311
rect 216733 568292 217446 568311
rect 217532 568326 217566 568347
rect 217888 568326 217922 568824
rect 217532 568292 217922 568326
rect 218008 568824 218398 568858
rect 218008 568326 218042 568824
rect 218088 568670 218106 568703
rect 218178 568679 218252 568824
rect 218178 568675 218267 568679
rect 218116 568674 218134 568675
rect 218178 568674 218280 568675
rect 218111 568663 218156 568674
rect 218122 568487 218156 568663
rect 218178 568487 218284 568674
rect 218178 568475 218280 568487
rect 218130 568474 218156 568475
rect 218158 568471 218267 568475
rect 218158 568446 218252 568471
rect 218178 568418 218252 568446
rect 218158 568404 218252 568418
rect 218158 568354 218248 568404
rect 218142 568340 218158 568342
rect 218199 568326 218233 568354
rect 218364 568326 218398 568824
rect 218008 568292 218398 568326
rect 216733 568242 217148 568292
rect 216733 567676 217460 568242
rect 217514 567676 217936 568242
rect 217990 567676 218412 568242
rect 216733 567652 218412 567676
rect 214734 567629 218412 567652
rect 218637 567676 218671 570924
rect 218751 567688 218785 570924
rect 218795 568404 218826 569414
rect 218823 568320 218826 568404
rect 218846 568506 222225 570924
rect 222286 568556 222320 571390
rect 222400 568506 222434 571390
rect 222612 572084 222657 573928
rect 222738 572154 222760 573370
rect 222612 569902 222646 572084
rect 222708 571790 222734 572140
rect 222762 572084 222807 573928
rect 222876 572370 222910 573928
rect 223236 573922 223254 573928
rect 223264 573894 223310 573928
rect 223320 573928 227296 573962
rect 223320 573922 223338 573928
rect 223270 572370 223304 573894
rect 222708 571316 222734 571604
rect 222762 569902 222796 572084
rect 222830 571732 223304 572370
rect 222864 571682 223076 571732
rect 222864 571648 223238 571682
rect 222864 571612 223076 571648
rect 223080 571612 223118 571618
rect 222864 571546 223118 571612
rect 222864 571386 223076 571546
rect 223079 571496 223124 571507
rect 222876 571168 222922 571386
rect 223002 571320 223036 571386
rect 223090 571320 223124 571496
rect 223080 571270 223118 571308
rect 223046 571236 223118 571270
rect 223204 571168 223238 571648
rect 222876 571134 223238 571168
rect 222574 569722 222608 569804
rect 222612 569680 222657 569902
rect 222762 569680 222807 569902
rect 222876 569748 222910 571134
rect 223270 569748 223304 571732
rect 223512 571690 223514 571778
rect 223708 569748 223742 573928
rect 223810 573922 223912 573928
rect 223810 573890 223868 573922
rect 223922 573894 227296 573928
rect 223822 573352 223856 573890
rect 223822 572136 223862 573352
rect 223888 572192 223890 573296
rect 223923 572720 227296 573894
rect 223923 572272 227324 572720
rect 223822 569902 223856 572136
rect 223860 571734 223862 571790
rect 223860 571478 223862 571534
rect 223860 571334 223862 571390
rect 223860 571078 223862 571134
rect 223822 569748 223867 569902
rect 223923 569748 227296 572272
rect 222612 568552 222646 569680
rect 222762 569242 222796 569680
rect 222738 569186 222796 569242
rect 222762 569042 222796 569186
rect 222818 569110 223756 569748
rect 223770 569110 227296 569748
rect 222876 569060 222910 569110
rect 223172 569060 223186 569110
rect 222738 568930 222796 569042
rect 222762 568556 222796 568930
rect 222872 569026 223222 569060
rect 222612 568544 222657 568552
rect 222872 568546 222910 569026
rect 223064 568958 223102 568996
rect 223030 568924 223102 568958
rect 222975 568874 223020 568885
rect 223063 568874 223108 568885
rect 223172 568882 223186 569026
rect 222986 568698 223020 568874
rect 223074 568698 223108 568874
rect 223064 568648 223102 568686
rect 223030 568614 223102 568648
rect 223188 568546 223222 569026
rect 222488 568506 222772 568544
rect 222872 568512 223222 568546
rect 218846 568472 222772 568506
rect 218846 568404 222225 568472
rect 222400 568404 222434 568472
rect 222544 568456 222658 568472
rect 222544 568404 222646 568456
rect 222876 568404 222910 568512
rect 218846 568370 222910 568404
rect 218846 568334 222225 568370
rect 218851 568320 218854 568334
rect 218823 568058 218826 568120
rect 218791 568012 218826 568058
rect 218851 568002 218854 568120
rect 218791 567984 218854 568002
rect 218857 567676 218902 568334
rect 219409 567688 219454 568334
rect 219515 567676 219560 568334
rect 219586 567676 219587 567880
rect 220024 567676 220028 567880
rect 220062 567676 220066 567880
rect 220067 567688 220112 568334
rect 220167 568002 220218 568334
rect 220173 567676 220218 568002
rect 218637 567629 218684 567676
rect 218844 567629 220219 567676
rect 220287 567629 220321 568334
rect 221804 567690 222225 568334
rect 222612 568058 222646 568370
rect 222606 567774 222646 568058
rect 222612 567690 222646 567774
rect 223270 567690 223304 569110
rect 223348 569026 223698 569060
rect 223348 568546 223382 569026
rect 223540 568958 223578 568996
rect 223506 568924 223578 568958
rect 223451 568874 223496 568885
rect 223539 568874 223584 568885
rect 223462 568698 223496 568874
rect 223550 568698 223584 568874
rect 223540 568648 223578 568686
rect 223506 568614 223578 568648
rect 223664 568546 223698 569026
rect 223348 568512 223698 568546
rect 221804 567652 222924 567690
rect 223242 567686 223304 567690
rect 223708 567690 223742 569110
rect 223822 569060 223856 569110
rect 223923 569060 227296 569110
rect 223822 569026 227296 569060
rect 223822 568982 223867 569026
rect 223923 568982 227296 569026
rect 223822 568964 223894 568982
rect 223822 568608 223858 568964
rect 223866 568882 223894 568964
rect 223922 568882 227296 568982
rect 223866 568608 223894 568688
rect 223822 568546 223894 568608
rect 223923 568546 227296 568882
rect 223822 568512 227296 568546
rect 227363 569048 227397 576518
rect 227477 576224 227511 576577
rect 228889 576543 228916 576645
rect 228917 576571 228944 576617
rect 227477 574872 227514 576224
rect 227363 568826 227408 569048
rect 227363 568542 227397 568826
rect 223822 568380 223894 568512
rect 223923 568483 227296 568512
rect 227477 568483 227511 574872
rect 228188 573154 228578 573188
rect 228188 572656 228222 573154
rect 228402 573086 228449 573133
rect 228364 573052 228449 573086
rect 228291 572993 228336 573004
rect 228419 572993 228464 573004
rect 228302 572817 228336 572993
rect 228430 572817 228464 572993
rect 228402 572758 228449 572805
rect 228364 572724 228449 572758
rect 228422 572720 228428 572724
rect 228434 572684 228440 572720
rect 228544 572656 228578 573154
rect 228188 572622 228578 572656
rect 228174 571952 228596 572572
rect 228867 571956 228901 576518
rect 228944 574878 228946 576230
rect 228944 572804 228962 573378
rect 228994 572678 230367 576679
rect 231850 576616 231884 576663
rect 232548 576632 232559 576643
rect 232571 576632 232582 576643
rect 232548 576616 232582 576632
rect 231850 576582 232582 576616
rect 231034 575574 231170 575684
rect 231034 575548 231186 575574
rect 231094 575116 231186 575548
rect 230972 572686 231434 573224
rect 228994 572422 230376 572678
rect 230390 572450 230432 572650
rect 230972 572620 231582 572686
rect 230972 572586 231644 572620
rect 231092 572536 231118 572570
rect 231370 572544 231644 572586
rect 231370 572536 231582 572544
rect 231030 572502 231582 572536
rect 228802 571870 228901 571956
rect 228752 571006 228778 571810
rect 228780 571006 228806 571810
rect 228867 571006 228901 571870
rect 228944 571810 228946 572358
rect 228994 571006 230367 572422
rect 231030 572022 231064 572502
rect 231118 572396 231152 572502
rect 231222 572434 231260 572472
rect 231172 572400 231186 572434
rect 231188 572400 231260 572434
rect 231118 572364 231158 572396
rect 231168 572392 231186 572396
rect 231222 572392 231244 572396
rect 231250 572364 231272 572396
rect 231118 572350 231152 572364
rect 231164 572350 231178 572361
rect 231221 572350 231266 572361
rect 231118 572174 231178 572350
rect 231232 572174 231266 572350
rect 231346 572238 231582 572502
rect 231742 572462 231746 572662
rect 231770 572434 231774 572690
rect 231118 572160 231152 572174
rect 231222 572160 231260 572162
rect 231118 572056 231158 572160
rect 231172 572074 231186 572132
rect 231222 572124 231266 572160
rect 231188 572090 231266 572124
rect 231222 572074 231238 572090
rect 231092 572046 231158 572056
rect 231250 572046 231266 572090
rect 231092 572022 231152 572046
rect 231346 572022 231380 572238
rect 231030 571988 231380 572022
rect 231742 571810 231766 572358
rect 231770 572062 231794 572386
rect 231770 571782 231798 572062
rect 231776 571776 231798 571782
rect 231222 571008 231224 571208
rect 228194 570980 230367 571006
rect 231250 570980 231252 571236
rect 228188 569582 228262 569912
rect 228188 569428 228394 569582
rect 228188 569258 228262 569428
rect 228218 568858 228243 568892
rect 223923 568449 227511 568483
rect 223923 568381 227296 568449
rect 227477 568433 227511 568449
rect 227477 568422 227488 568433
rect 227500 568422 227511 568433
rect 227680 568824 228070 568858
rect 227680 568433 227714 568824
rect 227894 568756 227941 568803
rect 227856 568722 227941 568756
rect 227783 568663 227828 568674
rect 227911 568663 227956 568674
rect 227794 568530 227828 568663
rect 227922 568530 227956 568663
rect 227782 568483 227840 568530
rect 227910 568483 227968 568530
rect 227756 568475 227994 568483
rect 227756 568466 227866 568475
rect 227884 568466 227994 568475
rect 227756 568449 227994 568466
rect 227680 568422 227691 568433
rect 227703 568422 227714 568433
rect 228036 568433 228070 568824
rect 228156 568824 228546 568858
rect 228156 568517 228190 568824
rect 228209 568526 228224 568824
rect 228370 568756 228417 568803
rect 228332 568722 228417 568756
rect 228236 568703 228243 568713
rect 228236 568701 228249 568703
rect 228232 568670 228249 568701
rect 228270 568675 228277 568679
rect 228264 568674 228277 568675
rect 228302 568674 228310 568675
rect 228232 568542 228243 568670
rect 228259 568663 228310 568674
rect 228236 568526 228243 568542
rect 228270 568530 228310 568663
rect 228156 568449 228215 568517
rect 228258 568483 228316 568530
rect 228330 568489 228338 568703
rect 228387 568663 228432 568674
rect 228398 568530 228432 568663
rect 228386 568483 228444 568530
rect 228258 568475 228470 568483
rect 228271 568466 228342 568475
rect 228360 568466 228470 568475
rect 228271 568464 228470 568466
rect 228262 568449 228470 568464
rect 227680 568388 227714 568415
rect 227840 568394 227910 568428
rect 228036 568422 228047 568433
rect 228059 568422 228070 568433
rect 228102 568420 228116 568443
rect 228036 568388 228070 568415
rect 228130 568392 228144 568443
rect 228156 568433 228190 568449
rect 228262 568443 228330 568449
rect 228156 568422 228167 568433
rect 228179 568422 228190 568433
rect 228290 568428 228330 568436
rect 228512 568433 228546 568824
rect 228752 568489 228778 570980
rect 228780 568489 228806 570980
rect 228867 568542 228901 570980
rect 228752 568436 228778 568443
rect 228290 568415 228386 568428
rect 228512 568422 228523 568433
rect 228535 568422 228546 568433
rect 228156 568388 228190 568415
rect 228316 568394 228386 568415
rect 228512 568388 228546 568415
rect 228780 568408 228806 568443
rect 228994 568404 230367 570980
rect 230418 568846 230432 570248
rect 231222 569408 231234 569608
rect 231250 569380 231262 569636
rect 231712 568782 231738 570240
rect 231740 568810 231766 570212
rect 231846 568810 231848 570212
rect 231850 568506 231884 576582
rect 231953 576532 231998 576543
rect 232423 576532 232468 576543
rect 231964 568556 231998 576532
rect 232208 572674 232420 572692
rect 232014 572244 232420 572674
rect 232014 572226 232226 572244
rect 232434 568556 232468 576532
rect 232548 575968 232582 576582
rect 232548 574864 232600 575968
rect 278619 575411 278653 580554
rect 280487 577149 280521 583647
rect 280963 583626 280997 583647
rect 281077 583644 281122 583647
rect 281077 583626 281111 583644
rect 280601 583610 280648 583626
rect 280589 583579 280648 583610
rect 280679 583585 280726 583626
rect 280662 583579 280726 583585
rect 280963 583579 281010 583626
rect 281077 583579 281124 583626
rect 281138 583598 281166 583647
rect 281259 583644 281304 583647
rect 281735 583644 281780 583647
rect 281259 583626 281293 583644
rect 281735 583626 281769 583644
rect 281259 583579 281306 583626
rect 281337 583579 281384 583626
rect 281735 583579 281782 583626
rect 281796 583598 281824 583647
rect 281852 583598 281880 583647
rect 281917 583644 281962 583647
rect 281917 583626 281951 583644
rect 281917 583579 281964 583626
rect 281995 583579 282042 583626
rect 280589 583545 280726 583579
rect 280769 583545 281384 583579
rect 281427 583545 282042 583579
rect 280589 583539 280691 583545
rect 280589 583498 280647 583539
rect 280718 583511 280719 583545
rect 280601 583254 280635 583498
rect 280696 583486 280741 583497
rect 280601 581790 280641 583254
rect 280658 581846 280669 583198
rect 280601 577310 280635 581790
rect 280645 577634 280676 579036
rect 280701 577606 280704 579064
rect 280707 577298 280741 583486
rect 280963 577298 280997 583545
rect 281077 577310 281111 583545
rect 281259 577310 281293 583545
rect 281354 583486 281399 583497
rect 281365 581488 281399 583486
rect 281296 581480 281508 581488
rect 281296 581040 281708 581480
rect 281365 577298 281399 581040
rect 281496 581032 281708 581040
rect 281735 577310 281769 583545
rect 281917 577310 281951 583545
rect 282012 583486 282057 583497
rect 282023 581480 282057 583486
rect 282137 581488 282171 583647
rect 282359 583644 282374 584750
rect 282137 581480 282354 581488
rect 281972 581040 282354 581480
rect 281972 581032 282184 581040
rect 282023 577298 282057 581032
rect 280695 577251 280754 577298
rect 280963 577251 281010 577298
rect 281353 577251 281412 577298
rect 282011 577251 282069 577298
rect 280663 577217 282069 577251
rect 280595 577155 280618 577211
rect 280695 577201 280753 577217
rect 280707 577149 280741 577183
rect 280963 577149 280997 577217
rect 281300 577204 281411 577217
rect 281353 577202 281411 577204
rect 281328 577201 281411 577202
rect 282011 577201 282069 577217
rect 281328 577149 281359 577201
rect 282054 577186 282069 577201
rect 282137 577251 282171 581032
rect 282393 577310 282427 585286
rect 282458 579612 282486 584962
rect 282514 579612 282542 584962
rect 282458 577257 282486 579426
rect 282514 577257 282542 579426
rect 282575 577310 282609 585286
rect 282826 581480 282830 581488
rect 282838 581040 282842 581480
rect 283051 580346 283085 585286
rect 283051 580156 283096 580346
rect 283128 580156 283156 584962
rect 283184 580156 283212 584962
rect 283233 580346 283267 585286
rect 283709 583722 283743 585286
rect 283836 583722 283864 584962
rect 283891 583722 283925 585286
rect 284005 583722 284039 585345
rect 283654 583686 284551 583722
rect 285558 583686 285592 585390
rect 286034 585384 286068 585431
rect 287534 585390 287562 585410
rect 287590 585390 287618 585422
rect 288198 585390 288226 585410
rect 288254 585390 288282 585410
rect 288906 585390 288934 585410
rect 289076 585400 289087 585411
rect 289099 585400 289110 585411
rect 289076 585384 289110 585400
rect 286034 585350 289110 585384
rect 286034 583686 286068 585350
rect 286137 585300 286182 585311
rect 286319 585300 286364 585311
rect 286795 585300 286840 585311
rect 286977 585300 287022 585311
rect 287453 585300 287498 585311
rect 286148 583686 286182 585300
rect 286224 583686 286252 584962
rect 286330 583686 286364 585300
rect 286806 583686 286840 585300
rect 286876 583686 286904 584962
rect 286932 583686 286960 584962
rect 286988 583686 287022 585300
rect 283654 583652 287242 583686
rect 283654 581480 284551 583652
rect 285558 581992 285592 583652
rect 286034 583622 286068 583652
rect 286148 583622 286182 583652
rect 285672 583615 285710 583622
rect 285660 583600 285710 583615
rect 285750 583618 285788 583622
rect 285660 583584 285718 583600
rect 285750 583590 285790 583618
rect 285726 583584 285790 583590
rect 286034 583584 286072 583622
rect 286148 583584 286186 583622
rect 286224 583610 286252 583652
rect 286330 583622 286364 583652
rect 286806 583622 286840 583652
rect 286330 583584 286368 583622
rect 286408 583584 286446 583622
rect 286806 583584 286844 583622
rect 286876 583616 286904 583652
rect 286932 583616 286960 583652
rect 286988 583622 287022 583652
rect 286988 583584 287026 583622
rect 287066 583584 287104 583622
rect 285660 583550 285790 583584
rect 285840 583550 286446 583584
rect 286498 583550 287104 583584
rect 285660 583544 285762 583550
rect 285660 583512 285718 583544
rect 285782 583516 285790 583550
rect 285672 582974 285706 583512
rect 285767 583500 285812 583511
rect 285672 582146 285712 582974
rect 283314 581032 284551 581480
rect 284680 581354 285142 581992
rect 285156 581354 285618 581992
rect 285672 581924 285717 582146
rect 285672 581768 285712 581924
rect 285738 581824 285740 582918
rect 285778 582146 285812 583500
rect 285778 581924 285823 582146
rect 285828 581966 285850 582048
rect 285738 581814 285772 581824
rect 285672 581758 285772 581768
rect 285672 581486 285706 581758
rect 283233 580156 283278 580346
rect 282848 580124 283278 580156
rect 282848 580122 283267 580124
rect 282848 579624 282882 580122
rect 283051 580101 283085 580122
rect 283051 580054 283098 580101
rect 283024 580020 283098 580054
rect 283051 579972 283085 580020
rect 283090 579972 283119 579977
rect 282951 579961 282996 579972
rect 282962 579785 282996 579961
rect 283051 579961 283124 579972
rect 283128 579968 283156 580122
rect 283184 579968 283267 580122
rect 283051 579773 283085 579961
rect 283090 579785 283124 579961
rect 283090 579773 283119 579785
rect 283051 579769 283119 579773
rect 283204 579772 283267 579968
rect 283051 579726 283098 579769
rect 283024 579692 283098 579726
rect 283051 579624 283085 579692
rect 283128 579624 283156 579772
rect 283184 579624 283267 579772
rect 282848 579590 283267 579624
rect 283051 579540 283085 579590
rect 283128 579540 283156 579590
rect 283184 579540 283212 579590
rect 283233 579540 283267 579590
rect 282834 578996 283267 579540
rect 282834 578920 283278 578996
rect 283051 578778 283096 578920
rect 283051 577310 283085 578778
rect 283128 577257 283156 578920
rect 283184 577257 283212 578920
rect 283233 578778 283278 578920
rect 283233 577310 283267 578778
rect 283654 577251 284551 581032
rect 284738 581270 285088 581304
rect 284738 580790 284772 581270
rect 284930 581202 284968 581240
rect 284896 581168 284968 581202
rect 284841 581118 284886 581129
rect 284929 581118 284974 581129
rect 284852 580942 284886 581118
rect 284940 580942 284974 581118
rect 284930 580892 284968 580930
rect 284896 580858 284968 580892
rect 285054 580790 285088 581270
rect 285120 580796 285122 581338
rect 285558 581304 285592 581354
rect 285214 581270 285592 581304
rect 284738 580756 285088 580790
rect 285214 580790 285248 581270
rect 285406 581202 285444 581240
rect 285372 581168 285444 581202
rect 285317 581118 285362 581129
rect 285405 581118 285450 581129
rect 285328 580942 285362 581118
rect 285416 580942 285450 581118
rect 285406 580892 285444 580930
rect 285372 580858 285444 580892
rect 285530 580790 285592 581270
rect 285214 580756 285592 580790
rect 282137 577217 284551 577251
rect 281365 577149 281399 577183
rect 282023 577149 282057 577183
rect 282137 577149 282171 577217
rect 282458 577204 282486 577211
rect 282514 577204 282542 577211
rect 283128 577204 283156 577211
rect 283184 577204 283212 577211
rect 283654 577149 284551 577217
rect 280487 577115 284551 577149
rect 285558 577172 285592 580756
rect 285672 581174 285712 581486
rect 285730 581372 285740 581430
rect 285728 581286 285740 581372
rect 285730 581230 285740 581286
rect 285672 580796 285706 581174
rect 285766 581156 285772 581182
rect 285710 581126 285712 581156
rect 285710 581100 285772 581126
rect 285778 580796 285812 581924
rect 285672 580578 285717 580796
rect 285778 580724 285823 580796
rect 285778 580638 285892 580724
rect 285778 580578 285823 580638
rect 285672 580522 285712 580578
rect 285672 577324 285706 580522
rect 285716 577608 285744 579010
rect 285778 577312 285812 580578
rect 286034 577312 286068 583550
rect 286148 577324 286182 583550
rect 286330 577324 286364 583550
rect 286425 583500 286470 583511
rect 286436 581460 286470 583500
rect 286392 581456 286604 581460
rect 286392 581012 286794 581456
rect 286436 577312 286470 581012
rect 286582 581008 286794 581012
rect 286806 577324 286840 583550
rect 286988 577324 287022 583550
rect 287083 583500 287128 583511
rect 287094 581456 287128 583500
rect 287208 581460 287242 583652
rect 287208 581456 287442 581460
rect 287058 581012 287442 581456
rect 287058 581008 287270 581012
rect 287094 577312 287128 581008
rect 285766 577274 285824 577312
rect 286034 577274 286072 577312
rect 286424 577274 286482 577312
rect 287082 577280 287140 577312
rect 287010 577274 287140 577280
rect 287208 577274 287242 581008
rect 287464 577324 287498 585300
rect 287534 577280 287562 585344
rect 287590 577324 287618 585344
rect 287635 585300 287680 585311
rect 288111 585300 288156 585311
rect 287646 577324 287680 585300
rect 287706 581454 287918 581460
rect 287706 581012 288110 581454
rect 287898 581006 288110 581012
rect 288122 577324 288156 585300
rect 288198 577280 288226 585344
rect 288254 577280 288282 585344
rect 288293 585300 288338 585311
rect 288769 585300 288814 585311
rect 288304 577324 288338 585300
rect 288374 581442 288586 581454
rect 288374 581006 288754 581442
rect 288542 580994 288754 581006
rect 288780 577324 288814 585300
rect 288850 583560 288878 584776
rect 288850 577400 288878 579092
rect 288906 577280 288934 585344
rect 288951 585300 288996 585311
rect 288962 577324 288996 585300
rect 289076 577274 289110 585350
rect 289207 583681 289622 585447
rect 291111 585379 291145 585417
rect 292761 585395 292772 585406
rect 292784 585395 292795 585406
rect 292761 585379 292795 585395
rect 290735 585345 293171 585379
rect 289972 583681 289978 584776
rect 290015 583681 290049 583715
rect 290673 583681 290707 583715
rect 291111 583681 291145 585345
rect 291214 585286 291270 585297
rect 291320 585286 291376 585297
rect 291872 585286 291928 585297
rect 291978 585286 292034 585297
rect 292530 585286 292586 585297
rect 292636 585286 292692 585297
rect 291225 583681 291270 585286
rect 291282 583681 291293 584962
rect 291331 583681 291376 585286
rect 291883 583681 291928 585286
rect 291989 584962 292034 585286
rect 291955 583681 291968 584962
rect 291983 583681 292034 584962
rect 292541 583681 292586 585286
rect 292604 583681 292609 584962
rect 292647 583681 292692 585286
rect 292761 583681 292795 585345
rect 289207 583647 292795 583681
rect 289207 583579 289622 583647
rect 289972 583640 289978 583647
rect 290015 583626 290049 583647
rect 290673 583626 290707 583647
rect 289987 583613 290049 583626
rect 290645 583613 290707 583626
rect 289987 583585 290055 583613
rect 290645 583585 290713 583613
rect 289981 583579 290055 583585
rect 290065 583579 290083 583585
rect 290639 583579 290713 583585
rect 290723 583579 290741 583585
rect 291111 583579 291145 583647
rect 291225 583644 291270 583647
rect 291282 583646 291293 583647
rect 291331 583644 291376 583647
rect 291883 583644 291928 583647
rect 291225 583626 291265 583644
rect 291331 583626 291365 583644
rect 291225 583595 291272 583626
rect 291213 583585 291272 583595
rect 291303 583585 291365 583626
rect 291883 583626 291917 583644
rect 291955 583640 291968 583647
rect 291983 583644 292034 583647
rect 292541 583644 292586 583647
rect 291983 583626 292024 583644
rect 291883 583595 291930 583626
rect 291213 583584 291365 583585
rect 291213 583579 291272 583584
rect 291297 583579 291365 583584
rect 291871 583585 291930 583595
rect 291961 583585 292024 583626
rect 292541 583626 292575 583644
rect 292576 583626 292581 583644
rect 292541 583595 292588 583626
rect 292604 583616 292609 583647
rect 292647 583644 292692 583647
rect 292647 583626 292681 583644
rect 291871 583584 292024 583585
rect 291871 583579 291930 583584
rect 291955 583579 292023 583584
rect 292529 583579 292588 583595
rect 292619 583585 292681 583626
rect 292613 583579 292681 583585
rect 289207 583545 290055 583579
rect 290061 583545 290713 583579
rect 290719 583545 291365 583579
rect 291377 583545 292023 583579
rect 292035 583545 292681 583579
rect 289207 578480 289622 583545
rect 289981 583539 289999 583545
rect 290009 583511 290055 583545
rect 290065 583539 290083 583545
rect 290639 583539 290657 583545
rect 290667 583511 290713 583545
rect 290723 583539 290741 583545
rect 290015 578480 290049 583511
rect 290673 578680 290707 583511
rect 290652 578480 290726 578680
rect 289207 578446 289920 578480
rect 289207 577948 289622 578446
rect 289744 578378 289791 578425
rect 289706 578344 289791 578378
rect 289633 578285 289678 578296
rect 289761 578285 289806 578296
rect 289644 578109 289678 578285
rect 289772 578109 289806 578285
rect 289744 578050 289791 578097
rect 289706 578016 289791 578050
rect 289886 577948 289920 578446
rect 289207 577914 289920 577948
rect 290006 578446 290396 578480
rect 290006 578384 290049 578446
rect 290006 577948 290040 578384
rect 290220 578378 290267 578425
rect 290182 578344 290267 578378
rect 290109 578285 290154 578296
rect 290237 578285 290282 578296
rect 290120 578109 290154 578285
rect 290248 578109 290282 578285
rect 290220 578050 290267 578097
rect 290182 578016 290267 578050
rect 290362 577948 290396 578446
rect 290006 577914 290396 577948
rect 290482 578446 290872 578480
rect 290482 577948 290516 578446
rect 290562 578292 290580 578325
rect 290652 578301 290726 578446
rect 290652 578297 290741 578301
rect 290590 578296 290608 578297
rect 290652 578296 290754 578297
rect 290585 578285 290630 578296
rect 290596 578109 290630 578285
rect 290652 578109 290758 578296
rect 290652 578097 290754 578109
rect 290604 578096 290630 578097
rect 290632 578093 290741 578097
rect 290632 578068 290726 578093
rect 290652 578040 290726 578068
rect 290632 578026 290726 578040
rect 290632 577976 290722 578026
rect 290616 577962 290632 577964
rect 290673 577948 290707 577976
rect 290838 577948 290872 578446
rect 290482 577914 290872 577948
rect 289207 577864 289622 577914
rect 289207 577298 289934 577864
rect 289988 577298 290410 577864
rect 290464 577298 290886 577864
rect 289207 577274 290886 577298
rect 285734 577251 290886 577274
rect 291111 577298 291145 583545
rect 291213 583498 291271 583545
rect 291297 583539 291315 583545
rect 291325 583511 291365 583545
rect 291225 583254 291259 583498
rect 291225 581790 291265 583254
rect 291282 581846 291293 583198
rect 291225 577310 291259 581790
rect 291297 577942 291300 579036
rect 291325 577942 291328 579064
rect 291297 577634 291300 577742
rect 291325 577606 291328 577742
rect 291331 577298 291365 583511
rect 291871 583498 291929 583545
rect 291955 583539 291973 583545
rect 291983 583511 292023 583545
rect 291444 581480 291656 581488
rect 291444 581040 291806 581480
rect 291594 581032 291806 581040
rect 291883 579058 291917 583498
rect 291883 577544 291923 579058
rect 291883 577310 291917 577544
rect 291989 577298 292023 583511
rect 292529 583498 292587 583545
rect 292613 583539 292631 583545
rect 292641 583511 292681 583545
rect 292120 581032 292452 581480
rect 292541 577310 292575 583498
rect 292576 581788 292581 583196
rect 292604 581816 292609 583168
rect 292647 579080 292681 583511
rect 292641 577566 292681 579080
rect 292647 577298 292681 577566
rect 292761 581488 292795 583647
rect 294278 583686 294699 585447
rect 296182 585384 296216 585431
rect 297832 585400 297843 585411
rect 297855 585400 297866 585411
rect 297832 585384 297866 585400
rect 296182 585350 297866 585384
rect 295086 583686 295120 583720
rect 295744 583686 295778 583720
rect 296182 583686 296216 585350
rect 296285 585300 296330 585311
rect 296391 585300 296436 585311
rect 296943 585300 296988 585311
rect 297049 585300 297094 585311
rect 297601 585300 297646 585311
rect 297707 585300 297752 585311
rect 296296 584774 296330 585300
rect 296296 583686 296336 584774
rect 296362 583686 296364 584718
rect 296402 583686 296436 585300
rect 296954 583686 296988 585300
rect 297060 584792 297094 585300
rect 297026 583686 297046 584736
rect 297054 583686 297102 584792
rect 297612 584748 297646 585300
rect 297612 583686 297652 584748
rect 297670 583686 297680 584720
rect 297718 583686 297752 585300
rect 297832 583686 297866 585350
rect 294278 583652 297866 583686
rect 294278 583584 294699 583652
rect 295086 583622 295120 583652
rect 295744 583622 295778 583652
rect 295058 583618 295120 583622
rect 295716 583618 295778 583622
rect 295058 583590 295126 583618
rect 295716 583590 295784 583618
rect 295052 583584 295126 583590
rect 295136 583584 295154 583590
rect 295710 583584 295784 583590
rect 295794 583584 295812 583590
rect 296182 583584 296216 583652
rect 296296 583600 296336 583652
rect 296362 583618 296364 583652
rect 296402 583622 296436 583652
rect 296374 583618 296436 583622
rect 296362 583614 296436 583618
rect 296284 583590 296342 583600
rect 296374 583590 296436 583614
rect 296954 583622 296988 583652
rect 297026 583632 297046 583652
rect 297054 583622 297102 583652
rect 296954 583600 296992 583622
rect 296284 583584 296436 583590
rect 296942 583590 297000 583600
rect 297032 583590 297102 583622
rect 297612 583600 297652 583652
rect 297670 583618 297680 583652
rect 297718 583622 297752 583652
rect 297690 583618 297752 583622
rect 297670 583616 297752 583618
rect 296942 583584 297102 583590
rect 297600 583590 297658 583600
rect 297690 583590 297752 583616
rect 297600 583588 297752 583590
rect 297600 583584 297658 583588
rect 297684 583584 297752 583588
rect 294278 583550 295126 583584
rect 295132 583550 295784 583584
rect 295790 583550 296436 583584
rect 296448 583550 297094 583584
rect 297106 583550 297752 583584
rect 293472 581922 293862 581956
rect 292761 581388 292978 581488
rect 293472 581480 293506 581922
rect 293686 581854 293733 581901
rect 293648 581820 293733 581854
rect 293575 581761 293620 581772
rect 293703 581761 293748 581772
rect 293586 581585 293620 581761
rect 293714 581585 293748 581761
rect 293686 581526 293733 581573
rect 293648 581516 293733 581526
rect 293622 581492 293733 581516
rect 293622 581480 293712 581492
rect 293462 581452 293712 581480
rect 293462 581424 293674 581452
rect 293828 581424 293862 581922
rect 294278 581480 294699 583550
rect 295052 583544 295070 583550
rect 295080 583516 295126 583550
rect 295136 583544 295154 583550
rect 295710 583544 295728 583550
rect 295738 583516 295784 583550
rect 295794 583544 295812 583550
rect 293462 581390 293862 581424
rect 294108 581460 294699 581480
rect 292761 581256 293014 581388
rect 293462 581340 293674 581390
rect 294108 581388 294884 581460
rect 292761 581040 292978 581256
rect 291111 577251 291158 577298
rect 291319 577251 291378 577298
rect 291977 577251 292036 577298
rect 292635 577251 292693 577298
rect 285734 577244 292693 577251
rect 285734 577240 290055 577244
rect 285666 577178 285694 577234
rect 285766 577224 285824 577240
rect 285778 577172 285812 577206
rect 286034 577172 286068 577240
rect 286424 577224 286482 577240
rect 287082 577224 287140 577240
rect 287094 577209 287140 577224
rect 286400 577172 286430 577180
rect 286436 577172 286470 577206
rect 286476 577172 286508 577180
rect 287094 577172 287128 577209
rect 287208 577172 287242 577240
rect 287534 577228 287562 577234
rect 288198 577222 288226 577234
rect 288254 577228 288282 577234
rect 288906 577222 288934 577234
rect 289076 577224 289110 577240
rect 289076 577213 289087 577224
rect 289099 577213 289110 577224
rect 289207 577217 290055 577240
rect 289207 577172 289622 577217
rect 289981 577211 289999 577217
rect 290009 577183 290055 577217
rect 290065 577217 290692 577244
rect 290695 577239 290713 577244
rect 290723 577239 292693 577244
rect 290695 577224 292693 577239
rect 290065 577211 290083 577217
rect 285558 577149 289622 577172
rect 290015 577149 290049 577183
rect 290673 577179 290683 577217
rect 290697 577179 290707 577224
rect 290735 577217 292693 577224
rect 291111 577149 291145 577217
rect 291319 577201 291377 577217
rect 291924 577211 292035 577217
rect 291977 577202 292035 577211
rect 291952 577201 292035 577202
rect 292635 577201 292693 577217
rect 291952 577183 291983 577201
rect 292678 577186 292693 577201
rect 292761 577149 292795 581040
rect 293458 580720 293880 581340
rect 294036 581312 294884 581388
rect 294108 581032 294884 581312
rect 294278 581012 294884 581032
rect 293472 580122 293862 580156
rect 293472 579624 293506 580122
rect 293686 580054 293733 580101
rect 293648 580020 293733 580054
rect 293828 580094 293862 580122
rect 293575 579961 293620 579972
rect 293703 579961 293748 579972
rect 293586 579785 293620 579961
rect 293714 579785 293748 579961
rect 293686 579764 293733 579773
rect 293556 579748 293634 579764
rect 293686 579748 293766 579764
rect 293686 579736 293733 579748
rect 293584 579720 293634 579736
rect 293686 579726 293738 579736
rect 293648 579720 293738 579726
rect 293648 579692 293733 579720
rect 293828 579686 293896 580094
rect 293828 579624 293862 579686
rect 293472 579590 293862 579624
rect 293458 578920 293880 579540
rect 294278 577274 294699 581012
rect 295086 577312 295120 583516
rect 295744 581992 295778 583516
rect 295304 581354 295778 581992
rect 295338 581304 295550 581354
rect 295338 581270 295712 581304
rect 295338 581234 295550 581270
rect 295554 581234 295592 581240
rect 295338 581168 295592 581234
rect 295338 581008 295550 581168
rect 295553 581118 295598 581129
rect 295362 580790 295396 581008
rect 295476 580942 295510 581008
rect 295564 580942 295598 581118
rect 295554 580892 295592 580930
rect 295520 580858 295592 580892
rect 295678 580790 295712 581270
rect 295362 580756 295712 580790
rect 295744 577312 295778 581354
rect 295986 581312 295988 581400
rect 295058 577308 295120 577312
rect 295716 577308 295778 577312
rect 296182 577312 296216 583550
rect 296284 583512 296342 583550
rect 296368 583544 296386 583550
rect 296396 583516 296436 583550
rect 296296 582974 296330 583512
rect 296296 581758 296336 582974
rect 296362 581814 296364 582918
rect 296296 577324 296330 581758
rect 296402 577312 296436 583516
rect 296942 583512 297000 583550
rect 297026 583544 297044 583550
rect 297054 583516 297094 583550
rect 296540 581454 296752 581460
rect 296540 581012 296866 581454
rect 296654 581006 296866 581012
rect 296954 579036 296988 583512
rect 296954 577522 296994 579036
rect 296954 577324 296988 577522
rect 297060 577312 297094 583516
rect 297600 583512 297658 583550
rect 297684 583544 297702 583550
rect 297712 583516 297752 583550
rect 297612 582948 297646 583512
rect 297612 581788 297652 582948
rect 297670 581816 297680 582920
rect 297206 581442 297418 581456
rect 297206 581008 297510 581442
rect 297298 580994 297510 581008
rect 297612 577324 297646 581788
rect 297718 579072 297752 583516
rect 297712 577558 297752 579072
rect 297718 577312 297752 577558
rect 295058 577280 295126 577308
rect 295716 577280 295784 577308
rect 295052 577274 295126 577280
rect 295136 577274 295154 577280
rect 295710 577274 295784 577280
rect 295794 577274 295812 577280
rect 296182 577274 296220 577312
rect 296390 577274 296448 577312
rect 297048 577274 297106 577312
rect 297706 577274 297764 577312
rect 297832 577274 297866 583652
rect 298910 578516 298984 578660
rect 298250 577878 298712 578516
rect 298726 577878 299188 578516
rect 300288 577962 300408 577982
rect 300594 577964 300834 578516
rect 300594 577962 300884 577964
rect 300282 577934 300436 577954
rect 300594 577936 300834 577962
rect 300594 577934 300912 577936
rect 300594 577878 300834 577934
rect 298304 577794 298654 577828
rect 298304 577766 298338 577794
rect 298270 577732 298338 577766
rect 298304 577314 298338 577732
rect 298496 577726 298534 577764
rect 298462 577692 298534 577726
rect 298407 577642 298452 577653
rect 298495 577642 298540 577653
rect 298418 577466 298452 577642
rect 298506 577466 298540 577642
rect 298496 577416 298534 577454
rect 298462 577382 298534 577416
rect 298620 577314 298654 577794
rect 298304 577280 298654 577314
rect 298780 577794 299130 577828
rect 298780 577314 298814 577794
rect 298904 577742 298928 577760
rect 298972 577742 299010 577764
rect 298904 577726 299010 577742
rect 298922 577692 299010 577726
rect 298922 577676 298974 577692
rect 298928 577654 298970 577676
rect 298982 577654 298996 577658
rect 298883 577642 298916 577653
rect 298928 577642 298962 577654
rect 298894 577578 298962 577642
rect 298974 577653 299012 577654
rect 298894 577466 298968 577578
rect 298928 577454 298968 577466
rect 298974 577466 299016 577653
rect 298974 577454 299012 577466
rect 298928 577450 298970 577454
rect 298904 577432 298970 577450
rect 298972 577432 299010 577454
rect 298904 577416 299010 577432
rect 298922 577382 299010 577416
rect 298922 577366 298974 577382
rect 298928 577324 298962 577348
rect 299096 577314 299130 577794
rect 298780 577280 299130 577314
rect 294278 577240 295126 577274
rect 295132 577240 295784 577274
rect 295790 577240 298242 577274
rect 298332 577240 298900 577274
rect 294278 577172 294699 577240
rect 295052 577234 295070 577240
rect 295080 577206 295126 577240
rect 295136 577234 295154 577240
rect 295674 577234 295728 577240
rect 295738 577216 295784 577240
rect 295794 577234 295838 577240
rect 295702 577206 295810 577216
rect 295086 577172 295120 577206
rect 295744 577172 295778 577206
rect 296182 577172 296216 577240
rect 296390 577224 296448 577240
rect 297048 577224 297106 577240
rect 297706 577224 297764 577240
rect 297749 577209 297764 577224
rect 297832 577172 297866 577240
rect 294278 577149 299638 577172
rect 285558 577138 299638 577149
rect 280049 576960 280083 576994
rect 279382 576926 279772 576960
rect 279382 576898 279416 576926
rect 279382 576490 279450 576898
rect 279596 576858 279643 576905
rect 279558 576824 279643 576858
rect 279485 576765 279530 576776
rect 279613 576765 279658 576776
rect 279496 576589 279530 576765
rect 279624 576589 279658 576765
rect 279596 576530 279643 576577
rect 279558 576496 279643 576530
rect 279382 576428 279416 576490
rect 279738 576428 279772 576926
rect 279382 576394 279772 576428
rect 279858 576926 280248 576960
rect 279858 576428 279892 576926
rect 280049 576892 280096 576905
rect 280049 576880 280106 576892
rect 280028 576824 280106 576880
rect 279938 576772 279956 576805
rect 280028 576781 280102 576824
rect 280028 576777 280117 576781
rect 279966 576776 279984 576777
rect 280028 576776 280130 576777
rect 279961 576765 280006 576776
rect 279972 576589 280006 576765
rect 280028 576770 280134 576776
rect 280028 576766 280140 576770
rect 280028 576589 280134 576766
rect 280028 576586 280130 576589
rect 280028 576577 280140 576586
rect 279980 576576 280006 576577
rect 280008 576573 280117 576577
rect 280008 576564 280102 576573
rect 280008 576548 280106 576564
rect 280028 576520 280106 576548
rect 280008 576496 280106 576520
rect 280008 576456 280102 576496
rect 279992 576442 280008 576444
rect 280028 576428 280102 576456
rect 280114 576428 280116 576573
rect 280214 576428 280248 576926
rect 279858 576394 280248 576428
rect 280028 576344 280102 576394
rect 278699 575760 278722 575834
rect 278727 575732 278750 575834
rect 279364 575724 279786 576344
rect 279840 575724 280262 576344
rect 282137 575411 282171 577115
rect 283654 577079 284551 577115
rect 286436 575524 286470 577138
rect 286700 576328 286704 576648
rect 286738 576328 286742 576648
rect 287094 575524 287128 577138
rect 287208 575434 287242 577138
rect 289207 577115 294699 577138
rect 289207 577102 289622 577115
rect 288102 576284 288342 576716
rect 287882 576264 287926 576284
rect 288102 576264 288402 576284
rect 288102 576250 288342 576264
rect 287882 576230 287892 576250
rect 288102 576230 288368 576250
rect 288102 576078 288342 576230
rect 292761 575411 292795 577115
rect 294278 577079 294699 577115
rect 295086 575524 295120 577138
rect 297060 575524 297094 577138
rect 297832 575434 297866 577138
rect 298726 576284 298966 576716
rect 298412 576264 298550 576284
rect 298726 576264 299026 576284
rect 298726 576250 298966 576264
rect 298446 576230 298516 576250
rect 298726 576230 298992 576250
rect 298726 576078 298966 576230
rect 278998 574982 279198 575026
rect 278970 574954 279226 574970
rect 232548 568506 232582 574864
rect 232632 569684 232656 569842
rect 232670 569722 232694 569804
rect 232966 569110 233428 569748
rect 233442 569110 233904 569748
rect 235975 569712 236009 571478
rect 236051 569722 236052 569804
rect 236089 569746 236090 569842
rect 236089 569712 236150 569746
rect 235936 569678 236212 569712
rect 235975 569610 236009 569678
rect 235982 569567 236009 569610
rect 236077 569576 236083 569657
rect 235941 569325 235970 569533
rect 235975 569291 236009 569567
rect 236089 569517 236123 569678
rect 236064 569341 236123 569517
rect 235982 569248 236009 569291
rect 236070 569258 236074 569284
rect 236077 569248 236083 569329
rect 235975 569214 236009 569248
rect 236089 569214 236123 569341
rect 235956 569194 236056 569214
rect 235975 569186 236009 569194
rect 235950 569180 236056 569186
rect 236089 569180 236150 569214
rect 236178 569180 236212 569678
rect 235936 569146 236212 569180
rect 236298 569678 236688 569712
rect 236298 569180 236332 569678
rect 236512 569610 236559 569657
rect 236474 569576 236559 569610
rect 236401 569517 236446 569528
rect 236529 569517 236574 569528
rect 236412 569341 236446 569517
rect 236540 569341 236574 569517
rect 236512 569282 236559 569329
rect 236474 569248 236559 569282
rect 236654 569180 236688 569678
rect 236298 569146 236688 569180
rect 236836 569168 236846 569518
rect 236864 569168 236874 569546
rect 235970 569134 236009 569146
rect 235975 569096 236009 569134
rect 233280 569060 233308 569094
rect 233020 569026 233370 569060
rect 232656 568552 232670 568574
rect 233020 568546 233054 569026
rect 233212 568958 233250 568996
rect 233178 568924 233250 568958
rect 233210 568916 233232 568920
rect 233123 568874 233168 568885
rect 233188 568882 233196 568912
rect 233238 568888 233260 568920
rect 233280 568912 233290 568924
rect 233216 568885 233224 568886
rect 233246 568885 233256 568888
rect 233211 568874 233256 568885
rect 233134 568698 233168 568874
rect 233222 568698 233256 568874
rect 233246 568686 233256 568698
rect 233212 568682 233256 568686
rect 233212 568648 233250 568682
rect 233280 568660 233294 568912
rect 233280 568648 233290 568660
rect 233178 568614 233250 568648
rect 233302 568580 233314 569026
rect 233280 568556 233314 568580
rect 233302 568552 233314 568556
rect 233336 568546 233370 569026
rect 232618 568512 232634 568540
rect 231850 568472 232582 568506
rect 232590 568506 232606 568512
rect 232590 568484 232610 568506
rect 232602 568472 232610 568484
rect 231850 568456 231884 568472
rect 231850 568445 231861 568456
rect 231873 568445 231884 568456
rect 232548 568456 232582 568472
rect 232548 568445 232559 568456
rect 232571 568445 232582 568456
rect 232636 568438 232644 568540
rect 233020 568512 233370 568546
rect 233496 569026 233846 569060
rect 233496 568546 233530 569026
rect 233688 568958 233726 568996
rect 233654 568924 233726 568958
rect 233599 568874 233644 568885
rect 233687 568874 233732 568885
rect 233610 568698 233644 568874
rect 233698 568698 233732 568874
rect 233688 568648 233726 568686
rect 233654 568614 233726 568648
rect 233812 568546 233846 569026
rect 233496 568512 233846 568546
rect 232684 568480 233252 568506
rect 232684 568472 233254 568480
rect 233302 568438 233318 568512
rect 233330 568466 233346 568512
rect 235939 568476 236226 569096
rect 236280 568476 236702 569096
rect 236836 568694 236846 568982
rect 236864 568666 236874 568982
rect 236111 568415 236138 568476
rect 236139 568443 236166 568476
rect 228994 568381 235306 568404
rect 223822 568334 223867 568380
rect 223923 568370 235306 568381
rect 223923 568347 230367 568370
rect 223822 567714 223856 568334
rect 223923 568311 227296 568347
rect 227814 568340 227934 568347
rect 228290 568340 228410 568342
rect 228994 568334 230367 568347
rect 227808 568326 227962 568332
rect 227714 568313 228036 568326
rect 228190 568313 228512 568326
rect 227808 568312 227962 568313
rect 228262 568312 228438 568313
rect 223822 567702 223862 567714
rect 223844 567690 223862 567702
rect 223928 567690 223962 568311
rect 224480 568002 224520 568311
rect 224480 567702 224514 568002
rect 224586 567690 224620 568311
rect 225138 567702 225172 568311
rect 225182 568002 225204 568084
rect 225238 568002 225278 568311
rect 225290 568160 225312 568311
rect 225244 567690 225278 568002
rect 223242 567658 223310 567686
rect 223236 567652 223310 567658
rect 223320 567652 223338 567658
rect 223708 567652 223746 567690
rect 223806 567658 223844 567690
rect 223862 567658 223872 567690
rect 223916 567652 223974 567690
rect 224574 567652 224632 567690
rect 225232 567652 225290 567690
rect 225358 567652 225392 568311
rect 225776 568256 226238 568311
rect 226252 568256 226714 568311
rect 228120 568256 228360 568311
rect 225638 568206 226100 568228
rect 225638 568172 226180 568206
rect 225638 567692 226100 568172
rect 226146 567692 226180 568172
rect 225638 567658 226180 567692
rect 226306 568172 226656 568206
rect 226306 567692 226340 568172
rect 226430 568120 226454 568138
rect 226498 568120 226536 568142
rect 226430 568104 226536 568120
rect 226448 568070 226536 568104
rect 226448 568054 226500 568070
rect 226454 568032 226496 568054
rect 226508 568032 226522 568036
rect 226409 568020 226442 568031
rect 226454 568020 226488 568032
rect 226420 567844 226488 568020
rect 226454 567832 226488 567844
rect 226500 568031 226538 568032
rect 226500 567844 226542 568031
rect 226580 568022 226604 568088
rect 226500 567832 226538 567844
rect 226454 567828 226496 567832
rect 226430 567810 226496 567828
rect 226498 567810 226536 567832
rect 226430 567794 226536 567810
rect 226448 567760 226536 567794
rect 226448 567744 226500 567760
rect 226454 567702 226488 567726
rect 226622 567692 226656 568172
rect 227296 568058 227496 568084
rect 227852 568062 227894 568084
rect 235024 568050 235096 568058
rect 235024 568048 235092 568050
rect 228370 568002 228384 568028
rect 235106 567830 235126 568009
rect 235106 567809 235136 567830
rect 226306 567658 226656 567692
rect 225638 567652 226100 567658
rect 214734 567622 220697 567629
rect 214734 567618 217575 567622
rect 213962 567550 213996 567584
rect 214620 567550 214654 567587
rect 214734 567550 214768 567618
rect 216602 567602 216636 567618
rect 216602 567591 216613 567602
rect 216625 567591 216636 567602
rect 216733 567595 217575 567618
rect 217603 567595 218218 567622
rect 216733 567550 217148 567595
rect 213084 567527 217148 567550
rect 217541 567527 217575 567595
rect 218199 567557 218209 567595
rect 218223 567557 218233 567622
rect 218261 567595 220697 567622
rect 221804 567618 222646 567652
rect 222674 567618 223310 567652
rect 223316 567624 226426 567652
rect 223316 567618 225290 567624
rect 218637 567527 218671 567595
rect 218845 567579 218903 567595
rect 219503 567579 219561 567595
rect 219548 567527 219549 567579
rect 219586 567560 219587 567595
rect 220024 567560 220028 567595
rect 220062 567560 220066 567595
rect 220161 567579 220219 567595
rect 220173 567564 220219 567579
rect 220173 567527 220207 567564
rect 220287 567527 220321 567595
rect 221804 567550 222225 567618
rect 222612 567564 222646 567618
rect 223200 567612 223254 567618
rect 223264 567594 223310 567618
rect 223320 567612 223364 567618
rect 223228 567584 223336 567594
rect 222578 567550 222588 567564
rect 222606 567550 222646 567564
rect 223270 567550 223304 567584
rect 223708 567550 223742 567618
rect 223806 567550 223844 567612
rect 223862 567550 223872 567612
rect 223916 567602 223974 567618
rect 224574 567602 224632 567618
rect 225232 567602 225290 567618
rect 225275 567587 225290 567602
rect 225358 567618 226426 567624
rect 225358 567550 225392 567618
rect 225638 567590 226100 567618
rect 221804 567527 227164 567550
rect 213084 567516 227164 567527
rect 206908 567304 207298 567338
rect 206908 567276 206942 567304
rect 206908 566868 206976 567276
rect 207122 567236 207169 567283
rect 207084 567202 207169 567236
rect 207011 567143 207056 567154
rect 207139 567143 207184 567154
rect 207022 566967 207056 567143
rect 207150 566967 207184 567143
rect 207122 566908 207169 566955
rect 207084 566874 207169 566908
rect 206908 566806 206942 566868
rect 207264 566806 207298 567304
rect 206908 566772 207298 566806
rect 207384 567304 207774 567338
rect 207384 566806 207418 567304
rect 207575 567283 207609 567304
rect 207575 567270 207622 567283
rect 207575 567258 207632 567270
rect 207554 567202 207632 567258
rect 207554 567159 207628 567202
rect 207554 567155 207643 567159
rect 207554 567154 207656 567155
rect 207487 567143 207532 567154
rect 207498 566967 207532 567143
rect 207554 566967 207660 567154
rect 207554 566955 207656 566967
rect 207554 566951 207643 566955
rect 207554 566942 207628 566951
rect 207554 566898 207632 566942
rect 207534 566874 207632 566898
rect 207534 566834 207628 566874
rect 207482 566814 207534 566822
rect 207554 566806 207628 566834
rect 207642 566814 207696 566850
rect 207640 566806 207642 566814
rect 207740 566806 207774 567304
rect 207384 566772 207774 566806
rect 207482 566758 207534 566772
rect 207554 566722 207628 566772
rect 207642 566758 207696 566772
rect 206225 566138 206248 566212
rect 206253 566110 206276 566212
rect 206890 566102 207312 566722
rect 207366 566102 207788 566722
rect 209549 565888 209583 567493
rect 209663 565789 209697 567493
rect 211180 567457 212077 567493
rect 211954 567456 211964 567457
rect 211982 567456 212020 567457
rect 212604 567148 212618 567456
rect 213962 565902 213996 567516
rect 214226 566706 214230 567026
rect 214264 566706 214268 567026
rect 214620 565902 214654 567516
rect 214734 565812 214768 567516
rect 216733 567493 222225 567516
rect 216733 567480 217148 567493
rect 215628 566662 215868 567094
rect 215408 566642 215452 566662
rect 215628 566642 215928 566662
rect 215628 566628 215868 566642
rect 215408 566608 215418 566628
rect 215628 566608 215894 566628
rect 215628 566456 215868 566608
rect 220173 565888 220207 567493
rect 220287 565789 220321 567493
rect 221804 567457 222225 567493
rect 222578 567456 222588 567516
rect 222606 567456 222646 567516
rect 222612 565902 222646 567456
rect 223228 567148 223242 567456
rect 223806 567148 223844 567516
rect 223862 567148 223872 567516
rect 224586 565902 224620 567516
rect 225358 565812 225392 567516
rect 225788 567506 225946 567516
rect 235072 567470 235130 567472
rect 235046 567436 235096 567438
rect 225850 567094 225884 567096
rect 225776 566956 226078 567094
rect 226252 566662 226492 567094
rect 225938 566642 226076 566662
rect 226252 566642 226552 566662
rect 226252 566628 226492 566642
rect 225972 566608 226042 566628
rect 226252 566608 226518 566628
rect 226252 566456 226492 566608
rect 143626 565727 149938 565750
rect 138687 565716 149938 565727
rect 138687 565693 144999 565716
rect 140016 565657 140986 565693
rect 143626 565680 144999 565693
rect 81984 565360 82184 565404
rect 87576 565360 87776 565404
rect 98910 565360 99110 565404
rect 140460 565396 140532 565404
rect 149656 565396 149728 565404
rect 140460 565394 140528 565396
rect 149656 565394 149724 565396
rect 206524 565360 206724 565404
rect 81956 565332 82212 565348
rect 87548 565332 87804 565348
rect 98882 565332 99138 565348
rect 134656 564906 134660 565226
rect 134694 564906 134698 565226
rect 149738 565176 149758 565355
rect 206496 565332 206752 565348
rect 149738 565155 149768 565176
rect 149704 564816 149762 564818
rect 149678 564782 149728 564784
<< metal2 >>
rect 524 -800 636 480
rect 1706 -800 1818 480
rect 2888 -800 3000 480
rect 4070 -800 4182 480
rect 5252 -800 5364 480
rect 6434 -800 6546 480
rect 7616 -800 7728 480
rect 8798 -800 8910 480
rect 9980 -800 10092 480
rect 11162 -800 11274 480
rect 12344 -800 12456 480
rect 13526 -800 13638 480
rect 14708 -800 14820 480
rect 15890 -800 16002 480
rect 17072 -800 17184 480
rect 18254 -800 18366 480
rect 19436 -800 19548 480
rect 20618 -800 20730 480
rect 21800 -800 21912 480
rect 22982 -800 23094 480
rect 24164 -800 24276 480
rect 25346 -800 25458 480
rect 26528 -800 26640 480
rect 27710 -800 27822 480
rect 28892 -800 29004 480
rect 30074 -800 30186 480
rect 31256 -800 31368 480
rect 32438 -800 32550 480
rect 33620 -800 33732 480
rect 34802 -800 34914 480
rect 35984 -800 36096 480
rect 37166 -800 37278 480
rect 38348 -800 38460 480
rect 39530 -800 39642 480
rect 40712 -800 40824 480
rect 41894 -800 42006 480
rect 43076 -800 43188 480
rect 44258 -800 44370 480
rect 45440 -800 45552 480
rect 46622 -800 46734 480
rect 47804 -800 47916 480
rect 48986 -800 49098 480
rect 50168 -800 50280 480
rect 51350 -800 51462 480
rect 52532 -800 52644 480
rect 53714 -800 53826 480
rect 54896 -800 55008 480
rect 56078 -800 56190 480
rect 57260 -800 57372 480
rect 58442 -800 58554 480
rect 59624 -800 59736 480
rect 60806 -800 60918 480
rect 61988 -800 62100 480
rect 63170 -800 63282 480
rect 64352 -800 64464 480
rect 65534 -800 65646 480
rect 66716 -800 66828 480
rect 67898 -800 68010 480
rect 69080 -800 69192 480
rect 70262 -800 70374 480
rect 71444 -800 71556 480
rect 72626 -800 72738 480
rect 73808 -800 73920 480
rect 74990 -800 75102 480
rect 76172 -800 76284 480
rect 77354 -800 77466 480
rect 78536 -800 78648 480
rect 79718 -800 79830 480
rect 80900 -800 81012 480
rect 82082 -800 82194 480
rect 83264 -800 83376 480
rect 84446 -800 84558 480
rect 85628 -800 85740 480
rect 86810 -800 86922 480
rect 87992 -800 88104 480
rect 89174 -800 89286 480
rect 90356 -800 90468 480
rect 91538 -800 91650 480
rect 92720 -800 92832 480
rect 93902 -800 94014 480
rect 95084 -800 95196 480
rect 96266 -800 96378 480
rect 97448 -800 97560 480
rect 98630 -800 98742 480
rect 99812 -800 99924 480
rect 100994 -800 101106 480
rect 102176 -800 102288 480
rect 103358 -800 103470 480
rect 104540 -800 104652 480
rect 105722 -800 105834 480
rect 106904 -800 107016 480
rect 108086 -800 108198 480
rect 109268 -800 109380 480
rect 110450 -800 110562 480
rect 111632 -800 111744 480
rect 112814 -800 112926 480
rect 113996 -800 114108 480
rect 115178 -800 115290 480
rect 116360 -800 116472 480
rect 117542 -800 117654 480
rect 118724 -800 118836 480
rect 119906 -800 120018 480
rect 121088 -800 121200 480
rect 122270 -800 122382 480
rect 123452 -800 123564 480
rect 124634 -800 124746 480
rect 125816 -800 125928 480
rect 126998 -800 127110 480
rect 128180 -800 128292 480
rect 129362 -800 129474 480
rect 130544 -800 130656 480
rect 131726 -800 131838 480
rect 132908 -800 133020 480
rect 134090 -800 134202 480
rect 135272 -800 135384 480
rect 136454 -800 136566 480
rect 137636 -800 137748 480
rect 138818 -800 138930 480
rect 140000 -800 140112 480
rect 141182 -800 141294 480
rect 142364 -800 142476 480
rect 143546 -800 143658 480
rect 144728 -800 144840 480
rect 145910 -800 146022 480
rect 147092 -800 147204 480
rect 148274 -800 148386 480
rect 149456 -800 149568 480
rect 150638 -800 150750 480
rect 151820 -800 151932 480
rect 153002 -800 153114 480
rect 154184 -800 154296 480
rect 155366 -800 155478 480
rect 156548 -800 156660 480
rect 157730 -800 157842 480
rect 158912 -800 159024 480
rect 160094 -800 160206 480
rect 161276 -800 161388 480
rect 162458 -800 162570 480
rect 163640 -800 163752 480
rect 164822 -800 164934 480
rect 166004 -800 166116 480
rect 167186 -800 167298 480
rect 168368 -800 168480 480
rect 169550 -800 169662 480
rect 170732 -800 170844 480
rect 171914 -800 172026 480
rect 173096 -800 173208 480
rect 174278 -800 174390 480
rect 175460 -800 175572 480
rect 176642 -800 176754 480
rect 177824 -800 177936 480
rect 179006 -800 179118 480
rect 180188 -800 180300 480
rect 181370 -800 181482 480
rect 182552 -800 182664 480
rect 183734 -800 183846 480
rect 184916 -800 185028 480
rect 186098 -800 186210 480
rect 187280 -800 187392 480
rect 188462 -800 188574 480
rect 189644 -800 189756 480
rect 190826 -800 190938 480
rect 192008 -800 192120 480
rect 193190 -800 193302 480
rect 194372 -800 194484 480
rect 195554 -800 195666 480
rect 196736 -800 196848 480
rect 197918 -800 198030 480
rect 199100 -800 199212 480
rect 200282 -800 200394 480
rect 201464 -800 201576 480
rect 202646 -800 202758 480
rect 203828 -800 203940 480
rect 205010 -800 205122 480
rect 206192 -800 206304 480
rect 207374 -800 207486 480
rect 208556 -800 208668 480
rect 209738 -800 209850 480
rect 210920 -800 211032 480
rect 212102 -800 212214 480
rect 213284 -800 213396 480
rect 214466 -800 214578 480
rect 215648 -800 215760 480
rect 216830 -800 216942 480
rect 218012 -800 218124 480
rect 219194 -800 219306 480
rect 220376 -800 220488 480
rect 221558 -800 221670 480
rect 222740 -800 222852 480
rect 223922 -800 224034 480
rect 225104 -800 225216 480
rect 226286 -800 226398 480
rect 227468 -800 227580 480
rect 228650 -800 228762 480
rect 229832 -800 229944 480
rect 231014 -800 231126 480
rect 232196 -800 232308 480
rect 233378 -800 233490 480
rect 234560 -800 234672 480
rect 235742 -800 235854 480
rect 236924 -800 237036 480
rect 238106 -800 238218 480
rect 239288 -800 239400 480
rect 240470 -800 240582 480
rect 241652 -800 241764 480
rect 242834 -800 242946 480
rect 244016 -800 244128 480
rect 245198 -800 245310 480
rect 246380 -800 246492 480
rect 247562 -800 247674 480
rect 248744 -800 248856 480
rect 249926 -800 250038 480
rect 251108 -800 251220 480
rect 252290 -800 252402 480
rect 253472 -800 253584 480
rect 254654 -800 254766 480
rect 255836 -800 255948 480
rect 257018 -800 257130 480
rect 258200 -800 258312 480
rect 259382 -800 259494 480
rect 260564 -800 260676 480
rect 261746 -800 261858 480
rect 262928 -800 263040 480
rect 264110 -800 264222 480
rect 265292 -800 265404 480
rect 266474 -800 266586 480
rect 267656 -800 267768 480
rect 268838 -800 268950 480
rect 270020 -800 270132 480
rect 271202 -800 271314 480
rect 272384 -800 272496 480
rect 273566 -800 273678 480
rect 274748 -800 274860 480
rect 275930 -800 276042 480
rect 277112 -800 277224 480
rect 278294 -800 278406 480
rect 279476 -800 279588 480
rect 280658 -800 280770 480
rect 281840 -800 281952 480
rect 283022 -800 283134 480
rect 284204 -800 284316 480
rect 285386 -800 285498 480
rect 286568 -800 286680 480
rect 287750 -800 287862 480
rect 288932 -800 289044 480
rect 290114 -800 290226 480
rect 291296 -800 291408 480
rect 292478 -800 292590 480
rect 293660 -800 293772 480
rect 294842 -800 294954 480
rect 296024 -800 296136 480
rect 297206 -800 297318 480
rect 298388 -800 298500 480
rect 299570 -800 299682 480
rect 300752 -800 300864 480
rect 301934 -800 302046 480
rect 303116 -800 303228 480
rect 304298 -800 304410 480
rect 305480 -800 305592 480
rect 306662 -800 306774 480
rect 307844 -800 307956 480
rect 309026 -800 309138 480
rect 310208 -800 310320 480
rect 311390 -800 311502 480
rect 312572 -800 312684 480
rect 313754 -800 313866 480
rect 314936 -800 315048 480
rect 316118 -800 316230 480
rect 317300 -800 317412 480
rect 318482 -800 318594 480
rect 319664 -800 319776 480
rect 320846 -800 320958 480
rect 322028 -800 322140 480
rect 323210 -800 323322 480
rect 324392 -800 324504 480
rect 325574 -800 325686 480
rect 326756 -800 326868 480
rect 327938 -800 328050 480
rect 329120 -800 329232 480
rect 330302 -800 330414 480
rect 331484 -800 331596 480
rect 332666 -800 332778 480
rect 333848 -800 333960 480
rect 335030 -800 335142 480
rect 336212 -800 336324 480
rect 337394 -800 337506 480
rect 338576 -800 338688 480
rect 339758 -800 339870 480
rect 340940 -800 341052 480
rect 342122 -800 342234 480
rect 343304 -800 343416 480
rect 344486 -800 344598 480
rect 345668 -800 345780 480
rect 346850 -800 346962 480
rect 348032 -800 348144 480
rect 349214 -800 349326 480
rect 350396 -800 350508 480
rect 351578 -800 351690 480
rect 352760 -800 352872 480
rect 353942 -800 354054 480
rect 355124 -800 355236 480
rect 356306 -800 356418 480
rect 357488 -800 357600 480
rect 358670 -800 358782 480
rect 359852 -800 359964 480
rect 361034 -800 361146 480
rect 362216 -800 362328 480
rect 363398 -800 363510 480
rect 364580 -800 364692 480
rect 365762 -800 365874 480
rect 366944 -800 367056 480
rect 368126 -800 368238 480
rect 369308 -800 369420 480
rect 370490 -800 370602 480
rect 371672 -800 371784 480
rect 372854 -800 372966 480
rect 374036 -800 374148 480
rect 375218 -800 375330 480
rect 376400 -800 376512 480
rect 377582 -800 377694 480
rect 378764 -800 378876 480
rect 379946 -800 380058 480
rect 381128 -800 381240 480
rect 382310 -800 382422 480
rect 383492 -800 383604 480
rect 384674 -800 384786 480
rect 385856 -800 385968 480
rect 387038 -800 387150 480
rect 388220 -800 388332 480
rect 389402 -800 389514 480
rect 390584 -800 390696 480
rect 391766 -800 391878 480
rect 392948 -800 393060 480
rect 394130 -800 394242 480
rect 395312 -800 395424 480
rect 396494 -800 396606 480
rect 397676 -800 397788 480
rect 398858 -800 398970 480
rect 400040 -800 400152 480
rect 401222 -800 401334 480
rect 402404 -800 402516 480
rect 403586 -800 403698 480
rect 404768 -800 404880 480
rect 405950 -800 406062 480
rect 407132 -800 407244 480
rect 408314 -800 408426 480
rect 409496 -800 409608 480
rect 410678 -800 410790 480
rect 411860 -800 411972 480
rect 413042 -800 413154 480
rect 414224 -800 414336 480
rect 415406 -800 415518 480
rect 416588 -800 416700 480
rect 417770 -800 417882 480
rect 418952 -800 419064 480
rect 420134 -800 420246 480
rect 421316 -800 421428 480
rect 422498 -800 422610 480
rect 423680 -800 423792 480
rect 424862 -800 424974 480
rect 426044 -800 426156 480
rect 427226 -800 427338 480
rect 428408 -800 428520 480
rect 429590 -800 429702 480
rect 430772 -800 430884 480
rect 431954 -800 432066 480
rect 433136 -800 433248 480
rect 434318 -800 434430 480
rect 435500 -800 435612 480
rect 436682 -800 436794 480
rect 437864 -800 437976 480
rect 439046 -800 439158 480
rect 440228 -800 440340 480
rect 441410 -800 441522 480
rect 442592 -800 442704 480
rect 443774 -800 443886 480
rect 444956 -800 445068 480
rect 446138 -800 446250 480
rect 447320 -800 447432 480
rect 448502 -800 448614 480
rect 449684 -800 449796 480
rect 450866 -800 450978 480
rect 452048 -800 452160 480
rect 453230 -800 453342 480
rect 454412 -800 454524 480
rect 455594 -800 455706 480
rect 456776 -800 456888 480
rect 457958 -800 458070 480
rect 459140 -800 459252 480
rect 460322 -800 460434 480
rect 461504 -800 461616 480
rect 462686 -800 462798 480
rect 463868 -800 463980 480
rect 465050 -800 465162 480
rect 466232 -800 466344 480
rect 467414 -800 467526 480
rect 468596 -800 468708 480
rect 469778 -800 469890 480
rect 470960 -800 471072 480
rect 472142 -800 472254 480
rect 473324 -800 473436 480
rect 474506 -800 474618 480
rect 475688 -800 475800 480
rect 476870 -800 476982 480
rect 478052 -800 478164 480
rect 479234 -800 479346 480
rect 480416 -800 480528 480
rect 481598 -800 481710 480
rect 482780 -800 482892 480
rect 483962 -800 484074 480
rect 485144 -800 485256 480
rect 486326 -800 486438 480
rect 487508 -800 487620 480
rect 488690 -800 488802 480
rect 489872 -800 489984 480
rect 491054 -800 491166 480
rect 492236 -800 492348 480
rect 493418 -800 493530 480
rect 494600 -800 494712 480
rect 495782 -800 495894 480
rect 496964 -800 497076 480
rect 498146 -800 498258 480
rect 499328 -800 499440 480
rect 500510 -800 500622 480
rect 501692 -800 501804 480
rect 502874 -800 502986 480
rect 504056 -800 504168 480
rect 505238 -800 505350 480
rect 506420 -800 506532 480
rect 507602 -800 507714 480
rect 508784 -800 508896 480
rect 509966 -800 510078 480
rect 511148 -800 511260 480
rect 512330 -800 512442 480
rect 513512 -800 513624 480
rect 514694 -800 514806 480
rect 515876 -800 515988 480
rect 517058 -800 517170 480
rect 518240 -800 518352 480
rect 519422 -800 519534 480
rect 520604 -800 520716 480
rect 521786 -800 521898 480
rect 522968 -800 523080 480
rect 524150 -800 524262 480
rect 525332 -800 525444 480
rect 526514 -800 526626 480
rect 527696 -800 527808 480
rect 528878 -800 528990 480
rect 530060 -800 530172 480
rect 531242 -800 531354 480
rect 532424 -800 532536 480
rect 533606 -800 533718 480
rect 534788 -800 534900 480
rect 535970 -800 536082 480
rect 537152 -800 537264 480
rect 538334 -800 538446 480
rect 539516 -800 539628 480
rect 540698 -800 540810 480
rect 541880 -800 541992 480
rect 543062 -800 543174 480
rect 544244 -800 544356 480
rect 545426 -800 545538 480
rect 546608 -800 546720 480
rect 547790 -800 547902 480
rect 548972 -800 549084 480
rect 550154 -800 550266 480
rect 551336 -800 551448 480
rect 552518 -800 552630 480
rect 553700 -800 553812 480
rect 554882 -800 554994 480
rect 556064 -800 556176 480
rect 557246 -800 557358 480
rect 558428 -800 558540 480
rect 559610 -800 559722 480
rect 560792 -800 560904 480
rect 561974 -800 562086 480
rect 563156 -800 563268 480
rect 564338 -800 564450 480
rect 565520 -800 565632 480
rect 566702 -800 566814 480
rect 567884 -800 567996 480
rect 569066 -800 569178 480
rect 570248 -800 570360 480
rect 571430 -800 571542 480
rect 572612 -800 572724 480
rect 573794 -800 573906 480
rect 574976 -800 575088 480
rect 576158 -800 576270 480
rect 577340 -800 577452 480
rect 578522 -800 578634 480
rect 579704 -800 579816 480
rect 580886 -800 580998 480
rect 582068 -800 582180 480
rect 583250 -800 583362 480
<< metal3 >>
rect 16194 702300 21194 704800
rect 68194 702300 73194 704800
rect 120194 702300 125194 704800
rect 165594 702300 170594 704800
rect 170894 702300 173094 704800
rect 173394 702300 175594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 222594 702300 224794 704800
rect 225094 702300 227294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 324294 702300 326494 704800
rect 326794 702300 328994 704800
rect 329294 702300 334294 704800
rect 413394 702300 418394 704800
rect 465394 702300 470394 704800
rect 510594 702340 515394 704800
rect 520594 702340 525394 704800
rect 566594 702300 571594 704800
rect -800 680242 1700 685242
rect 582300 677984 584800 682984
rect -800 643842 1660 648642
rect 582340 639784 584800 644584
rect -800 633842 1660 638642
rect 582340 629784 584800 634584
rect 583520 589472 584800 589584
rect 583520 588290 584800 588402
rect 583520 587108 584800 587220
rect 583520 585926 584800 586038
rect 583520 584744 584800 584856
rect 583520 583562 584800 583674
rect -800 559442 1660 564242
rect -800 549442 1660 554242
rect 582340 550562 584800 555362
rect 582340 540562 584800 545362
rect -800 511530 480 511642
rect -800 510348 480 510460
rect -800 509166 480 509278
rect -800 507984 480 508096
rect -800 506802 480 506914
rect -800 505620 480 505732
rect 583520 500050 584800 500162
rect 583520 498868 584800 498980
rect 583520 497686 584800 497798
rect 583520 496504 584800 496616
rect 583520 495322 584800 495434
rect 583520 494140 584800 494252
rect -800 468308 480 468420
rect -800 467126 480 467238
rect -800 465944 480 466056
rect -800 464762 480 464874
rect -800 463580 480 463692
rect -800 462398 480 462510
rect 583520 455628 584800 455740
rect 583520 454446 584800 454558
rect 583520 453264 584800 453376
rect 583520 452082 584800 452194
rect 583520 450900 584800 451012
rect 583520 449718 584800 449830
rect -800 425086 480 425198
rect -800 423904 480 424016
rect -800 422722 480 422834
rect -800 421540 480 421652
rect -800 420358 480 420470
rect -800 419176 480 419288
rect 583520 411206 584800 411318
rect 583520 410024 584800 410136
rect 583520 408842 584800 408954
rect 583520 407660 584800 407772
rect 583520 406478 584800 406590
rect 583520 405296 584800 405408
rect -800 381864 480 381976
rect -800 380682 480 380794
rect -800 379500 480 379612
rect -800 378318 480 378430
rect -800 377136 480 377248
rect -800 375954 480 376066
rect 583520 364784 584800 364896
rect 583520 363602 584800 363714
rect 583520 362420 584800 362532
rect 583520 361238 584800 361350
rect 583520 360056 584800 360168
rect 583520 358874 584800 358986
rect -800 338642 480 338754
rect -800 337460 480 337572
rect -800 336278 480 336390
rect -800 335096 480 335208
rect -800 333914 480 334026
rect -800 332732 480 332844
rect 583520 319562 584800 319674
rect 583520 318380 584800 318492
rect 583520 317198 584800 317310
rect 583520 316016 584800 316128
rect 583520 314834 584800 314946
rect 583520 313652 584800 313764
rect -800 295420 480 295532
rect -800 294238 480 294350
rect -800 293056 480 293168
rect -800 291874 480 291986
rect -800 290692 480 290804
rect -800 289510 480 289622
rect 583520 275140 584800 275252
rect 583520 273958 584800 274070
rect 583520 272776 584800 272888
rect 583520 271594 584800 271706
rect 583520 270412 584800 270524
rect 583520 269230 584800 269342
rect -800 252398 480 252510
rect -800 251216 480 251328
rect -800 250034 480 250146
rect -800 248852 480 248964
rect -800 247670 480 247782
rect -800 246488 480 246600
rect 582340 235230 584800 240030
rect 582340 225230 584800 230030
rect -800 214888 1660 219688
rect -800 204888 1660 209688
rect 582340 191430 584800 196230
rect 582340 181430 584800 186230
rect -800 172888 1660 177688
rect -800 162888 1660 167688
rect 582340 146830 584800 151630
rect 582340 136830 584800 141630
rect -800 124776 480 124888
rect -800 123594 480 123706
rect -800 122412 480 122524
rect -800 121230 480 121342
rect -800 120048 480 120160
rect -800 118866 480 118978
rect 583520 95118 584800 95230
rect 583520 93936 584800 94048
rect 583520 92754 584800 92866
rect 583520 91572 584800 91684
rect -800 81554 480 81666
rect -800 80372 480 80484
rect -800 79190 480 79302
rect -800 78008 480 78120
rect -800 76826 480 76938
rect -800 75644 480 75756
rect 583520 50460 584800 50572
rect 583520 49278 584800 49390
rect 583520 48096 584800 48208
rect 583520 46914 584800 47026
rect -800 38332 480 38444
rect -800 37150 480 37262
rect -800 35968 480 36080
rect -800 34786 480 34898
rect -800 33604 480 33716
rect -800 32422 480 32534
rect 583520 24002 584800 24114
rect 583520 22820 584800 22932
rect 583520 21638 584800 21750
rect 583520 20456 584800 20568
rect 583520 19274 584800 19386
rect 583520 18092 584800 18204
rect -800 16910 480 17022
rect 583520 16910 584800 17022
rect -800 15728 480 15840
rect 583520 15728 584800 15840
rect -800 14546 480 14658
rect 583520 14546 584800 14658
rect -800 13364 480 13476
rect 583520 13364 584800 13476
rect -800 12182 480 12294
rect 583520 12182 584800 12294
rect -800 11000 480 11112
rect 583520 11000 584800 11112
rect -800 9818 480 9930
rect 583520 9818 584800 9930
rect -800 8636 480 8748
rect 583520 8636 584800 8748
rect -800 7454 480 7566
rect 583520 7454 584800 7566
rect -800 6272 480 6384
rect 583520 6272 584800 6384
rect -800 5090 480 5202
rect 583520 5090 584800 5202
rect -800 3908 480 4020
rect 583520 3908 584800 4020
rect -800 2726 480 2838
rect 583520 2726 584800 2838
rect -800 1544 480 1656
rect 583520 1544 584800 1656
<< metal4 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
<< metal5 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
<< comment >>
rect -100 704000 584100 704100
rect -100 0 0 704000
rect 584000 0 584100 704000
rect -100 -100 584100 0
use sky130_fd_pr__res_generic_m3_DPAT6Q  R1
timestamp 1695461801
transform 1 0 1100 0 1 687
box -1100 -87 1100 87
use sky130_fd_pr__res_generic_m3_DPAT6Q  R2
timestamp 1695461801
transform 1 0 3300 0 1 687
box -1100 -87 1100 87
use sky130_fd_pr__res_generic_m3_DPAT6Q  R4
timestamp 1695461801
transform 1 0 5500 0 1 687
box -1100 -87 1100 87
use sky130_fd_pr__res_generic_m3_DPAT6Q  R5
timestamp 1695461801
transform 1 0 7700 0 1 687
box -1100 -87 1100 87
use sky130_fd_pr__res_generic_m3_DPAT6Q  R6
timestamp 1695461801
transform 1 0 9900 0 1 687
box -1100 -87 1100 87
use sky130_fd_pr__res_generic_m3_DPAT6Q  R7
timestamp 1695461801
transform 1 0 12100 0 1 687
box -1100 -87 1100 87
use sky130_fd_pr__res_generic_m3_2QNVX3  R8
timestamp 1695461801
transform 1 0 13256 0 1 706
box 0 0 1 1
use sky130_fd_pr__res_generic_m3_SS5VKG  R9
timestamp 1695461801
transform 1 0 13368 0 1 688
box -56 -88 56 88
use sky130_fd_pr__res_generic_m3_HK2ST4  R11
timestamp 1695461801
transform 1 0 13480 0 1 715
box -56 -115 56 115
use sky130_fd_pr__res_generic_m3_BHQV68  R12
timestamp 1695461801
transform 1 0 13592 0 1 717
box -56 -117 56 117
use ColROs  x3
timestamp 1695461801
transform 1 0 114976 0 1 573182
box -33468 -9022 186662 48942
<< labels >>
flabel metal3 s 583520 269230 584800 269342 0 FreeSans 1120 0 0 0 gpio_analog[0]
port 0 nsew signal bidirectional
flabel metal3 s -800 381864 480 381976 0 FreeSans 1120 0 0 0 gpio_analog[10]
port 1 nsew signal bidirectional
flabel metal3 s -800 338642 480 338754 0 FreeSans 1120 0 0 0 gpio_analog[11]
port 2 nsew signal bidirectional
flabel metal3 s -800 295420 480 295532 0 FreeSans 1120 0 0 0 gpio_analog[12]
port 3 nsew signal bidirectional
flabel metal3 s -800 252398 480 252510 0 FreeSans 1120 0 0 0 gpio_analog[13]
port 4 nsew signal bidirectional
flabel metal3 s -800 124776 480 124888 0 FreeSans 1120 0 0 0 gpio_analog[14]
port 5 nsew signal bidirectional
flabel metal3 s -800 81554 480 81666 0 FreeSans 1120 0 0 0 gpio_analog[15]
port 6 nsew signal bidirectional
flabel metal3 s -800 38332 480 38444 0 FreeSans 1120 0 0 0 gpio_analog[16]
port 7 nsew signal bidirectional
flabel metal3 s -800 16910 480 17022 0 FreeSans 1120 0 0 0 gpio_analog[17]
port 8 nsew signal bidirectional
flabel metal3 s 583520 313652 584800 313764 0 FreeSans 1120 0 0 0 gpio_analog[1]
port 9 nsew signal bidirectional
flabel metal3 s 583520 358874 584800 358986 0 FreeSans 1120 0 0 0 gpio_analog[2]
port 10 nsew signal bidirectional
flabel metal3 s 583520 405296 584800 405408 0 FreeSans 1120 0 0 0 gpio_analog[3]
port 11 nsew signal bidirectional
flabel metal3 s 583520 449718 584800 449830 0 FreeSans 1120 0 0 0 gpio_analog[4]
port 12 nsew signal bidirectional
flabel metal3 s 583520 494140 584800 494252 0 FreeSans 1120 0 0 0 gpio_analog[5]
port 13 nsew signal bidirectional
flabel metal3 s 583520 583562 584800 583674 0 FreeSans 1120 0 0 0 gpio_analog[6]
port 14 nsew signal bidirectional
flabel metal3 s -800 511530 480 511642 0 FreeSans 1120 0 0 0 gpio_analog[7]
port 15 nsew signal bidirectional
flabel metal3 s -800 468308 480 468420 0 FreeSans 1120 0 0 0 gpio_analog[8]
port 16 nsew signal bidirectional
flabel metal3 s -800 425086 480 425198 0 FreeSans 1120 0 0 0 gpio_analog[9]
port 17 nsew signal bidirectional
flabel metal3 s 583520 270412 584800 270524 0 FreeSans 1120 0 0 0 gpio_noesd[0]
port 18 nsew signal bidirectional
flabel metal3 s -800 380682 480 380794 0 FreeSans 1120 0 0 0 gpio_noesd[10]
port 19 nsew signal bidirectional
flabel metal3 s -800 337460 480 337572 0 FreeSans 1120 0 0 0 gpio_noesd[11]
port 20 nsew signal bidirectional
flabel metal3 s -800 294238 480 294350 0 FreeSans 1120 0 0 0 gpio_noesd[12]
port 21 nsew signal bidirectional
flabel metal3 s -800 251216 480 251328 0 FreeSans 1120 0 0 0 gpio_noesd[13]
port 22 nsew signal bidirectional
flabel metal3 s -800 123594 480 123706 0 FreeSans 1120 0 0 0 gpio_noesd[14]
port 23 nsew signal bidirectional
flabel metal3 s -800 80372 480 80484 0 FreeSans 1120 0 0 0 gpio_noesd[15]
port 24 nsew signal bidirectional
flabel metal3 s -800 37150 480 37262 0 FreeSans 1120 0 0 0 gpio_noesd[16]
port 25 nsew signal bidirectional
flabel metal3 s -800 15728 480 15840 0 FreeSans 1120 0 0 0 gpio_noesd[17]
port 26 nsew signal bidirectional
flabel metal3 s 583520 314834 584800 314946 0 FreeSans 1120 0 0 0 gpio_noesd[1]
port 27 nsew signal bidirectional
flabel metal3 s 583520 360056 584800 360168 0 FreeSans 1120 0 0 0 gpio_noesd[2]
port 28 nsew signal bidirectional
flabel metal3 s 583520 406478 584800 406590 0 FreeSans 1120 0 0 0 gpio_noesd[3]
port 29 nsew signal bidirectional
flabel metal3 s 583520 450900 584800 451012 0 FreeSans 1120 0 0 0 gpio_noesd[4]
port 30 nsew signal bidirectional
flabel metal3 s 583520 495322 584800 495434 0 FreeSans 1120 0 0 0 gpio_noesd[5]
port 31 nsew signal bidirectional
flabel metal3 s 583520 584744 584800 584856 0 FreeSans 1120 0 0 0 gpio_noesd[6]
port 32 nsew signal bidirectional
flabel metal3 s -800 510348 480 510460 0 FreeSans 1120 0 0 0 gpio_noesd[7]
port 33 nsew signal bidirectional
flabel metal3 s -800 467126 480 467238 0 FreeSans 1120 0 0 0 gpio_noesd[8]
port 34 nsew signal bidirectional
flabel metal3 s -800 423904 480 424016 0 FreeSans 1120 0 0 0 gpio_noesd[9]
port 35 nsew signal bidirectional
flabel metal3 s 582300 677984 584800 682984 0 FreeSans 1120 0 0 0 io_analog[0]
port 36 nsew signal bidirectional
flabel metal3 s 0 680242 1700 685242 0 FreeSans 1120 0 0 0 io_analog[10]
port 37 nsew signal bidirectional
flabel metal3 s 566594 702300 571594 704800 0 FreeSans 1920 180 0 0 io_analog[1]
port 38 nsew signal bidirectional
flabel metal3 s 465394 702300 470394 704800 0 FreeSans 1920 180 0 0 io_analog[2]
port 39 nsew signal bidirectional
flabel metal3 s 413394 702300 418394 704800 0 FreeSans 1920 180 0 0 io_analog[3]
port 40 nsew signal bidirectional
flabel metal3 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal4 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal5 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal3 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal4 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal5 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal3 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal4 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal5 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal3 s 120194 702300 125194 704800 0 FreeSans 1920 180 0 0 io_analog[7]
port 44 nsew signal bidirectional
flabel metal3 s 68194 702300 73194 704800 0 FreeSans 1920 180 0 0 io_analog[8]
port 45 nsew signal bidirectional
flabel metal3 s 16194 702300 21194 704800 0 FreeSans 1920 180 0 0 io_analog[9]
port 46 nsew signal bidirectional
flabel metal3 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal4 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal5 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal3 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal4 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal5 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal3 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal4 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal5 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal3 s 326794 702300 328994 704800 0 FreeSans 1920 180 0 0 io_clamp_high[0]
port 50 nsew signal bidirectional
flabel metal3 s 225094 702300 227294 704800 0 FreeSans 1920 180 0 0 io_clamp_high[1]
port 51 nsew signal bidirectional
flabel metal3 s 173394 702300 175594 704800 0 FreeSans 1920 180 0 0 io_clamp_high[2]
port 52 nsew signal bidirectional
flabel metal3 s 324294 702300 326494 704800 0 FreeSans 1920 180 0 0 io_clamp_low[0]
port 53 nsew signal bidirectional
flabel metal3 s 222594 702300 224794 704800 0 FreeSans 1920 180 0 0 io_clamp_low[1]
port 54 nsew signal bidirectional
flabel metal3 s 170894 702300 173094 704800 0 FreeSans 1920 180 0 0 io_clamp_low[2]
port 55 nsew signal bidirectional
flabel metal3 s 583520 2726 584800 2838 0 FreeSans 1120 0 0 0 io_in[0]
port 56 nsew signal input
flabel metal3 s 583520 408842 584800 408954 0 FreeSans 1120 0 0 0 io_in[10]
port 57 nsew signal input
flabel metal3 s 583520 453264 584800 453376 0 FreeSans 1120 0 0 0 io_in[11]
port 58 nsew signal input
flabel metal3 s 583520 497686 584800 497798 0 FreeSans 1120 0 0 0 io_in[12]
port 59 nsew signal input
flabel metal3 s 583520 587108 584800 587220 0 FreeSans 1120 0 0 0 io_in[13]
port 60 nsew signal input
flabel metal3 s -800 507984 480 508096 0 FreeSans 1120 0 0 0 io_in[14]
port 61 nsew signal input
flabel metal3 s -800 464762 480 464874 0 FreeSans 1120 0 0 0 io_in[15]
port 62 nsew signal input
flabel metal3 s -800 421540 480 421652 0 FreeSans 1120 0 0 0 io_in[16]
port 63 nsew signal input
flabel metal3 s -800 378318 480 378430 0 FreeSans 1120 0 0 0 io_in[17]
port 64 nsew signal input
flabel metal3 s -800 335096 480 335208 0 FreeSans 1120 0 0 0 io_in[18]
port 65 nsew signal input
flabel metal3 s -800 291874 480 291986 0 FreeSans 1120 0 0 0 io_in[19]
port 66 nsew signal input
flabel metal3 s 583520 7454 584800 7566 0 FreeSans 1120 0 0 0 io_in[1]
port 67 nsew signal input
flabel metal3 s -800 248852 480 248964 0 FreeSans 1120 0 0 0 io_in[20]
port 68 nsew signal input
flabel metal3 s -800 121230 480 121342 0 FreeSans 1120 0 0 0 io_in[21]
port 69 nsew signal input
flabel metal3 s -800 78008 480 78120 0 FreeSans 1120 0 0 0 io_in[22]
port 70 nsew signal input
flabel metal3 s -800 34786 480 34898 0 FreeSans 1120 0 0 0 io_in[23]
port 71 nsew signal input
flabel metal3 s -800 13364 480 13476 0 FreeSans 1120 0 0 0 io_in[24]
port 72 nsew signal input
flabel metal3 s -800 8636 480 8748 0 FreeSans 1120 0 0 0 io_in[25]
port 73 nsew signal input
flabel metal3 s -800 3908 480 4020 0 FreeSans 1120 0 0 0 io_in[26]
port 74 nsew signal input
flabel metal3 s 583520 12182 584800 12294 0 FreeSans 1120 0 0 0 io_in[2]
port 75 nsew signal input
flabel metal3 s 583520 16910 584800 17022 0 FreeSans 1120 0 0 0 io_in[3]
port 76 nsew signal input
flabel metal3 s 583520 21638 584800 21750 0 FreeSans 1120 0 0 0 io_in[4]
port 77 nsew signal input
flabel metal3 s 583520 48096 584800 48208 0 FreeSans 1120 0 0 0 io_in[5]
port 78 nsew signal input
flabel metal3 s 583520 92754 584800 92866 0 FreeSans 1120 0 0 0 io_in[6]
port 79 nsew signal input
flabel metal3 s 583520 272776 584800 272888 0 FreeSans 1120 0 0 0 io_in[7]
port 80 nsew signal input
flabel metal3 s 583520 317198 584800 317310 0 FreeSans 1120 0 0 0 io_in[8]
port 81 nsew signal input
flabel metal3 s 583520 362420 584800 362532 0 FreeSans 1120 0 0 0 io_in[9]
port 82 nsew signal input
flabel metal3 s 583520 1544 584800 1656 0 FreeSans 1120 0 0 0 io_in_3v3[0]
port 83 nsew signal input
flabel metal3 s 583520 407660 584800 407772 0 FreeSans 1120 0 0 0 io_in_3v3[10]
port 84 nsew signal input
flabel metal3 s 583520 452082 584800 452194 0 FreeSans 1120 0 0 0 io_in_3v3[11]
port 85 nsew signal input
flabel metal3 s 583520 496504 584800 496616 0 FreeSans 1120 0 0 0 io_in_3v3[12]
port 86 nsew signal input
flabel metal3 s 583520 585926 584800 586038 0 FreeSans 1120 0 0 0 io_in_3v3[13]
port 87 nsew signal input
flabel metal3 s -800 509166 480 509278 0 FreeSans 1120 0 0 0 io_in_3v3[14]
port 88 nsew signal input
flabel metal3 s -800 465944 480 466056 0 FreeSans 1120 0 0 0 io_in_3v3[15]
port 89 nsew signal input
flabel metal3 s -800 422722 480 422834 0 FreeSans 1120 0 0 0 io_in_3v3[16]
port 90 nsew signal input
flabel metal3 s -800 379500 480 379612 0 FreeSans 1120 0 0 0 io_in_3v3[17]
port 91 nsew signal input
flabel metal3 s -800 336278 480 336390 0 FreeSans 1120 0 0 0 io_in_3v3[18]
port 92 nsew signal input
flabel metal3 s -800 293056 480 293168 0 FreeSans 1120 0 0 0 io_in_3v3[19]
port 93 nsew signal input
flabel metal3 s 583520 6272 584800 6384 0 FreeSans 1120 0 0 0 io_in_3v3[1]
port 94 nsew signal input
flabel metal3 s -800 250034 480 250146 0 FreeSans 1120 0 0 0 io_in_3v3[20]
port 95 nsew signal input
flabel metal3 s -800 122412 480 122524 0 FreeSans 1120 0 0 0 io_in_3v3[21]
port 96 nsew signal input
flabel metal3 s -800 79190 480 79302 0 FreeSans 1120 0 0 0 io_in_3v3[22]
port 97 nsew signal input
flabel metal3 s -800 35968 480 36080 0 FreeSans 1120 0 0 0 io_in_3v3[23]
port 98 nsew signal input
flabel metal3 s -800 14546 480 14658 0 FreeSans 1120 0 0 0 io_in_3v3[24]
port 99 nsew signal input
flabel metal3 s -800 9818 480 9930 0 FreeSans 1120 0 0 0 io_in_3v3[25]
port 100 nsew signal input
flabel metal3 s -800 5090 480 5202 0 FreeSans 1120 0 0 0 io_in_3v3[26]
port 101 nsew signal input
flabel metal3 s 583520 11000 584800 11112 0 FreeSans 1120 0 0 0 io_in_3v3[2]
port 102 nsew signal input
flabel metal3 s 583520 15728 584800 15840 0 FreeSans 1120 0 0 0 io_in_3v3[3]
port 103 nsew signal input
flabel metal3 s 583520 20456 584800 20568 0 FreeSans 1120 0 0 0 io_in_3v3[4]
port 104 nsew signal input
flabel metal3 s 583520 46914 584800 47026 0 FreeSans 1120 0 0 0 io_in_3v3[5]
port 105 nsew signal input
flabel metal3 s 583520 91572 584800 91684 0 FreeSans 1120 0 0 0 io_in_3v3[6]
port 106 nsew signal input
flabel metal3 s 583520 271594 584800 271706 0 FreeSans 1120 0 0 0 io_in_3v3[7]
port 107 nsew signal input
flabel metal3 s 583520 316016 584800 316128 0 FreeSans 1120 0 0 0 io_in_3v3[8]
port 108 nsew signal input
flabel metal3 s 583520 361238 584800 361350 0 FreeSans 1120 0 0 0 io_in_3v3[9]
port 109 nsew signal input
flabel metal3 s 583520 5090 584800 5202 0 FreeSans 1120 0 0 0 io_oeb[0]
port 110 nsew signal tristate
flabel metal3 s 583520 411206 584800 411318 0 FreeSans 1120 0 0 0 io_oeb[10]
port 111 nsew signal tristate
flabel metal3 s 583520 455628 584800 455740 0 FreeSans 1120 0 0 0 io_oeb[11]
port 112 nsew signal tristate
flabel metal3 s 583520 500050 584800 500162 0 FreeSans 1120 0 0 0 io_oeb[12]
port 113 nsew signal tristate
flabel metal3 s 583520 589472 584800 589584 0 FreeSans 1120 0 0 0 io_oeb[13]
port 114 nsew signal tristate
flabel metal3 s -800 505620 480 505732 0 FreeSans 1120 0 0 0 io_oeb[14]
port 115 nsew signal tristate
flabel metal3 s -800 462398 480 462510 0 FreeSans 1120 0 0 0 io_oeb[15]
port 116 nsew signal tristate
flabel metal3 s -800 419176 480 419288 0 FreeSans 1120 0 0 0 io_oeb[16]
port 117 nsew signal tristate
flabel metal3 s -800 375954 480 376066 0 FreeSans 1120 0 0 0 io_oeb[17]
port 118 nsew signal tristate
flabel metal3 s -800 332732 480 332844 0 FreeSans 1120 0 0 0 io_oeb[18]
port 119 nsew signal tristate
flabel metal3 s -800 289510 480 289622 0 FreeSans 1120 0 0 0 io_oeb[19]
port 120 nsew signal tristate
flabel metal3 s 583520 9818 584800 9930 0 FreeSans 1120 0 0 0 io_oeb[1]
port 121 nsew signal tristate
flabel metal3 s -800 246488 480 246600 0 FreeSans 1120 0 0 0 io_oeb[20]
port 122 nsew signal tristate
flabel metal3 s -800 118866 480 118978 0 FreeSans 1120 0 0 0 io_oeb[21]
port 123 nsew signal tristate
flabel metal3 s -800 75644 480 75756 0 FreeSans 1120 0 0 0 io_oeb[22]
port 124 nsew signal tristate
flabel metal3 s -800 32422 480 32534 0 FreeSans 1120 0 0 0 io_oeb[23]
port 125 nsew signal tristate
flabel metal3 s -800 11000 480 11112 0 FreeSans 1120 0 0 0 io_oeb[24]
port 126 nsew signal tristate
flabel metal3 s -800 6272 480 6384 0 FreeSans 1120 0 0 0 io_oeb[25]
port 127 nsew signal tristate
flabel metal3 s -800 1544 480 1656 0 FreeSans 1120 0 0 0 io_oeb[26]
port 128 nsew signal tristate
flabel metal3 s 583520 14546 584800 14658 0 FreeSans 1120 0 0 0 io_oeb[2]
port 129 nsew signal tristate
flabel metal3 s 583520 19274 584800 19386 0 FreeSans 1120 0 0 0 io_oeb[3]
port 130 nsew signal tristate
flabel metal3 s 583520 24002 584800 24114 0 FreeSans 1120 0 0 0 io_oeb[4]
port 131 nsew signal tristate
flabel metal3 s 583520 50460 584800 50572 0 FreeSans 1120 0 0 0 io_oeb[5]
port 132 nsew signal tristate
flabel metal3 s 583520 95118 584800 95230 0 FreeSans 1120 0 0 0 io_oeb[6]
port 133 nsew signal tristate
flabel metal3 s 583520 275140 584800 275252 0 FreeSans 1120 0 0 0 io_oeb[7]
port 134 nsew signal tristate
flabel metal3 s 583520 319562 584800 319674 0 FreeSans 1120 0 0 0 io_oeb[8]
port 135 nsew signal tristate
flabel metal3 s 583520 364784 584800 364896 0 FreeSans 1120 0 0 0 io_oeb[9]
port 136 nsew signal tristate
flabel metal3 s 583520 3908 584800 4020 0 FreeSans 1120 0 0 0 io_out[0]
port 137 nsew signal tristate
flabel metal3 s 583520 410024 584800 410136 0 FreeSans 1120 0 0 0 io_out[10]
port 138 nsew signal tristate
flabel metal3 s 583520 454446 584800 454558 0 FreeSans 1120 0 0 0 io_out[11]
port 139 nsew signal tristate
flabel metal3 s 583520 498868 584800 498980 0 FreeSans 1120 0 0 0 io_out[12]
port 140 nsew signal tristate
flabel metal3 s 583520 588290 584800 588402 0 FreeSans 1120 0 0 0 io_out[13]
port 141 nsew signal tristate
flabel metal3 s -800 506802 480 506914 0 FreeSans 1120 0 0 0 io_out[14]
port 142 nsew signal tristate
flabel metal3 s -800 463580 480 463692 0 FreeSans 1120 0 0 0 io_out[15]
port 143 nsew signal tristate
flabel metal3 s -800 420358 480 420470 0 FreeSans 1120 0 0 0 io_out[16]
port 144 nsew signal tristate
flabel metal3 s -800 377136 480 377248 0 FreeSans 1120 0 0 0 io_out[17]
port 145 nsew signal tristate
flabel metal3 s -800 333914 480 334026 0 FreeSans 1120 0 0 0 io_out[18]
port 146 nsew signal tristate
flabel metal3 s -800 290692 480 290804 0 FreeSans 1120 0 0 0 io_out[19]
port 147 nsew signal tristate
flabel metal3 s 583520 8636 584800 8748 0 FreeSans 1120 0 0 0 io_out[1]
port 148 nsew signal tristate
flabel metal3 s -800 247670 480 247782 0 FreeSans 1120 0 0 0 io_out[20]
port 149 nsew signal tristate
flabel metal3 s -800 120048 480 120160 0 FreeSans 1120 0 0 0 io_out[21]
port 150 nsew signal tristate
flabel metal3 s -800 76826 480 76938 0 FreeSans 1120 0 0 0 io_out[22]
port 151 nsew signal tristate
flabel metal3 s -800 33604 480 33716 0 FreeSans 1120 0 0 0 io_out[23]
port 152 nsew signal tristate
flabel metal3 s -800 12182 480 12294 0 FreeSans 1120 0 0 0 io_out[24]
port 153 nsew signal tristate
flabel metal3 s -800 7454 480 7566 0 FreeSans 1120 0 0 0 io_out[25]
port 154 nsew signal tristate
flabel metal3 s -800 2726 480 2838 0 FreeSans 1120 0 0 0 io_out[26]
port 155 nsew signal tristate
flabel metal3 s 583520 13364 584800 13476 0 FreeSans 1120 0 0 0 io_out[2]
port 156 nsew signal tristate
flabel metal3 s 583520 18092 584800 18204 0 FreeSans 1120 0 0 0 io_out[3]
port 157 nsew signal tristate
flabel metal3 s 583520 22820 584800 22932 0 FreeSans 1120 0 0 0 io_out[4]
port 158 nsew signal tristate
flabel metal3 s 583520 49278 584800 49390 0 FreeSans 1120 0 0 0 io_out[5]
port 159 nsew signal tristate
flabel metal3 s 583520 93936 584800 94048 0 FreeSans 1120 0 0 0 io_out[6]
port 160 nsew signal tristate
flabel metal3 s 583520 273958 584800 274070 0 FreeSans 1120 0 0 0 io_out[7]
port 161 nsew signal tristate
flabel metal3 s 583520 318380 584800 318492 0 FreeSans 1120 0 0 0 io_out[8]
port 162 nsew signal tristate
flabel metal3 s 583520 363602 584800 363714 0 FreeSans 1120 0 0 0 io_out[9]
port 163 nsew signal tristate
flabel metal2 s 125816 -800 125928 480 0 FreeSans 1120 90 0 0 la_data_in[0]
port 164 nsew signal input
flabel metal2 s 480416 -800 480528 480 0 FreeSans 1120 90 0 0 la_data_in[100]
port 165 nsew signal input
flabel metal2 s 483962 -800 484074 480 0 FreeSans 1120 90 0 0 la_data_in[101]
port 166 nsew signal input
flabel metal2 s 487508 -800 487620 480 0 FreeSans 1120 90 0 0 la_data_in[102]
port 167 nsew signal input
flabel metal2 s 491054 -800 491166 480 0 FreeSans 1120 90 0 0 la_data_in[103]
port 168 nsew signal input
flabel metal2 s 494600 -800 494712 480 0 FreeSans 1120 90 0 0 la_data_in[104]
port 169 nsew signal input
flabel metal2 s 498146 -800 498258 480 0 FreeSans 1120 90 0 0 la_data_in[105]
port 170 nsew signal input
flabel metal2 s 501692 -800 501804 480 0 FreeSans 1120 90 0 0 la_data_in[106]
port 171 nsew signal input
flabel metal2 s 505238 -800 505350 480 0 FreeSans 1120 90 0 0 la_data_in[107]
port 172 nsew signal input
flabel metal2 s 508784 -800 508896 480 0 FreeSans 1120 90 0 0 la_data_in[108]
port 173 nsew signal input
flabel metal2 s 512330 -800 512442 480 0 FreeSans 1120 90 0 0 la_data_in[109]
port 174 nsew signal input
flabel metal2 s 161276 -800 161388 480 0 FreeSans 1120 90 0 0 la_data_in[10]
port 175 nsew signal input
flabel metal2 s 515876 -800 515988 480 0 FreeSans 1120 90 0 0 la_data_in[110]
port 176 nsew signal input
flabel metal2 s 519422 -800 519534 480 0 FreeSans 1120 90 0 0 la_data_in[111]
port 177 nsew signal input
flabel metal2 s 522968 -800 523080 480 0 FreeSans 1120 90 0 0 la_data_in[112]
port 178 nsew signal input
flabel metal2 s 526514 -800 526626 480 0 FreeSans 1120 90 0 0 la_data_in[113]
port 179 nsew signal input
flabel metal2 s 530060 -800 530172 480 0 FreeSans 1120 90 0 0 la_data_in[114]
port 180 nsew signal input
flabel metal2 s 533606 -800 533718 480 0 FreeSans 1120 90 0 0 la_data_in[115]
port 181 nsew signal input
flabel metal2 s 537152 -800 537264 480 0 FreeSans 1120 90 0 0 la_data_in[116]
port 182 nsew signal input
flabel metal2 s 540698 -800 540810 480 0 FreeSans 1120 90 0 0 la_data_in[117]
port 183 nsew signal input
flabel metal2 s 544244 -800 544356 480 0 FreeSans 1120 90 0 0 la_data_in[118]
port 184 nsew signal input
flabel metal2 s 547790 -800 547902 480 0 FreeSans 1120 90 0 0 la_data_in[119]
port 185 nsew signal input
flabel metal2 s 164822 -800 164934 480 0 FreeSans 1120 90 0 0 la_data_in[11]
port 186 nsew signal input
flabel metal2 s 551336 -800 551448 480 0 FreeSans 1120 90 0 0 la_data_in[120]
port 187 nsew signal input
flabel metal2 s 554882 -800 554994 480 0 FreeSans 1120 90 0 0 la_data_in[121]
port 188 nsew signal input
flabel metal2 s 558428 -800 558540 480 0 FreeSans 1120 90 0 0 la_data_in[122]
port 189 nsew signal input
flabel metal2 s 561974 -800 562086 480 0 FreeSans 1120 90 0 0 la_data_in[123]
port 190 nsew signal input
flabel metal2 s 565520 -800 565632 480 0 FreeSans 1120 90 0 0 la_data_in[124]
port 191 nsew signal input
flabel metal2 s 569066 -800 569178 480 0 FreeSans 1120 90 0 0 la_data_in[125]
port 192 nsew signal input
flabel metal2 s 572612 -800 572724 480 0 FreeSans 1120 90 0 0 la_data_in[126]
port 193 nsew signal input
flabel metal2 s 576158 -800 576270 480 0 FreeSans 1120 90 0 0 la_data_in[127]
port 194 nsew signal input
flabel metal2 s 168368 -800 168480 480 0 FreeSans 1120 90 0 0 la_data_in[12]
port 195 nsew signal input
flabel metal2 s 171914 -800 172026 480 0 FreeSans 1120 90 0 0 la_data_in[13]
port 196 nsew signal input
flabel metal2 s 175460 -800 175572 480 0 FreeSans 1120 90 0 0 la_data_in[14]
port 197 nsew signal input
flabel metal2 s 179006 -800 179118 480 0 FreeSans 1120 90 0 0 la_data_in[15]
port 198 nsew signal input
flabel metal2 s 182552 -800 182664 480 0 FreeSans 1120 90 0 0 la_data_in[16]
port 199 nsew signal input
flabel metal2 s 186098 -800 186210 480 0 FreeSans 1120 90 0 0 la_data_in[17]
port 200 nsew signal input
flabel metal2 s 189644 -800 189756 480 0 FreeSans 1120 90 0 0 la_data_in[18]
port 201 nsew signal input
flabel metal2 s 193190 -800 193302 480 0 FreeSans 1120 90 0 0 la_data_in[19]
port 202 nsew signal input
flabel metal2 s 129362 -800 129474 480 0 FreeSans 1120 90 0 0 la_data_in[1]
port 203 nsew signal input
flabel metal2 s 196736 -800 196848 480 0 FreeSans 1120 90 0 0 la_data_in[20]
port 204 nsew signal input
flabel metal2 s 200282 -800 200394 480 0 FreeSans 1120 90 0 0 la_data_in[21]
port 205 nsew signal input
flabel metal2 s 203828 -800 203940 480 0 FreeSans 1120 90 0 0 la_data_in[22]
port 206 nsew signal input
flabel metal2 s 207374 -800 207486 480 0 FreeSans 1120 90 0 0 la_data_in[23]
port 207 nsew signal input
flabel metal2 s 210920 -800 211032 480 0 FreeSans 1120 90 0 0 la_data_in[24]
port 208 nsew signal input
flabel metal2 s 214466 -800 214578 480 0 FreeSans 1120 90 0 0 la_data_in[25]
port 209 nsew signal input
flabel metal2 s 218012 -800 218124 480 0 FreeSans 1120 90 0 0 la_data_in[26]
port 210 nsew signal input
flabel metal2 s 221558 -800 221670 480 0 FreeSans 1120 90 0 0 la_data_in[27]
port 211 nsew signal input
flabel metal2 s 225104 -800 225216 480 0 FreeSans 1120 90 0 0 la_data_in[28]
port 212 nsew signal input
flabel metal2 s 228650 -800 228762 480 0 FreeSans 1120 90 0 0 la_data_in[29]
port 213 nsew signal input
flabel metal2 s 132908 -800 133020 480 0 FreeSans 1120 90 0 0 la_data_in[2]
port 214 nsew signal input
flabel metal2 s 232196 -800 232308 480 0 FreeSans 1120 90 0 0 la_data_in[30]
port 215 nsew signal input
flabel metal2 s 235742 -800 235854 480 0 FreeSans 1120 90 0 0 la_data_in[31]
port 216 nsew signal input
flabel metal2 s 239288 -800 239400 480 0 FreeSans 1120 90 0 0 la_data_in[32]
port 217 nsew signal input
flabel metal2 s 242834 -800 242946 480 0 FreeSans 1120 90 0 0 la_data_in[33]
port 218 nsew signal input
flabel metal2 s 246380 -800 246492 480 0 FreeSans 1120 90 0 0 la_data_in[34]
port 219 nsew signal input
flabel metal2 s 249926 -800 250038 480 0 FreeSans 1120 90 0 0 la_data_in[35]
port 220 nsew signal input
flabel metal2 s 253472 -800 253584 480 0 FreeSans 1120 90 0 0 la_data_in[36]
port 221 nsew signal input
flabel metal2 s 257018 -800 257130 480 0 FreeSans 1120 90 0 0 la_data_in[37]
port 222 nsew signal input
flabel metal2 s 260564 -800 260676 480 0 FreeSans 1120 90 0 0 la_data_in[38]
port 223 nsew signal input
flabel metal2 s 264110 -800 264222 480 0 FreeSans 1120 90 0 0 la_data_in[39]
port 224 nsew signal input
flabel metal2 s 136454 -800 136566 480 0 FreeSans 1120 90 0 0 la_data_in[3]
port 225 nsew signal input
flabel metal2 s 267656 -800 267768 480 0 FreeSans 1120 90 0 0 la_data_in[40]
port 226 nsew signal input
flabel metal2 s 271202 -800 271314 480 0 FreeSans 1120 90 0 0 la_data_in[41]
port 227 nsew signal input
flabel metal2 s 274748 -800 274860 480 0 FreeSans 1120 90 0 0 la_data_in[42]
port 228 nsew signal input
flabel metal2 s 278294 -800 278406 480 0 FreeSans 1120 90 0 0 la_data_in[43]
port 229 nsew signal input
flabel metal2 s 281840 -800 281952 480 0 FreeSans 1120 90 0 0 la_data_in[44]
port 230 nsew signal input
flabel metal2 s 285386 -800 285498 480 0 FreeSans 1120 90 0 0 la_data_in[45]
port 231 nsew signal input
flabel metal2 s 288932 -800 289044 480 0 FreeSans 1120 90 0 0 la_data_in[46]
port 232 nsew signal input
flabel metal2 s 292478 -800 292590 480 0 FreeSans 1120 90 0 0 la_data_in[47]
port 233 nsew signal input
flabel metal2 s 296024 -800 296136 480 0 FreeSans 1120 90 0 0 la_data_in[48]
port 234 nsew signal input
flabel metal2 s 299570 -800 299682 480 0 FreeSans 1120 90 0 0 la_data_in[49]
port 235 nsew signal input
flabel metal2 s 140000 -800 140112 480 0 FreeSans 1120 90 0 0 la_data_in[4]
port 236 nsew signal input
flabel metal2 s 303116 -800 303228 480 0 FreeSans 1120 90 0 0 la_data_in[50]
port 237 nsew signal input
flabel metal2 s 306662 -800 306774 480 0 FreeSans 1120 90 0 0 la_data_in[51]
port 238 nsew signal input
flabel metal2 s 310208 -800 310320 480 0 FreeSans 1120 90 0 0 la_data_in[52]
port 239 nsew signal input
flabel metal2 s 313754 -800 313866 480 0 FreeSans 1120 90 0 0 la_data_in[53]
port 240 nsew signal input
flabel metal2 s 317300 -800 317412 480 0 FreeSans 1120 90 0 0 la_data_in[54]
port 241 nsew signal input
flabel metal2 s 320846 -800 320958 480 0 FreeSans 1120 90 0 0 la_data_in[55]
port 242 nsew signal input
flabel metal2 s 324392 -800 324504 480 0 FreeSans 1120 90 0 0 la_data_in[56]
port 243 nsew signal input
flabel metal2 s 327938 -800 328050 480 0 FreeSans 1120 90 0 0 la_data_in[57]
port 244 nsew signal input
flabel metal2 s 331484 -800 331596 480 0 FreeSans 1120 90 0 0 la_data_in[58]
port 245 nsew signal input
flabel metal2 s 335030 -800 335142 480 0 FreeSans 1120 90 0 0 la_data_in[59]
port 246 nsew signal input
flabel metal2 s 143546 -800 143658 480 0 FreeSans 1120 90 0 0 la_data_in[5]
port 247 nsew signal input
flabel metal2 s 338576 -800 338688 480 0 FreeSans 1120 90 0 0 la_data_in[60]
port 248 nsew signal input
flabel metal2 s 342122 -800 342234 480 0 FreeSans 1120 90 0 0 la_data_in[61]
port 249 nsew signal input
flabel metal2 s 345668 -800 345780 480 0 FreeSans 1120 90 0 0 la_data_in[62]
port 250 nsew signal input
flabel metal2 s 349214 -800 349326 480 0 FreeSans 1120 90 0 0 la_data_in[63]
port 251 nsew signal input
flabel metal2 s 352760 -800 352872 480 0 FreeSans 1120 90 0 0 la_data_in[64]
port 252 nsew signal input
flabel metal2 s 356306 -800 356418 480 0 FreeSans 1120 90 0 0 la_data_in[65]
port 253 nsew signal input
flabel metal2 s 359852 -800 359964 480 0 FreeSans 1120 90 0 0 la_data_in[66]
port 254 nsew signal input
flabel metal2 s 363398 -800 363510 480 0 FreeSans 1120 90 0 0 la_data_in[67]
port 255 nsew signal input
flabel metal2 s 366944 -800 367056 480 0 FreeSans 1120 90 0 0 la_data_in[68]
port 256 nsew signal input
flabel metal2 s 370490 -800 370602 480 0 FreeSans 1120 90 0 0 la_data_in[69]
port 257 nsew signal input
flabel metal2 s 147092 -800 147204 480 0 FreeSans 1120 90 0 0 la_data_in[6]
port 258 nsew signal input
flabel metal2 s 374036 -800 374148 480 0 FreeSans 1120 90 0 0 la_data_in[70]
port 259 nsew signal input
flabel metal2 s 377582 -800 377694 480 0 FreeSans 1120 90 0 0 la_data_in[71]
port 260 nsew signal input
flabel metal2 s 381128 -800 381240 480 0 FreeSans 1120 90 0 0 la_data_in[72]
port 261 nsew signal input
flabel metal2 s 384674 -800 384786 480 0 FreeSans 1120 90 0 0 la_data_in[73]
port 262 nsew signal input
flabel metal2 s 388220 -800 388332 480 0 FreeSans 1120 90 0 0 la_data_in[74]
port 263 nsew signal input
flabel metal2 s 391766 -800 391878 480 0 FreeSans 1120 90 0 0 la_data_in[75]
port 264 nsew signal input
flabel metal2 s 395312 -800 395424 480 0 FreeSans 1120 90 0 0 la_data_in[76]
port 265 nsew signal input
flabel metal2 s 398858 -800 398970 480 0 FreeSans 1120 90 0 0 la_data_in[77]
port 266 nsew signal input
flabel metal2 s 402404 -800 402516 480 0 FreeSans 1120 90 0 0 la_data_in[78]
port 267 nsew signal input
flabel metal2 s 405950 -800 406062 480 0 FreeSans 1120 90 0 0 la_data_in[79]
port 268 nsew signal input
flabel metal2 s 150638 -800 150750 480 0 FreeSans 1120 90 0 0 la_data_in[7]
port 269 nsew signal input
flabel metal2 s 409496 -800 409608 480 0 FreeSans 1120 90 0 0 la_data_in[80]
port 270 nsew signal input
flabel metal2 s 413042 -800 413154 480 0 FreeSans 1120 90 0 0 la_data_in[81]
port 271 nsew signal input
flabel metal2 s 416588 -800 416700 480 0 FreeSans 1120 90 0 0 la_data_in[82]
port 272 nsew signal input
flabel metal2 s 420134 -800 420246 480 0 FreeSans 1120 90 0 0 la_data_in[83]
port 273 nsew signal input
flabel metal2 s 423680 -800 423792 480 0 FreeSans 1120 90 0 0 la_data_in[84]
port 274 nsew signal input
flabel metal2 s 427226 -800 427338 480 0 FreeSans 1120 90 0 0 la_data_in[85]
port 275 nsew signal input
flabel metal2 s 430772 -800 430884 480 0 FreeSans 1120 90 0 0 la_data_in[86]
port 276 nsew signal input
flabel metal2 s 434318 -800 434430 480 0 FreeSans 1120 90 0 0 la_data_in[87]
port 277 nsew signal input
flabel metal2 s 437864 -800 437976 480 0 FreeSans 1120 90 0 0 la_data_in[88]
port 278 nsew signal input
flabel metal2 s 441410 -800 441522 480 0 FreeSans 1120 90 0 0 la_data_in[89]
port 279 nsew signal input
flabel metal2 s 154184 -800 154296 480 0 FreeSans 1120 90 0 0 la_data_in[8]
port 280 nsew signal input
flabel metal2 s 444956 -800 445068 480 0 FreeSans 1120 90 0 0 la_data_in[90]
port 281 nsew signal input
flabel metal2 s 448502 -800 448614 480 0 FreeSans 1120 90 0 0 la_data_in[91]
port 282 nsew signal input
flabel metal2 s 452048 -800 452160 480 0 FreeSans 1120 90 0 0 la_data_in[92]
port 283 nsew signal input
flabel metal2 s 455594 -800 455706 480 0 FreeSans 1120 90 0 0 la_data_in[93]
port 284 nsew signal input
flabel metal2 s 459140 -800 459252 480 0 FreeSans 1120 90 0 0 la_data_in[94]
port 285 nsew signal input
flabel metal2 s 462686 -800 462798 480 0 FreeSans 1120 90 0 0 la_data_in[95]
port 286 nsew signal input
flabel metal2 s 466232 -800 466344 480 0 FreeSans 1120 90 0 0 la_data_in[96]
port 287 nsew signal input
flabel metal2 s 469778 -800 469890 480 0 FreeSans 1120 90 0 0 la_data_in[97]
port 288 nsew signal input
flabel metal2 s 473324 -800 473436 480 0 FreeSans 1120 90 0 0 la_data_in[98]
port 289 nsew signal input
flabel metal2 s 476870 -800 476982 480 0 FreeSans 1120 90 0 0 la_data_in[99]
port 290 nsew signal input
flabel metal2 s 157730 -800 157842 480 0 FreeSans 1120 90 0 0 la_data_in[9]
port 291 nsew signal input
flabel metal2 s 126998 -800 127110 480 0 FreeSans 1120 90 0 0 la_data_out[0]
port 292 nsew signal tristate
flabel metal2 s 481598 -800 481710 480 0 FreeSans 1120 90 0 0 la_data_out[100]
port 293 nsew signal tristate
flabel metal2 s 485144 -800 485256 480 0 FreeSans 1120 90 0 0 la_data_out[101]
port 294 nsew signal tristate
flabel metal2 s 488690 -800 488802 480 0 FreeSans 1120 90 0 0 la_data_out[102]
port 295 nsew signal tristate
flabel metal2 s 492236 -800 492348 480 0 FreeSans 1120 90 0 0 la_data_out[103]
port 296 nsew signal tristate
flabel metal2 s 495782 -800 495894 480 0 FreeSans 1120 90 0 0 la_data_out[104]
port 297 nsew signal tristate
flabel metal2 s 499328 -800 499440 480 0 FreeSans 1120 90 0 0 la_data_out[105]
port 298 nsew signal tristate
flabel metal2 s 502874 -800 502986 480 0 FreeSans 1120 90 0 0 la_data_out[106]
port 299 nsew signal tristate
flabel metal2 s 506420 -800 506532 480 0 FreeSans 1120 90 0 0 la_data_out[107]
port 300 nsew signal tristate
flabel metal2 s 509966 -800 510078 480 0 FreeSans 1120 90 0 0 la_data_out[108]
port 301 nsew signal tristate
flabel metal2 s 513512 -800 513624 480 0 FreeSans 1120 90 0 0 la_data_out[109]
port 302 nsew signal tristate
flabel metal2 s 162458 -800 162570 480 0 FreeSans 1120 90 0 0 la_data_out[10]
port 303 nsew signal tristate
flabel metal2 s 517058 -800 517170 480 0 FreeSans 1120 90 0 0 la_data_out[110]
port 304 nsew signal tristate
flabel metal2 s 520604 -800 520716 480 0 FreeSans 1120 90 0 0 la_data_out[111]
port 305 nsew signal tristate
flabel metal2 s 524150 -800 524262 480 0 FreeSans 1120 90 0 0 la_data_out[112]
port 306 nsew signal tristate
flabel metal2 s 527696 -800 527808 480 0 FreeSans 1120 90 0 0 la_data_out[113]
port 307 nsew signal tristate
flabel metal2 s 531242 -800 531354 480 0 FreeSans 1120 90 0 0 la_data_out[114]
port 308 nsew signal tristate
flabel metal2 s 534788 -800 534900 480 0 FreeSans 1120 90 0 0 la_data_out[115]
port 309 nsew signal tristate
flabel metal2 s 538334 -800 538446 480 0 FreeSans 1120 90 0 0 la_data_out[116]
port 310 nsew signal tristate
flabel metal2 s 541880 -800 541992 480 0 FreeSans 1120 90 0 0 la_data_out[117]
port 311 nsew signal tristate
flabel metal2 s 545426 -800 545538 480 0 FreeSans 1120 90 0 0 la_data_out[118]
port 312 nsew signal tristate
flabel metal2 s 548972 -800 549084 480 0 FreeSans 1120 90 0 0 la_data_out[119]
port 313 nsew signal tristate
flabel metal2 s 166004 -800 166116 480 0 FreeSans 1120 90 0 0 la_data_out[11]
port 314 nsew signal tristate
flabel metal2 s 552518 -800 552630 480 0 FreeSans 1120 90 0 0 la_data_out[120]
port 315 nsew signal tristate
flabel metal2 s 556064 -800 556176 480 0 FreeSans 1120 90 0 0 la_data_out[121]
port 316 nsew signal tristate
flabel metal2 s 559610 -800 559722 480 0 FreeSans 1120 90 0 0 la_data_out[122]
port 317 nsew signal tristate
flabel metal2 s 563156 -800 563268 480 0 FreeSans 1120 90 0 0 la_data_out[123]
port 318 nsew signal tristate
flabel metal2 s 566702 -800 566814 480 0 FreeSans 1120 90 0 0 la_data_out[124]
port 319 nsew signal tristate
flabel metal2 s 570248 -800 570360 480 0 FreeSans 1120 90 0 0 la_data_out[125]
port 320 nsew signal tristate
flabel metal2 s 573794 -800 573906 480 0 FreeSans 1120 90 0 0 la_data_out[126]
port 321 nsew signal tristate
flabel metal2 s 577340 -800 577452 480 0 FreeSans 1120 90 0 0 la_data_out[127]
port 322 nsew signal tristate
flabel metal2 s 169550 -800 169662 480 0 FreeSans 1120 90 0 0 la_data_out[12]
port 323 nsew signal tristate
flabel metal2 s 173096 -800 173208 480 0 FreeSans 1120 90 0 0 la_data_out[13]
port 324 nsew signal tristate
flabel metal2 s 176642 -800 176754 480 0 FreeSans 1120 90 0 0 la_data_out[14]
port 325 nsew signal tristate
flabel metal2 s 180188 -800 180300 480 0 FreeSans 1120 90 0 0 la_data_out[15]
port 326 nsew signal tristate
flabel metal2 s 183734 -800 183846 480 0 FreeSans 1120 90 0 0 la_data_out[16]
port 327 nsew signal tristate
flabel metal2 s 187280 -800 187392 480 0 FreeSans 1120 90 0 0 la_data_out[17]
port 328 nsew signal tristate
flabel metal2 s 190826 -800 190938 480 0 FreeSans 1120 90 0 0 la_data_out[18]
port 329 nsew signal tristate
flabel metal2 s 194372 -800 194484 480 0 FreeSans 1120 90 0 0 la_data_out[19]
port 330 nsew signal tristate
flabel metal2 s 130544 -800 130656 480 0 FreeSans 1120 90 0 0 la_data_out[1]
port 331 nsew signal tristate
flabel metal2 s 197918 -800 198030 480 0 FreeSans 1120 90 0 0 la_data_out[20]
port 332 nsew signal tristate
flabel metal2 s 201464 -800 201576 480 0 FreeSans 1120 90 0 0 la_data_out[21]
port 333 nsew signal tristate
flabel metal2 s 205010 -800 205122 480 0 FreeSans 1120 90 0 0 la_data_out[22]
port 334 nsew signal tristate
flabel metal2 s 208556 -800 208668 480 0 FreeSans 1120 90 0 0 la_data_out[23]
port 335 nsew signal tristate
flabel metal2 s 212102 -800 212214 480 0 FreeSans 1120 90 0 0 la_data_out[24]
port 336 nsew signal tristate
flabel metal2 s 215648 -800 215760 480 0 FreeSans 1120 90 0 0 la_data_out[25]
port 337 nsew signal tristate
flabel metal2 s 219194 -800 219306 480 0 FreeSans 1120 90 0 0 la_data_out[26]
port 338 nsew signal tristate
flabel metal2 s 222740 -800 222852 480 0 FreeSans 1120 90 0 0 la_data_out[27]
port 339 nsew signal tristate
flabel metal2 s 226286 -800 226398 480 0 FreeSans 1120 90 0 0 la_data_out[28]
port 340 nsew signal tristate
flabel metal2 s 229832 -800 229944 480 0 FreeSans 1120 90 0 0 la_data_out[29]
port 341 nsew signal tristate
flabel metal2 s 134090 -800 134202 480 0 FreeSans 1120 90 0 0 la_data_out[2]
port 342 nsew signal tristate
flabel metal2 s 233378 -800 233490 480 0 FreeSans 1120 90 0 0 la_data_out[30]
port 343 nsew signal tristate
flabel metal2 s 236924 -800 237036 480 0 FreeSans 1120 90 0 0 la_data_out[31]
port 344 nsew signal tristate
flabel metal2 s 240470 -800 240582 480 0 FreeSans 1120 90 0 0 la_data_out[32]
port 345 nsew signal tristate
flabel metal2 s 244016 -800 244128 480 0 FreeSans 1120 90 0 0 la_data_out[33]
port 346 nsew signal tristate
flabel metal2 s 247562 -800 247674 480 0 FreeSans 1120 90 0 0 la_data_out[34]
port 347 nsew signal tristate
flabel metal2 s 251108 -800 251220 480 0 FreeSans 1120 90 0 0 la_data_out[35]
port 348 nsew signal tristate
flabel metal2 s 254654 -800 254766 480 0 FreeSans 1120 90 0 0 la_data_out[36]
port 349 nsew signal tristate
flabel metal2 s 258200 -800 258312 480 0 FreeSans 1120 90 0 0 la_data_out[37]
port 350 nsew signal tristate
flabel metal2 s 261746 -800 261858 480 0 FreeSans 1120 90 0 0 la_data_out[38]
port 351 nsew signal tristate
flabel metal2 s 265292 -800 265404 480 0 FreeSans 1120 90 0 0 la_data_out[39]
port 352 nsew signal tristate
flabel metal2 s 137636 -800 137748 480 0 FreeSans 1120 90 0 0 la_data_out[3]
port 353 nsew signal tristate
flabel metal2 s 268838 -800 268950 480 0 FreeSans 1120 90 0 0 la_data_out[40]
port 354 nsew signal tristate
flabel metal2 s 272384 -800 272496 480 0 FreeSans 1120 90 0 0 la_data_out[41]
port 355 nsew signal tristate
flabel metal2 s 275930 -800 276042 480 0 FreeSans 1120 90 0 0 la_data_out[42]
port 356 nsew signal tristate
flabel metal2 s 279476 -800 279588 480 0 FreeSans 1120 90 0 0 la_data_out[43]
port 357 nsew signal tristate
flabel metal2 s 283022 -800 283134 480 0 FreeSans 1120 90 0 0 la_data_out[44]
port 358 nsew signal tristate
flabel metal2 s 286568 -800 286680 480 0 FreeSans 1120 90 0 0 la_data_out[45]
port 359 nsew signal tristate
flabel metal2 s 290114 -800 290226 480 0 FreeSans 1120 90 0 0 la_data_out[46]
port 360 nsew signal tristate
flabel metal2 s 293660 -800 293772 480 0 FreeSans 1120 90 0 0 la_data_out[47]
port 361 nsew signal tristate
flabel metal2 s 297206 -800 297318 480 0 FreeSans 1120 90 0 0 la_data_out[48]
port 362 nsew signal tristate
flabel metal2 s 300752 -800 300864 480 0 FreeSans 1120 90 0 0 la_data_out[49]
port 363 nsew signal tristate
flabel metal2 s 141182 -800 141294 480 0 FreeSans 1120 90 0 0 la_data_out[4]
port 364 nsew signal tristate
flabel metal2 s 304298 -800 304410 480 0 FreeSans 1120 90 0 0 la_data_out[50]
port 365 nsew signal tristate
flabel metal2 s 307844 -800 307956 480 0 FreeSans 1120 90 0 0 la_data_out[51]
port 366 nsew signal tristate
flabel metal2 s 311390 -800 311502 480 0 FreeSans 1120 90 0 0 la_data_out[52]
port 367 nsew signal tristate
flabel metal2 s 314936 -800 315048 480 0 FreeSans 1120 90 0 0 la_data_out[53]
port 368 nsew signal tristate
flabel metal2 s 318482 -800 318594 480 0 FreeSans 1120 90 0 0 la_data_out[54]
port 369 nsew signal tristate
flabel metal2 s 322028 -800 322140 480 0 FreeSans 1120 90 0 0 la_data_out[55]
port 370 nsew signal tristate
flabel metal2 s 325574 -800 325686 480 0 FreeSans 1120 90 0 0 la_data_out[56]
port 371 nsew signal tristate
flabel metal2 s 329120 -800 329232 480 0 FreeSans 1120 90 0 0 la_data_out[57]
port 372 nsew signal tristate
flabel metal2 s 332666 -800 332778 480 0 FreeSans 1120 90 0 0 la_data_out[58]
port 373 nsew signal tristate
flabel metal2 s 336212 -800 336324 480 0 FreeSans 1120 90 0 0 la_data_out[59]
port 374 nsew signal tristate
flabel metal2 s 144728 -800 144840 480 0 FreeSans 1120 90 0 0 la_data_out[5]
port 375 nsew signal tristate
flabel metal2 s 339758 -800 339870 480 0 FreeSans 1120 90 0 0 la_data_out[60]
port 376 nsew signal tristate
flabel metal2 s 343304 -800 343416 480 0 FreeSans 1120 90 0 0 la_data_out[61]
port 377 nsew signal tristate
flabel metal2 s 346850 -800 346962 480 0 FreeSans 1120 90 0 0 la_data_out[62]
port 378 nsew signal tristate
flabel metal2 s 350396 -800 350508 480 0 FreeSans 1120 90 0 0 la_data_out[63]
port 379 nsew signal tristate
flabel metal2 s 353942 -800 354054 480 0 FreeSans 1120 90 0 0 la_data_out[64]
port 380 nsew signal tristate
flabel metal2 s 357488 -800 357600 480 0 FreeSans 1120 90 0 0 la_data_out[65]
port 381 nsew signal tristate
flabel metal2 s 361034 -800 361146 480 0 FreeSans 1120 90 0 0 la_data_out[66]
port 382 nsew signal tristate
flabel metal2 s 364580 -800 364692 480 0 FreeSans 1120 90 0 0 la_data_out[67]
port 383 nsew signal tristate
flabel metal2 s 368126 -800 368238 480 0 FreeSans 1120 90 0 0 la_data_out[68]
port 384 nsew signal tristate
flabel metal2 s 371672 -800 371784 480 0 FreeSans 1120 90 0 0 la_data_out[69]
port 385 nsew signal tristate
flabel metal2 s 148274 -800 148386 480 0 FreeSans 1120 90 0 0 la_data_out[6]
port 386 nsew signal tristate
flabel metal2 s 375218 -800 375330 480 0 FreeSans 1120 90 0 0 la_data_out[70]
port 387 nsew signal tristate
flabel metal2 s 378764 -800 378876 480 0 FreeSans 1120 90 0 0 la_data_out[71]
port 388 nsew signal tristate
flabel metal2 s 382310 -800 382422 480 0 FreeSans 1120 90 0 0 la_data_out[72]
port 389 nsew signal tristate
flabel metal2 s 385856 -800 385968 480 0 FreeSans 1120 90 0 0 la_data_out[73]
port 390 nsew signal tristate
flabel metal2 s 389402 -800 389514 480 0 FreeSans 1120 90 0 0 la_data_out[74]
port 391 nsew signal tristate
flabel metal2 s 392948 -800 393060 480 0 FreeSans 1120 90 0 0 la_data_out[75]
port 392 nsew signal tristate
flabel metal2 s 396494 -800 396606 480 0 FreeSans 1120 90 0 0 la_data_out[76]
port 393 nsew signal tristate
flabel metal2 s 400040 -800 400152 480 0 FreeSans 1120 90 0 0 la_data_out[77]
port 394 nsew signal tristate
flabel metal2 s 403586 -800 403698 480 0 FreeSans 1120 90 0 0 la_data_out[78]
port 395 nsew signal tristate
flabel metal2 s 407132 -800 407244 480 0 FreeSans 1120 90 0 0 la_data_out[79]
port 396 nsew signal tristate
flabel metal2 s 151820 -800 151932 480 0 FreeSans 1120 90 0 0 la_data_out[7]
port 397 nsew signal tristate
flabel metal2 s 410678 -800 410790 480 0 FreeSans 1120 90 0 0 la_data_out[80]
port 398 nsew signal tristate
flabel metal2 s 414224 -800 414336 480 0 FreeSans 1120 90 0 0 la_data_out[81]
port 399 nsew signal tristate
flabel metal2 s 417770 -800 417882 480 0 FreeSans 1120 90 0 0 la_data_out[82]
port 400 nsew signal tristate
flabel metal2 s 421316 -800 421428 480 0 FreeSans 1120 90 0 0 la_data_out[83]
port 401 nsew signal tristate
flabel metal2 s 424862 -800 424974 480 0 FreeSans 1120 90 0 0 la_data_out[84]
port 402 nsew signal tristate
flabel metal2 s 428408 -800 428520 480 0 FreeSans 1120 90 0 0 la_data_out[85]
port 403 nsew signal tristate
flabel metal2 s 431954 -800 432066 480 0 FreeSans 1120 90 0 0 la_data_out[86]
port 404 nsew signal tristate
flabel metal2 s 435500 -800 435612 480 0 FreeSans 1120 90 0 0 la_data_out[87]
port 405 nsew signal tristate
flabel metal2 s 439046 -800 439158 480 0 FreeSans 1120 90 0 0 la_data_out[88]
port 406 nsew signal tristate
flabel metal2 s 442592 -800 442704 480 0 FreeSans 1120 90 0 0 la_data_out[89]
port 407 nsew signal tristate
flabel metal2 s 155366 -800 155478 480 0 FreeSans 1120 90 0 0 la_data_out[8]
port 408 nsew signal tristate
flabel metal2 s 446138 -800 446250 480 0 FreeSans 1120 90 0 0 la_data_out[90]
port 409 nsew signal tristate
flabel metal2 s 449684 -800 449796 480 0 FreeSans 1120 90 0 0 la_data_out[91]
port 410 nsew signal tristate
flabel metal2 s 453230 -800 453342 480 0 FreeSans 1120 90 0 0 la_data_out[92]
port 411 nsew signal tristate
flabel metal2 s 456776 -800 456888 480 0 FreeSans 1120 90 0 0 la_data_out[93]
port 412 nsew signal tristate
flabel metal2 s 460322 -800 460434 480 0 FreeSans 1120 90 0 0 la_data_out[94]
port 413 nsew signal tristate
flabel metal2 s 463868 -800 463980 480 0 FreeSans 1120 90 0 0 la_data_out[95]
port 414 nsew signal tristate
flabel metal2 s 467414 -800 467526 480 0 FreeSans 1120 90 0 0 la_data_out[96]
port 415 nsew signal tristate
flabel metal2 s 470960 -800 471072 480 0 FreeSans 1120 90 0 0 la_data_out[97]
port 416 nsew signal tristate
flabel metal2 s 474506 -800 474618 480 0 FreeSans 1120 90 0 0 la_data_out[98]
port 417 nsew signal tristate
flabel metal2 s 478052 -800 478164 480 0 FreeSans 1120 90 0 0 la_data_out[99]
port 418 nsew signal tristate
flabel metal2 s 158912 -800 159024 480 0 FreeSans 1120 90 0 0 la_data_out[9]
port 419 nsew signal tristate
flabel metal2 s 128180 -800 128292 480 0 FreeSans 1120 90 0 0 la_oenb[0]
port 420 nsew signal input
flabel metal2 s 482780 -800 482892 480 0 FreeSans 1120 90 0 0 la_oenb[100]
port 421 nsew signal input
flabel metal2 s 486326 -800 486438 480 0 FreeSans 1120 90 0 0 la_oenb[101]
port 422 nsew signal input
flabel metal2 s 489872 -800 489984 480 0 FreeSans 1120 90 0 0 la_oenb[102]
port 423 nsew signal input
flabel metal2 s 493418 -800 493530 480 0 FreeSans 1120 90 0 0 la_oenb[103]
port 424 nsew signal input
flabel metal2 s 496964 -800 497076 480 0 FreeSans 1120 90 0 0 la_oenb[104]
port 425 nsew signal input
flabel metal2 s 500510 -800 500622 480 0 FreeSans 1120 90 0 0 la_oenb[105]
port 426 nsew signal input
flabel metal2 s 504056 -800 504168 480 0 FreeSans 1120 90 0 0 la_oenb[106]
port 427 nsew signal input
flabel metal2 s 507602 -800 507714 480 0 FreeSans 1120 90 0 0 la_oenb[107]
port 428 nsew signal input
flabel metal2 s 511148 -800 511260 480 0 FreeSans 1120 90 0 0 la_oenb[108]
port 429 nsew signal input
flabel metal2 s 514694 -800 514806 480 0 FreeSans 1120 90 0 0 la_oenb[109]
port 430 nsew signal input
flabel metal2 s 163640 -800 163752 480 0 FreeSans 1120 90 0 0 la_oenb[10]
port 431 nsew signal input
flabel metal2 s 518240 -800 518352 480 0 FreeSans 1120 90 0 0 la_oenb[110]
port 432 nsew signal input
flabel metal2 s 521786 -800 521898 480 0 FreeSans 1120 90 0 0 la_oenb[111]
port 433 nsew signal input
flabel metal2 s 525332 -800 525444 480 0 FreeSans 1120 90 0 0 la_oenb[112]
port 434 nsew signal input
flabel metal2 s 528878 -800 528990 480 0 FreeSans 1120 90 0 0 la_oenb[113]
port 435 nsew signal input
flabel metal2 s 532424 -800 532536 480 0 FreeSans 1120 90 0 0 la_oenb[114]
port 436 nsew signal input
flabel metal2 s 535970 -800 536082 480 0 FreeSans 1120 90 0 0 la_oenb[115]
port 437 nsew signal input
flabel metal2 s 539516 -800 539628 480 0 FreeSans 1120 90 0 0 la_oenb[116]
port 438 nsew signal input
flabel metal2 s 543062 -800 543174 480 0 FreeSans 1120 90 0 0 la_oenb[117]
port 439 nsew signal input
flabel metal2 s 546608 -800 546720 480 0 FreeSans 1120 90 0 0 la_oenb[118]
port 440 nsew signal input
flabel metal2 s 550154 -800 550266 480 0 FreeSans 1120 90 0 0 la_oenb[119]
port 441 nsew signal input
flabel metal2 s 167186 -800 167298 480 0 FreeSans 1120 90 0 0 la_oenb[11]
port 442 nsew signal input
flabel metal2 s 553700 -800 553812 480 0 FreeSans 1120 90 0 0 la_oenb[120]
port 443 nsew signal input
flabel metal2 s 557246 -800 557358 480 0 FreeSans 1120 90 0 0 la_oenb[121]
port 444 nsew signal input
flabel metal2 s 560792 -800 560904 480 0 FreeSans 1120 90 0 0 la_oenb[122]
port 445 nsew signal input
flabel metal2 s 564338 -800 564450 480 0 FreeSans 1120 90 0 0 la_oenb[123]
port 446 nsew signal input
flabel metal2 s 567884 -800 567996 480 0 FreeSans 1120 90 0 0 la_oenb[124]
port 447 nsew signal input
flabel metal2 s 571430 -800 571542 480 0 FreeSans 1120 90 0 0 la_oenb[125]
port 448 nsew signal input
flabel metal2 s 574976 -800 575088 480 0 FreeSans 1120 90 0 0 la_oenb[126]
port 449 nsew signal input
flabel metal2 s 578522 -800 578634 480 0 FreeSans 1120 90 0 0 la_oenb[127]
port 450 nsew signal input
flabel metal2 s 170732 -800 170844 480 0 FreeSans 1120 90 0 0 la_oenb[12]
port 451 nsew signal input
flabel metal2 s 174278 -800 174390 480 0 FreeSans 1120 90 0 0 la_oenb[13]
port 452 nsew signal input
flabel metal2 s 177824 -800 177936 480 0 FreeSans 1120 90 0 0 la_oenb[14]
port 453 nsew signal input
flabel metal2 s 181370 -800 181482 480 0 FreeSans 1120 90 0 0 la_oenb[15]
port 454 nsew signal input
flabel metal2 s 184916 -800 185028 480 0 FreeSans 1120 90 0 0 la_oenb[16]
port 455 nsew signal input
flabel metal2 s 188462 -800 188574 480 0 FreeSans 1120 90 0 0 la_oenb[17]
port 456 nsew signal input
flabel metal2 s 192008 -800 192120 480 0 FreeSans 1120 90 0 0 la_oenb[18]
port 457 nsew signal input
flabel metal2 s 195554 -800 195666 480 0 FreeSans 1120 90 0 0 la_oenb[19]
port 458 nsew signal input
flabel metal2 s 131726 -800 131838 480 0 FreeSans 1120 90 0 0 la_oenb[1]
port 459 nsew signal input
flabel metal2 s 199100 -800 199212 480 0 FreeSans 1120 90 0 0 la_oenb[20]
port 460 nsew signal input
flabel metal2 s 202646 -800 202758 480 0 FreeSans 1120 90 0 0 la_oenb[21]
port 461 nsew signal input
flabel metal2 s 206192 -800 206304 480 0 FreeSans 1120 90 0 0 la_oenb[22]
port 462 nsew signal input
flabel metal2 s 209738 -800 209850 480 0 FreeSans 1120 90 0 0 la_oenb[23]
port 463 nsew signal input
flabel metal2 s 213284 -800 213396 480 0 FreeSans 1120 90 0 0 la_oenb[24]
port 464 nsew signal input
flabel metal2 s 216830 -800 216942 480 0 FreeSans 1120 90 0 0 la_oenb[25]
port 465 nsew signal input
flabel metal2 s 220376 -800 220488 480 0 FreeSans 1120 90 0 0 la_oenb[26]
port 466 nsew signal input
flabel metal2 s 223922 -800 224034 480 0 FreeSans 1120 90 0 0 la_oenb[27]
port 467 nsew signal input
flabel metal2 s 227468 -800 227580 480 0 FreeSans 1120 90 0 0 la_oenb[28]
port 468 nsew signal input
flabel metal2 s 231014 -800 231126 480 0 FreeSans 1120 90 0 0 la_oenb[29]
port 469 nsew signal input
flabel metal2 s 135272 -800 135384 480 0 FreeSans 1120 90 0 0 la_oenb[2]
port 470 nsew signal input
flabel metal2 s 234560 -800 234672 480 0 FreeSans 1120 90 0 0 la_oenb[30]
port 471 nsew signal input
flabel metal2 s 238106 -800 238218 480 0 FreeSans 1120 90 0 0 la_oenb[31]
port 472 nsew signal input
flabel metal2 s 241652 -800 241764 480 0 FreeSans 1120 90 0 0 la_oenb[32]
port 473 nsew signal input
flabel metal2 s 245198 -800 245310 480 0 FreeSans 1120 90 0 0 la_oenb[33]
port 474 nsew signal input
flabel metal2 s 248744 -800 248856 480 0 FreeSans 1120 90 0 0 la_oenb[34]
port 475 nsew signal input
flabel metal2 s 252290 -800 252402 480 0 FreeSans 1120 90 0 0 la_oenb[35]
port 476 nsew signal input
flabel metal2 s 255836 -800 255948 480 0 FreeSans 1120 90 0 0 la_oenb[36]
port 477 nsew signal input
flabel metal2 s 259382 -800 259494 480 0 FreeSans 1120 90 0 0 la_oenb[37]
port 478 nsew signal input
flabel metal2 s 262928 -800 263040 480 0 FreeSans 1120 90 0 0 la_oenb[38]
port 479 nsew signal input
flabel metal2 s 266474 -800 266586 480 0 FreeSans 1120 90 0 0 la_oenb[39]
port 480 nsew signal input
flabel metal2 s 138818 -800 138930 480 0 FreeSans 1120 90 0 0 la_oenb[3]
port 481 nsew signal input
flabel metal2 s 270020 -800 270132 480 0 FreeSans 1120 90 0 0 la_oenb[40]
port 482 nsew signal input
flabel metal2 s 273566 -800 273678 480 0 FreeSans 1120 90 0 0 la_oenb[41]
port 483 nsew signal input
flabel metal2 s 277112 -800 277224 480 0 FreeSans 1120 90 0 0 la_oenb[42]
port 484 nsew signal input
flabel metal2 s 280658 -800 280770 480 0 FreeSans 1120 90 0 0 la_oenb[43]
port 485 nsew signal input
flabel metal2 s 284204 -800 284316 480 0 FreeSans 1120 90 0 0 la_oenb[44]
port 486 nsew signal input
flabel metal2 s 287750 -800 287862 480 0 FreeSans 1120 90 0 0 la_oenb[45]
port 487 nsew signal input
flabel metal2 s 291296 -800 291408 480 0 FreeSans 1120 90 0 0 la_oenb[46]
port 488 nsew signal input
flabel metal2 s 294842 -800 294954 480 0 FreeSans 1120 90 0 0 la_oenb[47]
port 489 nsew signal input
flabel metal2 s 298388 -800 298500 480 0 FreeSans 1120 90 0 0 la_oenb[48]
port 490 nsew signal input
flabel metal2 s 301934 -800 302046 480 0 FreeSans 1120 90 0 0 la_oenb[49]
port 491 nsew signal input
flabel metal2 s 142364 -800 142476 480 0 FreeSans 1120 90 0 0 la_oenb[4]
port 492 nsew signal input
flabel metal2 s 305480 -800 305592 480 0 FreeSans 1120 90 0 0 la_oenb[50]
port 493 nsew signal input
flabel metal2 s 309026 -800 309138 480 0 FreeSans 1120 90 0 0 la_oenb[51]
port 494 nsew signal input
flabel metal2 s 312572 -800 312684 480 0 FreeSans 1120 90 0 0 la_oenb[52]
port 495 nsew signal input
flabel metal2 s 316118 -800 316230 480 0 FreeSans 1120 90 0 0 la_oenb[53]
port 496 nsew signal input
flabel metal2 s 319664 -800 319776 480 0 FreeSans 1120 90 0 0 la_oenb[54]
port 497 nsew signal input
flabel metal2 s 323210 -800 323322 480 0 FreeSans 1120 90 0 0 la_oenb[55]
port 498 nsew signal input
flabel metal2 s 326756 -800 326868 480 0 FreeSans 1120 90 0 0 la_oenb[56]
port 499 nsew signal input
flabel metal2 s 330302 -800 330414 480 0 FreeSans 1120 90 0 0 la_oenb[57]
port 500 nsew signal input
flabel metal2 s 333848 -800 333960 480 0 FreeSans 1120 90 0 0 la_oenb[58]
port 501 nsew signal input
flabel metal2 s 337394 -800 337506 480 0 FreeSans 1120 90 0 0 la_oenb[59]
port 502 nsew signal input
flabel metal2 s 145910 -800 146022 480 0 FreeSans 1120 90 0 0 la_oenb[5]
port 503 nsew signal input
flabel metal2 s 340940 -800 341052 480 0 FreeSans 1120 90 0 0 la_oenb[60]
port 504 nsew signal input
flabel metal2 s 344486 -800 344598 480 0 FreeSans 1120 90 0 0 la_oenb[61]
port 505 nsew signal input
flabel metal2 s 348032 -800 348144 480 0 FreeSans 1120 90 0 0 la_oenb[62]
port 506 nsew signal input
flabel metal2 s 351578 -800 351690 480 0 FreeSans 1120 90 0 0 la_oenb[63]
port 507 nsew signal input
flabel metal2 s 355124 -800 355236 480 0 FreeSans 1120 90 0 0 la_oenb[64]
port 508 nsew signal input
flabel metal2 s 358670 -800 358782 480 0 FreeSans 1120 90 0 0 la_oenb[65]
port 509 nsew signal input
flabel metal2 s 362216 -800 362328 480 0 FreeSans 1120 90 0 0 la_oenb[66]
port 510 nsew signal input
flabel metal2 s 365762 -800 365874 480 0 FreeSans 1120 90 0 0 la_oenb[67]
port 511 nsew signal input
flabel metal2 s 369308 -800 369420 480 0 FreeSans 1120 90 0 0 la_oenb[68]
port 512 nsew signal input
flabel metal2 s 372854 -800 372966 480 0 FreeSans 1120 90 0 0 la_oenb[69]
port 513 nsew signal input
flabel metal2 s 149456 -800 149568 480 0 FreeSans 1120 90 0 0 la_oenb[6]
port 514 nsew signal input
flabel metal2 s 376400 -800 376512 480 0 FreeSans 1120 90 0 0 la_oenb[70]
port 515 nsew signal input
flabel metal2 s 379946 -800 380058 480 0 FreeSans 1120 90 0 0 la_oenb[71]
port 516 nsew signal input
flabel metal2 s 383492 -800 383604 480 0 FreeSans 1120 90 0 0 la_oenb[72]
port 517 nsew signal input
flabel metal2 s 387038 -800 387150 480 0 FreeSans 1120 90 0 0 la_oenb[73]
port 518 nsew signal input
flabel metal2 s 390584 -800 390696 480 0 FreeSans 1120 90 0 0 la_oenb[74]
port 519 nsew signal input
flabel metal2 s 394130 -800 394242 480 0 FreeSans 1120 90 0 0 la_oenb[75]
port 520 nsew signal input
flabel metal2 s 397676 -800 397788 480 0 FreeSans 1120 90 0 0 la_oenb[76]
port 521 nsew signal input
flabel metal2 s 401222 -800 401334 480 0 FreeSans 1120 90 0 0 la_oenb[77]
port 522 nsew signal input
flabel metal2 s 404768 -800 404880 480 0 FreeSans 1120 90 0 0 la_oenb[78]
port 523 nsew signal input
flabel metal2 s 408314 -800 408426 480 0 FreeSans 1120 90 0 0 la_oenb[79]
port 524 nsew signal input
flabel metal2 s 153002 -800 153114 480 0 FreeSans 1120 90 0 0 la_oenb[7]
port 525 nsew signal input
flabel metal2 s 411860 -800 411972 480 0 FreeSans 1120 90 0 0 la_oenb[80]
port 526 nsew signal input
flabel metal2 s 415406 -800 415518 480 0 FreeSans 1120 90 0 0 la_oenb[81]
port 527 nsew signal input
flabel metal2 s 418952 -800 419064 480 0 FreeSans 1120 90 0 0 la_oenb[82]
port 528 nsew signal input
flabel metal2 s 422498 -800 422610 480 0 FreeSans 1120 90 0 0 la_oenb[83]
port 529 nsew signal input
flabel metal2 s 426044 -800 426156 480 0 FreeSans 1120 90 0 0 la_oenb[84]
port 530 nsew signal input
flabel metal2 s 429590 -800 429702 480 0 FreeSans 1120 90 0 0 la_oenb[85]
port 531 nsew signal input
flabel metal2 s 433136 -800 433248 480 0 FreeSans 1120 90 0 0 la_oenb[86]
port 532 nsew signal input
flabel metal2 s 436682 -800 436794 480 0 FreeSans 1120 90 0 0 la_oenb[87]
port 533 nsew signal input
flabel metal2 s 440228 -800 440340 480 0 FreeSans 1120 90 0 0 la_oenb[88]
port 534 nsew signal input
flabel metal2 s 443774 -800 443886 480 0 FreeSans 1120 90 0 0 la_oenb[89]
port 535 nsew signal input
flabel metal2 s 156548 -800 156660 480 0 FreeSans 1120 90 0 0 la_oenb[8]
port 536 nsew signal input
flabel metal2 s 447320 -800 447432 480 0 FreeSans 1120 90 0 0 la_oenb[90]
port 537 nsew signal input
flabel metal2 s 450866 -800 450978 480 0 FreeSans 1120 90 0 0 la_oenb[91]
port 538 nsew signal input
flabel metal2 s 454412 -800 454524 480 0 FreeSans 1120 90 0 0 la_oenb[92]
port 539 nsew signal input
flabel metal2 s 457958 -800 458070 480 0 FreeSans 1120 90 0 0 la_oenb[93]
port 540 nsew signal input
flabel metal2 s 461504 -800 461616 480 0 FreeSans 1120 90 0 0 la_oenb[94]
port 541 nsew signal input
flabel metal2 s 465050 -800 465162 480 0 FreeSans 1120 90 0 0 la_oenb[95]
port 542 nsew signal input
flabel metal2 s 468596 -800 468708 480 0 FreeSans 1120 90 0 0 la_oenb[96]
port 543 nsew signal input
flabel metal2 s 472142 -800 472254 480 0 FreeSans 1120 90 0 0 la_oenb[97]
port 544 nsew signal input
flabel metal2 s 475688 -800 475800 480 0 FreeSans 1120 90 0 0 la_oenb[98]
port 545 nsew signal input
flabel metal2 s 479234 -800 479346 480 0 FreeSans 1120 90 0 0 la_oenb[99]
port 546 nsew signal input
flabel metal2 s 160094 -800 160206 480 0 FreeSans 1120 90 0 0 la_oenb[9]
port 547 nsew signal input
flabel metal2 s 579704 -800 579816 480 0 FreeSans 1120 90 0 0 user_clock2
port 548 nsew signal input
flabel metal2 s 580886 -800 580998 480 0 FreeSans 1120 90 0 0 user_irq[0]
port 549 nsew signal tristate
flabel metal2 s 582068 -800 582180 480 0 FreeSans 1120 90 0 0 user_irq[1]
port 550 nsew signal tristate
flabel metal2 s 583250 -800 583362 480 0 FreeSans 1120 90 0 0 user_irq[2]
port 551 nsew signal tristate
flabel metal3 s 582340 639784 584800 644584 0 FreeSans 1120 0 0 0 vccd1
port 552 nsew signal bidirectional
flabel metal3 s 582340 629784 584800 634584 0 FreeSans 1120 0 0 0 vccd1
port 553 nsew signal bidirectional
flabel metal3 s 0 643842 1660 648642 0 FreeSans 1120 0 0 0 vccd2
port 554 nsew signal bidirectional
flabel metal3 s 0 633842 1660 638642 0 FreeSans 1120 0 0 0 vccd2
port 555 nsew signal bidirectional
flabel metal3 s 582340 540562 584800 545362 0 FreeSans 1120 0 0 0 vdda1
port 556 nsew signal bidirectional
flabel metal3 s 582340 550562 584800 555362 0 FreeSans 1120 0 0 0 vdda1
port 557 nsew signal bidirectional
flabel metal3 s 582340 235230 584800 240030 0 FreeSans 1120 0 0 0 vdda1
port 558 nsew signal bidirectional
flabel metal3 s 582340 225230 584800 230030 0 FreeSans 1120 0 0 0 vdda1
port 559 nsew signal bidirectional
flabel metal3 s 0 204888 1660 209688 0 FreeSans 1120 0 0 0 vdda2
port 560 nsew signal bidirectional
flabel metal3 s 0 214888 1660 219688 0 FreeSans 1120 0 0 0 vdda2
port 561 nsew signal bidirectional
flabel metal3 s 520594 702340 525394 704800 0 FreeSans 1920 180 0 0 vssa1
port 562 nsew signal bidirectional
flabel metal3 s 510594 702340 515394 704800 0 FreeSans 1920 180 0 0 vssa1
port 563 nsew signal bidirectional
flabel metal3 s 582340 146830 584800 151630 0 FreeSans 1120 0 0 0 vssa1
port 564 nsew signal bidirectional
flabel metal3 s 582340 136830 584800 141630 0 FreeSans 1120 0 0 0 vssa1
port 565 nsew signal bidirectional
flabel metal3 s 0 559442 1660 564242 0 FreeSans 1120 0 0 0 vssa2
port 566 nsew signal bidirectional
flabel metal3 s 0 549442 1660 554242 0 FreeSans 1120 0 0 0 vssa2
port 567 nsew signal bidirectional
flabel metal3 s 582340 191430 584800 196230 0 FreeSans 1120 0 0 0 vssd1
port 568 nsew signal bidirectional
flabel metal3 s 582340 181430 584800 186230 0 FreeSans 1120 0 0 0 vssd1
port 569 nsew signal bidirectional
flabel metal3 s 0 172888 1660 177688 0 FreeSans 1120 0 0 0 vssd2
port 570 nsew signal bidirectional
flabel metal3 s 0 162888 1660 167688 0 FreeSans 1120 0 0 0 vssd2
port 571 nsew signal bidirectional
flabel metal2 s 524 -800 636 480 0 FreeSans 1120 90 0 0 wb_clk_i
port 572 nsew signal input
flabel metal2 s 1706 -800 1818 480 0 FreeSans 1120 90 0 0 wb_rst_i
port 573 nsew signal input
flabel metal2 s 2888 -800 3000 480 0 FreeSans 1120 90 0 0 wbs_ack_o
port 574 nsew signal tristate
flabel metal2 s 7616 -800 7728 480 0 FreeSans 1120 90 0 0 wbs_adr_i[0]
port 575 nsew signal input
flabel metal2 s 47804 -800 47916 480 0 FreeSans 1120 90 0 0 wbs_adr_i[10]
port 576 nsew signal input
flabel metal2 s 51350 -800 51462 480 0 FreeSans 1120 90 0 0 wbs_adr_i[11]
port 577 nsew signal input
flabel metal2 s 54896 -800 55008 480 0 FreeSans 1120 90 0 0 wbs_adr_i[12]
port 578 nsew signal input
flabel metal2 s 58442 -800 58554 480 0 FreeSans 1120 90 0 0 wbs_adr_i[13]
port 579 nsew signal input
flabel metal2 s 61988 -800 62100 480 0 FreeSans 1120 90 0 0 wbs_adr_i[14]
port 580 nsew signal input
flabel metal2 s 65534 -800 65646 480 0 FreeSans 1120 90 0 0 wbs_adr_i[15]
port 581 nsew signal input
flabel metal2 s 69080 -800 69192 480 0 FreeSans 1120 90 0 0 wbs_adr_i[16]
port 582 nsew signal input
flabel metal2 s 72626 -800 72738 480 0 FreeSans 1120 90 0 0 wbs_adr_i[17]
port 583 nsew signal input
flabel metal2 s 76172 -800 76284 480 0 FreeSans 1120 90 0 0 wbs_adr_i[18]
port 584 nsew signal input
flabel metal2 s 79718 -800 79830 480 0 FreeSans 1120 90 0 0 wbs_adr_i[19]
port 585 nsew signal input
flabel metal2 s 12344 -800 12456 480 0 FreeSans 1120 90 0 0 wbs_adr_i[1]
port 586 nsew signal input
flabel metal2 s 83264 -800 83376 480 0 FreeSans 1120 90 0 0 wbs_adr_i[20]
port 587 nsew signal input
flabel metal2 s 86810 -800 86922 480 0 FreeSans 1120 90 0 0 wbs_adr_i[21]
port 588 nsew signal input
flabel metal2 s 90356 -800 90468 480 0 FreeSans 1120 90 0 0 wbs_adr_i[22]
port 589 nsew signal input
flabel metal2 s 93902 -800 94014 480 0 FreeSans 1120 90 0 0 wbs_adr_i[23]
port 590 nsew signal input
flabel metal2 s 97448 -800 97560 480 0 FreeSans 1120 90 0 0 wbs_adr_i[24]
port 591 nsew signal input
flabel metal2 s 100994 -800 101106 480 0 FreeSans 1120 90 0 0 wbs_adr_i[25]
port 592 nsew signal input
flabel metal2 s 104540 -800 104652 480 0 FreeSans 1120 90 0 0 wbs_adr_i[26]
port 593 nsew signal input
flabel metal2 s 108086 -800 108198 480 0 FreeSans 1120 90 0 0 wbs_adr_i[27]
port 594 nsew signal input
flabel metal2 s 111632 -800 111744 480 0 FreeSans 1120 90 0 0 wbs_adr_i[28]
port 595 nsew signal input
flabel metal2 s 115178 -800 115290 480 0 FreeSans 1120 90 0 0 wbs_adr_i[29]
port 596 nsew signal input
flabel metal2 s 17072 -800 17184 480 0 FreeSans 1120 90 0 0 wbs_adr_i[2]
port 597 nsew signal input
flabel metal2 s 118724 -800 118836 480 0 FreeSans 1120 90 0 0 wbs_adr_i[30]
port 598 nsew signal input
flabel metal2 s 122270 -800 122382 480 0 FreeSans 1120 90 0 0 wbs_adr_i[31]
port 599 nsew signal input
flabel metal2 s 21800 -800 21912 480 0 FreeSans 1120 90 0 0 wbs_adr_i[3]
port 600 nsew signal input
flabel metal2 s 26528 -800 26640 480 0 FreeSans 1120 90 0 0 wbs_adr_i[4]
port 601 nsew signal input
flabel metal2 s 30074 -800 30186 480 0 FreeSans 1120 90 0 0 wbs_adr_i[5]
port 602 nsew signal input
flabel metal2 s 33620 -800 33732 480 0 FreeSans 1120 90 0 0 wbs_adr_i[6]
port 603 nsew signal input
flabel metal2 s 37166 -800 37278 480 0 FreeSans 1120 90 0 0 wbs_adr_i[7]
port 604 nsew signal input
flabel metal2 s 40712 -800 40824 480 0 FreeSans 1120 90 0 0 wbs_adr_i[8]
port 605 nsew signal input
flabel metal2 s 44258 -800 44370 480 0 FreeSans 1120 90 0 0 wbs_adr_i[9]
port 606 nsew signal input
flabel metal2 s 4070 -800 4182 480 0 FreeSans 1120 90 0 0 wbs_cyc_i
port 607 nsew signal input
flabel metal2 s 8798 -800 8910 480 0 FreeSans 1120 90 0 0 wbs_dat_i[0]
port 608 nsew signal input
flabel metal2 s 48986 -800 49098 480 0 FreeSans 1120 90 0 0 wbs_dat_i[10]
port 609 nsew signal input
flabel metal2 s 52532 -800 52644 480 0 FreeSans 1120 90 0 0 wbs_dat_i[11]
port 610 nsew signal input
flabel metal2 s 56078 -800 56190 480 0 FreeSans 1120 90 0 0 wbs_dat_i[12]
port 611 nsew signal input
flabel metal2 s 59624 -800 59736 480 0 FreeSans 1120 90 0 0 wbs_dat_i[13]
port 612 nsew signal input
flabel metal2 s 63170 -800 63282 480 0 FreeSans 1120 90 0 0 wbs_dat_i[14]
port 613 nsew signal input
flabel metal2 s 66716 -800 66828 480 0 FreeSans 1120 90 0 0 wbs_dat_i[15]
port 614 nsew signal input
flabel metal2 s 70262 -800 70374 480 0 FreeSans 1120 90 0 0 wbs_dat_i[16]
port 615 nsew signal input
flabel metal2 s 73808 -800 73920 480 0 FreeSans 1120 90 0 0 wbs_dat_i[17]
port 616 nsew signal input
flabel metal2 s 77354 -800 77466 480 0 FreeSans 1120 90 0 0 wbs_dat_i[18]
port 617 nsew signal input
flabel metal2 s 80900 -800 81012 480 0 FreeSans 1120 90 0 0 wbs_dat_i[19]
port 618 nsew signal input
flabel metal2 s 13526 -800 13638 480 0 FreeSans 1120 90 0 0 wbs_dat_i[1]
port 619 nsew signal input
flabel metal2 s 84446 -800 84558 480 0 FreeSans 1120 90 0 0 wbs_dat_i[20]
port 620 nsew signal input
flabel metal2 s 87992 -800 88104 480 0 FreeSans 1120 90 0 0 wbs_dat_i[21]
port 621 nsew signal input
flabel metal2 s 91538 -800 91650 480 0 FreeSans 1120 90 0 0 wbs_dat_i[22]
port 622 nsew signal input
flabel metal2 s 95084 -800 95196 480 0 FreeSans 1120 90 0 0 wbs_dat_i[23]
port 623 nsew signal input
flabel metal2 s 98630 -800 98742 480 0 FreeSans 1120 90 0 0 wbs_dat_i[24]
port 624 nsew signal input
flabel metal2 s 102176 -800 102288 480 0 FreeSans 1120 90 0 0 wbs_dat_i[25]
port 625 nsew signal input
flabel metal2 s 105722 -800 105834 480 0 FreeSans 1120 90 0 0 wbs_dat_i[26]
port 626 nsew signal input
flabel metal2 s 109268 -800 109380 480 0 FreeSans 1120 90 0 0 wbs_dat_i[27]
port 627 nsew signal input
flabel metal2 s 112814 -800 112926 480 0 FreeSans 1120 90 0 0 wbs_dat_i[28]
port 628 nsew signal input
flabel metal2 s 116360 -800 116472 480 0 FreeSans 1120 90 0 0 wbs_dat_i[29]
port 629 nsew signal input
flabel metal2 s 18254 -800 18366 480 0 FreeSans 1120 90 0 0 wbs_dat_i[2]
port 630 nsew signal input
flabel metal2 s 119906 -800 120018 480 0 FreeSans 1120 90 0 0 wbs_dat_i[30]
port 631 nsew signal input
flabel metal2 s 123452 -800 123564 480 0 FreeSans 1120 90 0 0 wbs_dat_i[31]
port 632 nsew signal input
flabel metal2 s 22982 -800 23094 480 0 FreeSans 1120 90 0 0 wbs_dat_i[3]
port 633 nsew signal input
flabel metal2 s 27710 -800 27822 480 0 FreeSans 1120 90 0 0 wbs_dat_i[4]
port 634 nsew signal input
flabel metal2 s 31256 -800 31368 480 0 FreeSans 1120 90 0 0 wbs_dat_i[5]
port 635 nsew signal input
flabel metal2 s 34802 -800 34914 480 0 FreeSans 1120 90 0 0 wbs_dat_i[6]
port 636 nsew signal input
flabel metal2 s 38348 -800 38460 480 0 FreeSans 1120 90 0 0 wbs_dat_i[7]
port 637 nsew signal input
flabel metal2 s 41894 -800 42006 480 0 FreeSans 1120 90 0 0 wbs_dat_i[8]
port 638 nsew signal input
flabel metal2 s 45440 -800 45552 480 0 FreeSans 1120 90 0 0 wbs_dat_i[9]
port 639 nsew signal input
flabel metal2 s 9980 -800 10092 480 0 FreeSans 1120 90 0 0 wbs_dat_o[0]
port 640 nsew signal tristate
flabel metal2 s 50168 -800 50280 480 0 FreeSans 1120 90 0 0 wbs_dat_o[10]
port 641 nsew signal tristate
flabel metal2 s 53714 -800 53826 480 0 FreeSans 1120 90 0 0 wbs_dat_o[11]
port 642 nsew signal tristate
flabel metal2 s 57260 -800 57372 480 0 FreeSans 1120 90 0 0 wbs_dat_o[12]
port 643 nsew signal tristate
flabel metal2 s 60806 -800 60918 480 0 FreeSans 1120 90 0 0 wbs_dat_o[13]
port 644 nsew signal tristate
flabel metal2 s 64352 -800 64464 480 0 FreeSans 1120 90 0 0 wbs_dat_o[14]
port 645 nsew signal tristate
flabel metal2 s 67898 -800 68010 480 0 FreeSans 1120 90 0 0 wbs_dat_o[15]
port 646 nsew signal tristate
flabel metal2 s 71444 -800 71556 480 0 FreeSans 1120 90 0 0 wbs_dat_o[16]
port 647 nsew signal tristate
flabel metal2 s 74990 -800 75102 480 0 FreeSans 1120 90 0 0 wbs_dat_o[17]
port 648 nsew signal tristate
flabel metal2 s 78536 -800 78648 480 0 FreeSans 1120 90 0 0 wbs_dat_o[18]
port 649 nsew signal tristate
flabel metal2 s 82082 -800 82194 480 0 FreeSans 1120 90 0 0 wbs_dat_o[19]
port 650 nsew signal tristate
flabel metal2 s 14708 -800 14820 480 0 FreeSans 1120 90 0 0 wbs_dat_o[1]
port 651 nsew signal tristate
flabel metal2 s 85628 -800 85740 480 0 FreeSans 1120 90 0 0 wbs_dat_o[20]
port 652 nsew signal tristate
flabel metal2 s 89174 -800 89286 480 0 FreeSans 1120 90 0 0 wbs_dat_o[21]
port 653 nsew signal tristate
flabel metal2 s 92720 -800 92832 480 0 FreeSans 1120 90 0 0 wbs_dat_o[22]
port 654 nsew signal tristate
flabel metal2 s 96266 -800 96378 480 0 FreeSans 1120 90 0 0 wbs_dat_o[23]
port 655 nsew signal tristate
flabel metal2 s 99812 -800 99924 480 0 FreeSans 1120 90 0 0 wbs_dat_o[24]
port 656 nsew signal tristate
flabel metal2 s 103358 -800 103470 480 0 FreeSans 1120 90 0 0 wbs_dat_o[25]
port 657 nsew signal tristate
flabel metal2 s 106904 -800 107016 480 0 FreeSans 1120 90 0 0 wbs_dat_o[26]
port 658 nsew signal tristate
flabel metal2 s 110450 -800 110562 480 0 FreeSans 1120 90 0 0 wbs_dat_o[27]
port 659 nsew signal tristate
flabel metal2 s 113996 -800 114108 480 0 FreeSans 1120 90 0 0 wbs_dat_o[28]
port 660 nsew signal tristate
flabel metal2 s 117542 -800 117654 480 0 FreeSans 1120 90 0 0 wbs_dat_o[29]
port 661 nsew signal tristate
flabel metal2 s 19436 -800 19548 480 0 FreeSans 1120 90 0 0 wbs_dat_o[2]
port 662 nsew signal tristate
flabel metal2 s 121088 -800 121200 480 0 FreeSans 1120 90 0 0 wbs_dat_o[30]
port 663 nsew signal tristate
flabel metal2 s 124634 -800 124746 480 0 FreeSans 1120 90 0 0 wbs_dat_o[31]
port 664 nsew signal tristate
flabel metal2 s 24164 -800 24276 480 0 FreeSans 1120 90 0 0 wbs_dat_o[3]
port 665 nsew signal tristate
flabel metal2 s 28892 -800 29004 480 0 FreeSans 1120 90 0 0 wbs_dat_o[4]
port 666 nsew signal tristate
flabel metal2 s 32438 -800 32550 480 0 FreeSans 1120 90 0 0 wbs_dat_o[5]
port 667 nsew signal tristate
flabel metal2 s 35984 -800 36096 480 0 FreeSans 1120 90 0 0 wbs_dat_o[6]
port 668 nsew signal tristate
flabel metal2 s 39530 -800 39642 480 0 FreeSans 1120 90 0 0 wbs_dat_o[7]
port 669 nsew signal tristate
flabel metal2 s 43076 -800 43188 480 0 FreeSans 1120 90 0 0 wbs_dat_o[8]
port 670 nsew signal tristate
flabel metal2 s 46622 -800 46734 480 0 FreeSans 1120 90 0 0 wbs_dat_o[9]
port 671 nsew signal tristate
flabel metal2 s 11162 -800 11274 480 0 FreeSans 1120 90 0 0 wbs_sel_i[0]
port 672 nsew signal input
flabel metal2 s 15890 -800 16002 480 0 FreeSans 1120 90 0 0 wbs_sel_i[1]
port 673 nsew signal input
flabel metal2 s 20618 -800 20730 480 0 FreeSans 1120 90 0 0 wbs_sel_i[2]
port 674 nsew signal input
flabel metal2 s 25346 -800 25458 480 0 FreeSans 1120 90 0 0 wbs_sel_i[3]
port 675 nsew signal input
flabel metal2 s 5252 -800 5364 480 0 FreeSans 1120 90 0 0 wbs_stb_i
port 676 nsew signal input
flabel metal2 s 6434 -800 6546 480 0 FreeSans 1120 90 0 0 wbs_we_i
port 677 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
