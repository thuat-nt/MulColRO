** sch_path: /run/media/thuat/build/cmos/MulColRO/xschem/user_analog_project_wrapper.sch
.subckt user_analog_project_wrapper vdda1 vdda2 vssa1 vssa2 vccd1 vccd2 vssd1 vssd2 wb_clk_i
+ wb_rst_i wbs_stb_i wbs_cyc_i wbs_we_i wbs_sel_i[3] wbs_sel_i[2] wbs_sel_i[1] wbs_sel_i[0] wbs_dat_i[31]
+ wbs_dat_i[30] wbs_dat_i[29] wbs_dat_i[28] wbs_dat_i[27] wbs_dat_i[26] wbs_dat_i[25] wbs_dat_i[24] wbs_dat_i[23]
+ wbs_dat_i[22] wbs_dat_i[21] wbs_dat_i[20] wbs_dat_i[19] wbs_dat_i[18] wbs_dat_i[17] wbs_dat_i[16] wbs_dat_i[15]
+ wbs_dat_i[14] wbs_dat_i[13] wbs_dat_i[12] wbs_dat_i[11] wbs_dat_i[10] wbs_dat_i[9] wbs_dat_i[8] wbs_dat_i[7]
+ wbs_dat_i[6] wbs_dat_i[5] wbs_dat_i[4] wbs_dat_i[3] wbs_dat_i[2] wbs_dat_i[1] wbs_dat_i[0] wbs_adr_i[31]
+ wbs_adr_i[30] wbs_adr_i[29] wbs_adr_i[28] wbs_adr_i[27] wbs_adr_i[26] wbs_adr_i[25] wbs_adr_i[24] wbs_adr_i[23]
+ wbs_adr_i[22] wbs_adr_i[21] wbs_adr_i[20] wbs_adr_i[19] wbs_adr_i[18] wbs_adr_i[17] wbs_adr_i[16] wbs_adr_i[15]
+ wbs_adr_i[14] wbs_adr_i[13] wbs_adr_i[12] wbs_adr_i[11] wbs_adr_i[10] wbs_adr_i[9] wbs_adr_i[8] wbs_adr_i[7]
+ wbs_adr_i[6] wbs_adr_i[5] wbs_adr_i[4] wbs_adr_i[3] wbs_adr_i[2] wbs_adr_i[1] wbs_adr_i[0] wbs_ack_o
+ wbs_dat_o[31] wbs_dat_o[30] wbs_dat_o[29] wbs_dat_o[28] wbs_dat_o[27] wbs_dat_o[26] wbs_dat_o[25] wbs_dat_o[24]
+ wbs_dat_o[23] wbs_dat_o[22] wbs_dat_o[21] wbs_dat_o[20] wbs_dat_o[19] wbs_dat_o[18] wbs_dat_o[17] wbs_dat_o[16]
+ wbs_dat_o[15] wbs_dat_o[14] wbs_dat_o[13] wbs_dat_o[12] wbs_dat_o[11] wbs_dat_o[10] wbs_dat_o[9] wbs_dat_o[8]
+ wbs_dat_o[7] wbs_dat_o[6] wbs_dat_o[5] wbs_dat_o[4] wbs_dat_o[3] wbs_dat_o[2] wbs_dat_o[1] wbs_dat_o[0]
+ la_data_in[127] la_data_in[126] la_data_in[125] la_data_in[124] la_data_in[123] la_data_in[122] la_data_in[121]
+ la_data_in[120] la_data_in[119] la_data_in[118] la_data_in[117] la_data_in[116] la_data_in[115] la_data_in[114]
+ la_data_in[113] la_data_in[112] la_data_in[111] la_data_in[110] la_data_in[109] la_data_in[108] la_data_in[107]
+ la_data_in[106] la_data_in[105] la_data_in[104] la_data_in[103] la_data_in[102] la_data_in[101] la_data_in[100]
+ la_data_in[99] la_data_in[98] la_data_in[97] la_data_in[96] la_data_in[95] la_data_in[94] la_data_in[93]
+ la_data_in[92] la_data_in[91] la_data_in[90] la_data_in[89] la_data_in[88] la_data_in[87] la_data_in[86]
+ la_data_in[85] la_data_in[84] la_data_in[83] la_data_in[82] la_data_in[81] la_data_in[80] la_data_in[79]
+ la_data_in[78] la_data_in[77] la_data_in[76] la_data_in[75] la_data_in[74] la_data_in[73] la_data_in[72]
+ la_data_in[71] la_data_in[70] la_data_in[69] la_data_in[68] la_data_in[67] la_data_in[66] la_data_in[65]
+ la_data_in[64] la_data_in[63] la_data_in[62] la_data_in[61] la_data_in[60] la_data_in[59] la_data_in[58]
+ la_data_in[57] la_data_in[56] la_data_in[55] la_data_in[54] la_data_in[53] la_data_in[52] la_data_in[51]
+ la_data_in[50] la_data_in[49] la_data_in[48] la_data_in[47] la_data_in[46] la_data_in[45] la_data_in[44]
+ la_data_in[43] la_data_in[42] la_data_in[41] la_data_in[40] la_data_in[39] la_data_in[38] la_data_in[37]
+ la_data_in[36] la_data_in[35] la_data_in[34] la_data_in[33] la_data_in[32] la_data_in[31] la_data_in[30]
+ la_data_in[29] la_data_in[28] la_data_in[27] la_data_in[26] la_data_in[25] la_data_in[24] la_data_in[23]
+ la_data_in[22] la_data_in[21] la_data_in[20] la_data_in[19] la_data_in[18] la_data_in[17] la_data_in[16]
+ la_data_in[15] la_data_in[14] la_data_in[13] la_data_in[12] la_data_in[11] la_data_in[10] la_data_in[9]
+ la_data_in[8] la_data_in[7] la_data_in[6] la_data_in[5] la_data_in[4] la_data_in[3] la_data_in[2] la_data_in[1]
+ la_data_in[0] la_data_out[127] la_data_out[126] la_data_out[125] la_data_out[124] la_data_out[123]
+ la_data_out[122] la_data_out[121] la_data_out[120] la_data_out[119] la_data_out[118] la_data_out[117]
+ la_data_out[116] la_data_out[115] la_data_out[114] la_data_out[113] la_data_out[112] la_data_out[111]
+ la_data_out[110] la_data_out[109] la_data_out[108] la_data_out[107] la_data_out[106] la_data_out[105]
+ la_data_out[104] la_data_out[103] la_data_out[102] la_data_out[101] la_data_out[100] la_data_out[99] la_data_out[98]
+ la_data_out[97] la_data_out[96] la_data_out[95] la_data_out[94] la_data_out[93] la_data_out[92] la_data_out[91]
+ la_data_out[90] la_data_out[89] la_data_out[88] la_data_out[87] la_data_out[86] la_data_out[85] la_data_out[84]
+ la_data_out[83] la_data_out[82] la_data_out[81] la_data_out[80] la_data_out[79] la_data_out[78] la_data_out[77]
+ la_data_out[76] la_data_out[75] la_data_out[74] la_data_out[73] la_data_out[72] la_data_out[71] la_data_out[70]
+ la_data_out[69] la_data_out[68] la_data_out[67] la_data_out[66] la_data_out[65] la_data_out[64] la_data_out[63]
+ la_data_out[62] la_data_out[61] la_data_out[60] la_data_out[59] la_data_out[58] la_data_out[57] la_data_out[56]
+ la_data_out[55] la_data_out[54] la_data_out[53] la_data_out[52] la_data_out[51] la_data_out[50] la_data_out[49]
+ la_data_out[48] la_data_out[47] la_data_out[46] la_data_out[45] la_data_out[44] la_data_out[43] la_data_out[42]
+ la_data_out[41] la_data_out[40] la_data_out[39] la_data_out[38] la_data_out[37] la_data_out[36] la_data_out[35]
+ la_data_out[34] la_data_out[33] la_data_out[32] la_data_out[31] la_data_out[30] la_data_out[29] la_data_out[28]
+ la_data_out[27] la_data_out[26] la_data_out[25] la_data_out[24] la_data_out[23] la_data_out[22] la_data_out[21]
+ la_data_out[20] la_data_out[19] la_data_out[18] la_data_out[17] la_data_out[16] la_data_out[15] la_data_out[14]
+ la_data_out[13] la_data_out[12] la_data_out[11] la_data_out[10] la_data_out[9] la_data_out[8] la_data_out[7]
+ la_data_out[6] la_data_out[5] la_data_out[4] la_data_out[3] la_data_out[2] la_data_out[1] la_data_out[0] io_in[26]
+ io_in[25] io_in[24] io_in[23] io_in[22] io_in[21] io_in[20] io_in[19] io_in[18] io_in[17] io_in[16] io_in[15]
+ io_in[14] io_in[13] io_in[12] io_in[11] io_in[10] io_in[9] io_in[8] io_in[7] io_in[6] io_in[5] io_in[4]
+ io_in[3] io_in[2] io_in[1] io_in[0] io_in_3v3[26] io_in_3v3[25] io_in_3v3[24] io_in_3v3[23] io_in_3v3[22]
+ io_in_3v3[21] io_in_3v3[20] io_in_3v3[19] io_in_3v3[18] io_in_3v3[17] io_in_3v3[16] io_in_3v3[15] io_in_3v3[14]
+ io_in_3v3[13] io_in_3v3[12] io_in_3v3[11] io_in_3v3[10] io_in_3v3[9] io_in_3v3[8] io_in_3v3[7] io_in_3v3[6]
+ io_in_3v3[5] io_in_3v3[4] io_in_3v3[3] io_in_3v3[2] io_in_3v3[1] io_in_3v3[0] user_clock2 io_out[26] io_out[25]
+ io_out[24] io_out[23] io_out[22] io_out[21] io_out[20] io_out[19] io_out[18] io_out[17] io_out[16] io_out[15]
+ io_out[14] io_out[13] io_out[12] io_out[11] io_out[10] io_out[9] io_out[8] io_out[7] io_out[6] io_out[5]
+ io_out[4] io_out[3] io_out[2] io_out[1] io_out[0] io_oeb[26] io_oeb[25] io_oeb[24] io_oeb[23] io_oeb[22]
+ io_oeb[21] io_oeb[20] io_oeb[19] io_oeb[18] io_oeb[17] io_oeb[16] io_oeb[15] io_oeb[14] io_oeb[13] io_oeb[12]
+ io_oeb[11] io_oeb[10] io_oeb[9] io_oeb[8] io_oeb[7] io_oeb[6] io_oeb[5] io_oeb[4] io_oeb[3] io_oeb[2]
+ io_oeb[1] io_oeb[0] gpio_analog[17] gpio_analog[16] gpio_analog[15] gpio_analog[14] gpio_analog[13]
+ gpio_analog[12] gpio_analog[11] gpio_analog[10] gpio_analog[9] gpio_analog[8] gpio_analog[7] gpio_analog[6]
+ gpio_analog[5] gpio_analog[4] gpio_analog[3] gpio_analog[2] gpio_analog[1] gpio_analog[0] gpio_noesd[17]
+ gpio_noesd[16] gpio_noesd[15] gpio_noesd[14] gpio_noesd[13] gpio_noesd[12] gpio_noesd[11] gpio_noesd[10]
+ gpio_noesd[9] gpio_noesd[8] gpio_noesd[7] gpio_noesd[6] gpio_noesd[5] gpio_noesd[4] gpio_noesd[3] gpio_noesd[2]
+ gpio_noesd[1] gpio_noesd[0] io_analog[10] io_analog[9] io_analog[8] io_analog[7] io_analog[6] io_analog[5]
+ io_analog[4] io_analog[3] io_analog[2] io_analog[1] io_analog[0] io_clamp_high[2] io_clamp_high[1]
+ io_clamp_high[0] io_clamp_low[2] io_clamp_low[1] io_clamp_low[0] user_irq[2] user_irq[1] user_irq[0] la_oenb[127]
+ la_oenb[126] la_oenb[125] la_oenb[124] la_oenb[123] la_oenb[122] la_oenb[121] la_oenb[120] la_oenb[119]
+ la_oenb[118] la_oenb[117] la_oenb[116] la_oenb[115] la_oenb[114] la_oenb[113] la_oenb[112] la_oenb[111]
+ la_oenb[110] la_oenb[109] la_oenb[108] la_oenb[107] la_oenb[106] la_oenb[105] la_oenb[104] la_oenb[103]
+ la_oenb[102] la_oenb[101] la_oenb[100] la_oenb[99] la_oenb[98] la_oenb[97] la_oenb[96] la_oenb[95] la_oenb[94]
+ la_oenb[93] la_oenb[92] la_oenb[91] la_oenb[90] la_oenb[89] la_oenb[88] la_oenb[87] la_oenb[86] la_oenb[85]
+ la_oenb[84] la_oenb[83] la_oenb[82] la_oenb[81] la_oenb[80] la_oenb[79] la_oenb[78] la_oenb[77] la_oenb[76]
+ la_oenb[75] la_oenb[74] la_oenb[73] la_oenb[72] la_oenb[71] la_oenb[70] la_oenb[69] la_oenb[68] la_oenb[67]
+ la_oenb[66] la_oenb[65] la_oenb[64] la_oenb[63] la_oenb[62] la_oenb[61] la_oenb[60] la_oenb[59] la_oenb[58]
+ la_oenb[57] la_oenb[56] la_oenb[55] la_oenb[54] la_oenb[53] la_oenb[52] la_oenb[51] la_oenb[50] la_oenb[49]
+ la_oenb[48] la_oenb[47] la_oenb[46] la_oenb[45] la_oenb[44] la_oenb[43] la_oenb[42] la_oenb[41] la_oenb[40]
+ la_oenb[39] la_oenb[38] la_oenb[37] la_oenb[36] la_oenb[35] la_oenb[34] la_oenb[33] la_oenb[32] la_oenb[31]
+ la_oenb[30] la_oenb[29] la_oenb[28] la_oenb[27] la_oenb[26] la_oenb[25] la_oenb[24] la_oenb[23] la_oenb[22]
+ la_oenb[21] la_oenb[20] la_oenb[19] la_oenb[18] la_oenb[17] la_oenb[16] la_oenb[15] la_oenb[14] la_oenb[13]
+ la_oenb[12] la_oenb[11] la_oenb[10] la_oenb[9] la_oenb[8] la_oenb[7] la_oenb[6] la_oenb[5] la_oenb[4]
+ la_oenb[3] la_oenb[2] la_oenb[1] la_oenb[0] vdda1
*.PININFO vdda1:B vdda2:B vssa1:B vssa2:B vccd1:B vccd2:B vssd1:B vssd2:B wb_clk_i:I wb_rst_i:I
*+ wbs_stb_i:I wbs_cyc_i:I wbs_we_i:I wbs_sel_i[3:0]:I wbs_dat_i[31:0]:I wbs_adr_i[31:0]:I wbs_ack_o:O
*+ wbs_dat_o[31:0]:O la_data_in[127:0]:I la_data_out[127:0]:O io_in[26:0]:I io_in_3v3[26:0]:I user_clock2:I
*+ io_out[26:0]:O io_oeb[26:0]:O gpio_analog[17:0]:B gpio_noesd[17:0]:B io_analog[10:0]:B io_clamp_high[2:0]:B
*+ io_clamp_low[2:0]:B user_irq[2:0]:O la_oenb[127:0]:I vdda1:B
R1 vssd1 io_clamp_low[2] sky130_fd_pr__res_generic_m3 W=11 L=0.25 m=1
R2 vssd1 io_clamp_high[2] sky130_fd_pr__res_generic_m3 W=11 L=0.25 m=1
R4 vssd1 io_clamp_low[1] sky130_fd_pr__res_generic_m3 W=11 L=0.25 m=1
R5 vssd1 io_clamp_high[1] sky130_fd_pr__res_generic_m3 W=11 L=0.25 m=1
R6 vssd1 io_clamp_low[0] sky130_fd_pr__res_generic_m3 W=11 L=0.25 m=1
R7 vssd1 io_clamp_high[0] sky130_fd_pr__res_generic_m3 W=11 L=0.25 m=1
x3 vccd1 vssd1 gpio_analog[6] io_analog[0] gpio_analog[5] gpio_analog[4] gpio_analog[3]
+ gpio_analog[2] gpio_analog[1] io_in[7] io_in[6] io_in[5] io_in[4] io_in[3] io_in[2] io_in[1] ColROs
XR[12] io_oeb[13] vccd1 R_0_125
XR[11] io_oeb[12] vccd1 R_0_125
XR[10] io_oeb[11] vccd1 R_0_125
XR[9] io_oeb[10] vccd1 R_0_125
XR[8] io_oeb[9] vccd1 R_0_125
XR[7] io_oeb[8] vccd1 R_0_125
XR[6] io_oeb[7] vccd1 R_0_125
XR[5] io_oeb[6] vccd1 R_0_125
XR[4] io_oeb[5] vccd1 R_0_125
XR[3] io_oeb[4] vccd1 R_0_125
XR[2] io_oeb[3] vccd1 R_0_125
XR[1] io_oeb[2] vccd1 R_0_125
XR[0] io_oeb[1] vccd1 R_0_125
.ends

* expanding   symbol:  ColROs.sym # of pins=16
** sym_path: /run/media/thuat/build/cmos/MulColRO/xschem/ColROs.sym
** sch_path: /run/media/thuat/build/cmos/MulColRO/xschem/ColROs.sch
.subckt ColROs VDD GROUND AIn0 AOut AIn1 AIn2 AIn3 AIn4 AIn5 REG0 REG1 REG2 REG3 REG4 REG5 REG6
*.PININFO AOut:O REG1:I REG2:I REG3:I REG0:I REG5:I REG6:I REG4:I AIn0:I AIn1:I AIn2:I AIn3:I AIn4:I
*+ AIn5:I GROUND:I VDD:I
x1 AIn3 net1 AIn0 AIn1 AIn2 diffamp
x2 REG3 REG2 net1 net2 AIn4 REG0 AIn5 REG1 REG5 REG4 integrator
x7 AIn4 net3 AOut buffer
x3 REG6 net2 net3 net1 mux2_1
.ends


* expanding   symbol:  R_0_125/R_0_125.sym # of pins=2
** sym_path: /run/media/thuat/build/cmos/MulColRO/xschem/R_0_125/R_0_125.sym
** sch_path: /run/media/thuat/build/cmos/MulColRO/xschem/R_0_125/R_0_125.sch
.subckt R_0_125 out in
*.PININFO in:I out:O
R1 in out sky130_fd_pr__res_generic_m1 W=10 L=10 m=1
.ends


* expanding   symbol:  diffamp/diffamp.sym # of pins=5
** sym_path: /run/media/thuat/build/cmos/MulColRO/xschem/diffamp/diffamp.sym
** sch_path: /run/media/thuat/build/cmos/MulColRO/xschem/diffamp/diffamp.sch
.subckt diffamp PCAS OUT REF PIX GM_BIAS
*.PININFO PCAS:I PIX:I REF:I GM_BIAS:I OUT:O
XM17 net4 GM_BIAS GND sky130_fd_pr__nfet_01v8_lvt L=15 W=20 nf=2 m=1
XM8 net2 net1 VDD sky130_fd_pr__pfet_01v8_lvt L=15 W=90 nf=3 m=1
XM1 net3 net1 VDD sky130_fd_pr__pfet_01v8_lvt L=15 W=90 nf=3 m=1
XM2 OUT PCAS net2 sky130_fd_pr__pfet_01v8_lvt L=3 W=90 nf=3 m=1
XM4 net1 PCAS net3 sky130_fd_pr__pfet_01v8_lvt L=3 W=90 nf=3 m=1
XM5 OUT PIX net4 sky130_fd_pr__nfet_01v8_lvt L=3.5 W=800 nf=35 m=1
XM6 net1 REF net4 sky130_fd_pr__nfet_01v8_lvt L=3.5 W=800 nf=35 m=1
.ends


* expanding   symbol:  Integrator/integrator.sym # of pins=10
** sym_path: /run/media/thuat/build/cmos/MulColRO/xschem/Integrator/integrator.sym
** sch_path: /run/media/thuat/build/cmos/MulColRO/xschem/Integrator/integrator.sch
.subckt integrator sw2 sw1 intin intout opbias en Vtune rst sw4 sw3
*.PININFO intin:I Vtune:I intout:O opbias:I sw1:I sw2:I rst:I en:I sw3:I sw4:I
XC1 net4 intout sky130_fd_pr__cap_mim_m3_1 W=50 L=50 m=1
XC2 net3 intout sky130_fd_pr__cap_mim_m3_1 W=50 L=50 m=1
x9 sw2 net3 net2 switch
x1 sw1 net4 net2 switch
x3 Vtune intin curr_mir
x4 opbias net1 net2 intout opamp
x5 rst intout net2 switch
x6 en net1 GND switch
x7 net5 en not
x2 net5 net2 intin switch
XC3 net6 intout sky130_fd_pr__cap_mim_m3_1 W=50 L=50 m=1
x10 sw3 net6 net2 switch
XC4 net7 intout sky130_fd_pr__cap_mim_m3_1 W=50 L=50 m=1
x8 sw4 net7 net2 switch
.ends


* expanding   symbol:  buffer/buffer.sym # of pins=3
** sym_path: /run/media/thuat/build/cmos/MulColRO/xschem/buffer/buffer.sym
** sch_path: /run/media/thuat/build/cmos/MulColRO/xschem/buffer/buffer.sch
.subckt buffer opbias in out
*.PININFO in:I opbias:I out:O
x1 opbias in out out opamp
.ends


* expanding   symbol:  mux2_1/mux2_1.sym # of pins=4
** sym_path: /run/media/thuat/build/cmos/MulColRO/xschem/mux2_1/mux2_1.sym
** sch_path: /run/media/thuat/build/cmos/MulColRO/xschem/mux2_1/mux2_1.sch
.subckt mux2_1 SEL0 IN1 OUT IN0
*.PININFO SEL0:I OUT:O IN1:I IN0:I
x1 net1 SEL0 not
x6 SEL0 OUT IN1 switch
x5 net1 OUT IN0 switch
.ends


* expanding   symbol:  switch/switch.sym # of pins=3
** sym_path: /run/media/thuat/build/cmos/MulColRO/xschem/switch/switch.sym
** sch_path: /run/media/thuat/build/cmos/MulColRO/xschem/switch/switch.sch
.subckt switch toggle out in
*.PININFO toggle:I in:I out:O
x1 net1 toggle not
XM26 out net1 in sky130_fd_pr__pfet_01v8_lvt L=3 W=200 nf=5 m=1
XM17 in toggle out sky130_fd_pr__nfet_01v8_lvt L=3 W=200 nf=5 m=1
.ends


* expanding   symbol:  current_mirror/curr_mir.sym # of pins=2
** sym_path: /run/media/thuat/build/cmos/MulColRO/xschem/current_mirror/curr_mir.sym
** sch_path: /run/media/thuat/build/cmos/MulColRO/xschem/current_mirror/curr_mir.sch
.subckt curr_mir Vtune Ib
*.PININFO Vtune:I Ib:B
XM1 net1 net1 GND GND sky130_fd_pr__nfet_01v8_lvt L=2 W=50 nf=1 m=1
XM2 Ib net1 GND GND sky130_fd_pr__nfet_01v8_lvt L=25 W=4 nf=1 m=1
XM10 net1 Vtune VDD VDD sky130_fd_pr__pfet_01v8_lvt L=10 W=10 nf=1 m=1
.ends


* expanding   symbol:  opamp/opamp.sym # of pins=4
** sym_path: /run/media/thuat/build/cmos/MulColRO/xschem/opamp/opamp.sym
** sch_path: /run/media/thuat/build/cmos/MulColRO/xschem/opamp/opamp.sch
.subckt opamp opbias inp inn out
*.PININFO inp:I inn:I opbias:I out:O
XC1 net5 out sky130_fd_pr__cap_mim_m3_1 W=2 L=4 m=1
XC2 out net4 sky130_fd_pr__cap_mim_m3_1 W=2 L=4 m=1
XM26 net2 opbias VDD sky130_fd_pr__pfet_01v8_lvt L=3 W=10 nf=4 m=1
XM3 net1 net1 VDD sky130_fd_pr__pfet_01v8_lvt L=3 W=10 nf=2 m=1
XM4 net5 net1 VDD sky130_fd_pr__pfet_01v8_lvt L=3 W=10 nf=2 m=1
XM10 out net5 VDD sky130_fd_pr__pfet_01v8_lvt L=3 W=100 nf=5 m=1
XM17 out net4 GND sky130_fd_pr__nfet_01v8_lvt L=3 W=80 nf=5 m=1
XM19 net4 net3 GND sky130_fd_pr__nfet_01v8_lvt L=3 W=5 nf=1 m=1
XM20 net3 net3 GND sky130_fd_pr__nfet_01v8_lvt L=3 W=5 nf=1 m=1
XM2 net1 net4 GND GND sky130_fd_pr__nfet_01v8_lvt L=3 W=8 nf=1 m=1
XM5 net5 net3 GND GND sky130_fd_pr__nfet_01v8_lvt L=3 W=8 nf=1 m=1
XM1 net3 inn net2 sky130_fd_pr__pfet_01v8_lvt L=3 W=15 nf=3 m=1
XM6 net4 inp net2 sky130_fd_pr__pfet_01v8_lvt L=3 W=15 nf=3 m=1
.ends


* expanding   symbol:  not/not.sym # of pins=2
** sym_path: /run/media/thuat/build/cmos/MulColRO/xschem/not/not.sym
** sch_path: /run/media/thuat/build/cmos/MulColRO/xschem/not/not.sch
.subckt not out in
*.PININFO in:I out:O
XM10 out in VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=1 nf=1 m=1
XM1 out in GND GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 m=1
.ends

.GLOBAL GND
.GLOBAL VDD
.end
