magic
tech sky130A
timestamp 1695443368
<< metal1 >>
rect 0 0 100 100
rect 0 -200 100 -100
rect 0 -400 100 -300
use opamp  x1
timestamp 1695442520
transform 1 0 0 0 1 900
box 3034 622 9644 4507
<< labels >>
flabel metal1 0 0 100 100 0 FreeSans 128 0 0 0 opbias
port 0 nsew
flabel metal1 0 -200 100 -100 0 FreeSans 128 0 0 0 in
port 1 nsew
flabel metal1 0 -400 100 -300 0 FreeSans 128 0 0 0 out
port 2 nsew
<< end >>
