magic
tech sky130A
magscale 1 2
timestamp 1694848836
<< nwell >>
rect -4115 -2711 4115 2711
<< pmoslvt >>
rect -3919 -2492 -3319 2492
rect -3261 -2492 -2661 2492
rect -2603 -2492 -2003 2492
rect -1945 -2492 -1345 2492
rect -1287 -2492 -687 2492
rect -629 -2492 -29 2492
rect 29 -2492 629 2492
rect 687 -2492 1287 2492
rect 1345 -2492 1945 2492
rect 2003 -2492 2603 2492
rect 2661 -2492 3261 2492
rect 3319 -2492 3919 2492
<< pdiff >>
rect -3977 2480 -3919 2492
rect -3977 -2480 -3965 2480
rect -3931 -2480 -3919 2480
rect -3977 -2492 -3919 -2480
rect -3319 2480 -3261 2492
rect -3319 -2480 -3307 2480
rect -3273 -2480 -3261 2480
rect -3319 -2492 -3261 -2480
rect -2661 2480 -2603 2492
rect -2661 -2480 -2649 2480
rect -2615 -2480 -2603 2480
rect -2661 -2492 -2603 -2480
rect -2003 2480 -1945 2492
rect -2003 -2480 -1991 2480
rect -1957 -2480 -1945 2480
rect -2003 -2492 -1945 -2480
rect -1345 2480 -1287 2492
rect -1345 -2480 -1333 2480
rect -1299 -2480 -1287 2480
rect -1345 -2492 -1287 -2480
rect -687 2480 -629 2492
rect -687 -2480 -675 2480
rect -641 -2480 -629 2480
rect -687 -2492 -629 -2480
rect -29 2480 29 2492
rect -29 -2480 -17 2480
rect 17 -2480 29 2480
rect -29 -2492 29 -2480
rect 629 2480 687 2492
rect 629 -2480 641 2480
rect 675 -2480 687 2480
rect 629 -2492 687 -2480
rect 1287 2480 1345 2492
rect 1287 -2480 1299 2480
rect 1333 -2480 1345 2480
rect 1287 -2492 1345 -2480
rect 1945 2480 2003 2492
rect 1945 -2480 1957 2480
rect 1991 -2480 2003 2480
rect 1945 -2492 2003 -2480
rect 2603 2480 2661 2492
rect 2603 -2480 2615 2480
rect 2649 -2480 2661 2480
rect 2603 -2492 2661 -2480
rect 3261 2480 3319 2492
rect 3261 -2480 3273 2480
rect 3307 -2480 3319 2480
rect 3261 -2492 3319 -2480
rect 3919 2480 3977 2492
rect 3919 -2480 3931 2480
rect 3965 -2480 3977 2480
rect 3919 -2492 3977 -2480
<< pdiffc >>
rect -3965 -2480 -3931 2480
rect -3307 -2480 -3273 2480
rect -2649 -2480 -2615 2480
rect -1991 -2480 -1957 2480
rect -1333 -2480 -1299 2480
rect -675 -2480 -641 2480
rect -17 -2480 17 2480
rect 641 -2480 675 2480
rect 1299 -2480 1333 2480
rect 1957 -2480 1991 2480
rect 2615 -2480 2649 2480
rect 3273 -2480 3307 2480
rect 3931 -2480 3965 2480
<< nsubdiff >>
rect -4079 2641 -3983 2675
rect 3983 2641 4079 2675
rect -4079 2579 -4045 2641
rect 4045 2579 4079 2641
rect -4079 -2641 -4045 -2579
rect 4045 -2641 4079 -2579
rect -4079 -2675 -3983 -2641
rect 3983 -2675 4079 -2641
<< nsubdiffcont >>
rect -3983 2641 3983 2675
rect -4079 -2579 -4045 2579
rect 4045 -2579 4079 2579
rect -3983 -2675 3983 -2641
<< poly >>
rect -3919 2573 -3319 2589
rect -3919 2539 -3903 2573
rect -3335 2539 -3319 2573
rect -3919 2492 -3319 2539
rect -3261 2573 -2661 2589
rect -3261 2539 -3245 2573
rect -2677 2539 -2661 2573
rect -3261 2492 -2661 2539
rect -2603 2573 -2003 2589
rect -2603 2539 -2587 2573
rect -2019 2539 -2003 2573
rect -2603 2492 -2003 2539
rect -1945 2573 -1345 2589
rect -1945 2539 -1929 2573
rect -1361 2539 -1345 2573
rect -1945 2492 -1345 2539
rect -1287 2573 -687 2589
rect -1287 2539 -1271 2573
rect -703 2539 -687 2573
rect -1287 2492 -687 2539
rect -629 2573 -29 2589
rect -629 2539 -613 2573
rect -45 2539 -29 2573
rect -629 2492 -29 2539
rect 29 2573 629 2589
rect 29 2539 45 2573
rect 613 2539 629 2573
rect 29 2492 629 2539
rect 687 2573 1287 2589
rect 687 2539 703 2573
rect 1271 2539 1287 2573
rect 687 2492 1287 2539
rect 1345 2573 1945 2589
rect 1345 2539 1361 2573
rect 1929 2539 1945 2573
rect 1345 2492 1945 2539
rect 2003 2573 2603 2589
rect 2003 2539 2019 2573
rect 2587 2539 2603 2573
rect 2003 2492 2603 2539
rect 2661 2573 3261 2589
rect 2661 2539 2677 2573
rect 3245 2539 3261 2573
rect 2661 2492 3261 2539
rect 3319 2573 3919 2589
rect 3319 2539 3335 2573
rect 3903 2539 3919 2573
rect 3319 2492 3919 2539
rect -3919 -2539 -3319 -2492
rect -3919 -2573 -3903 -2539
rect -3335 -2573 -3319 -2539
rect -3919 -2589 -3319 -2573
rect -3261 -2539 -2661 -2492
rect -3261 -2573 -3245 -2539
rect -2677 -2573 -2661 -2539
rect -3261 -2589 -2661 -2573
rect -2603 -2539 -2003 -2492
rect -2603 -2573 -2587 -2539
rect -2019 -2573 -2003 -2539
rect -2603 -2589 -2003 -2573
rect -1945 -2539 -1345 -2492
rect -1945 -2573 -1929 -2539
rect -1361 -2573 -1345 -2539
rect -1945 -2589 -1345 -2573
rect -1287 -2539 -687 -2492
rect -1287 -2573 -1271 -2539
rect -703 -2573 -687 -2539
rect -1287 -2589 -687 -2573
rect -629 -2539 -29 -2492
rect -629 -2573 -613 -2539
rect -45 -2573 -29 -2539
rect -629 -2589 -29 -2573
rect 29 -2539 629 -2492
rect 29 -2573 45 -2539
rect 613 -2573 629 -2539
rect 29 -2589 629 -2573
rect 687 -2539 1287 -2492
rect 687 -2573 703 -2539
rect 1271 -2573 1287 -2539
rect 687 -2589 1287 -2573
rect 1345 -2539 1945 -2492
rect 1345 -2573 1361 -2539
rect 1929 -2573 1945 -2539
rect 1345 -2589 1945 -2573
rect 2003 -2539 2603 -2492
rect 2003 -2573 2019 -2539
rect 2587 -2573 2603 -2539
rect 2003 -2589 2603 -2573
rect 2661 -2539 3261 -2492
rect 2661 -2573 2677 -2539
rect 3245 -2573 3261 -2539
rect 2661 -2589 3261 -2573
rect 3319 -2539 3919 -2492
rect 3319 -2573 3335 -2539
rect 3903 -2573 3919 -2539
rect 3319 -2589 3919 -2573
<< polycont >>
rect -3903 2539 -3335 2573
rect -3245 2539 -2677 2573
rect -2587 2539 -2019 2573
rect -1929 2539 -1361 2573
rect -1271 2539 -703 2573
rect -613 2539 -45 2573
rect 45 2539 613 2573
rect 703 2539 1271 2573
rect 1361 2539 1929 2573
rect 2019 2539 2587 2573
rect 2677 2539 3245 2573
rect 3335 2539 3903 2573
rect -3903 -2573 -3335 -2539
rect -3245 -2573 -2677 -2539
rect -2587 -2573 -2019 -2539
rect -1929 -2573 -1361 -2539
rect -1271 -2573 -703 -2539
rect -613 -2573 -45 -2539
rect 45 -2573 613 -2539
rect 703 -2573 1271 -2539
rect 1361 -2573 1929 -2539
rect 2019 -2573 2587 -2539
rect 2677 -2573 3245 -2539
rect 3335 -2573 3903 -2539
<< locali >>
rect -4079 2641 -3983 2675
rect 3983 2641 4079 2675
rect -4079 2579 -4045 2641
rect 4045 2579 4079 2641
rect -3919 2539 -3903 2573
rect -3335 2539 -3319 2573
rect -3261 2539 -3245 2573
rect -2677 2539 -2661 2573
rect -2603 2539 -2587 2573
rect -2019 2539 -2003 2573
rect -1945 2539 -1929 2573
rect -1361 2539 -1345 2573
rect -1287 2539 -1271 2573
rect -703 2539 -687 2573
rect -629 2539 -613 2573
rect -45 2539 -29 2573
rect 29 2539 45 2573
rect 613 2539 629 2573
rect 687 2539 703 2573
rect 1271 2539 1287 2573
rect 1345 2539 1361 2573
rect 1929 2539 1945 2573
rect 2003 2539 2019 2573
rect 2587 2539 2603 2573
rect 2661 2539 2677 2573
rect 3245 2539 3261 2573
rect 3319 2539 3335 2573
rect 3903 2539 3919 2573
rect -3965 2480 -3931 2496
rect -3965 -2496 -3931 -2480
rect -3307 2480 -3273 2496
rect -3307 -2496 -3273 -2480
rect -2649 2480 -2615 2496
rect -2649 -2496 -2615 -2480
rect -1991 2480 -1957 2496
rect -1991 -2496 -1957 -2480
rect -1333 2480 -1299 2496
rect -1333 -2496 -1299 -2480
rect -675 2480 -641 2496
rect -675 -2496 -641 -2480
rect -17 2480 17 2496
rect -17 -2496 17 -2480
rect 641 2480 675 2496
rect 641 -2496 675 -2480
rect 1299 2480 1333 2496
rect 1299 -2496 1333 -2480
rect 1957 2480 1991 2496
rect 1957 -2496 1991 -2480
rect 2615 2480 2649 2496
rect 2615 -2496 2649 -2480
rect 3273 2480 3307 2496
rect 3273 -2496 3307 -2480
rect 3931 2480 3965 2496
rect 3931 -2496 3965 -2480
rect -3919 -2573 -3903 -2539
rect -3335 -2573 -3319 -2539
rect -3261 -2573 -3245 -2539
rect -2677 -2573 -2661 -2539
rect -2603 -2573 -2587 -2539
rect -2019 -2573 -2003 -2539
rect -1945 -2573 -1929 -2539
rect -1361 -2573 -1345 -2539
rect -1287 -2573 -1271 -2539
rect -703 -2573 -687 -2539
rect -629 -2573 -613 -2539
rect -45 -2573 -29 -2539
rect 29 -2573 45 -2539
rect 613 -2573 629 -2539
rect 687 -2573 703 -2539
rect 1271 -2573 1287 -2539
rect 1345 -2573 1361 -2539
rect 1929 -2573 1945 -2539
rect 2003 -2573 2019 -2539
rect 2587 -2573 2603 -2539
rect 2661 -2573 2677 -2539
rect 3245 -2573 3261 -2539
rect 3319 -2573 3335 -2539
rect 3903 -2573 3919 -2539
rect -4079 -2641 -4045 -2579
rect 4045 -2641 4079 -2579
rect -4079 -2675 -3983 -2641
rect 3983 -2675 4079 -2641
<< viali >>
rect -3903 2539 -3335 2573
rect -3245 2539 -2677 2573
rect -2587 2539 -2019 2573
rect -1929 2539 -1361 2573
rect -1271 2539 -703 2573
rect -613 2539 -45 2573
rect 45 2539 613 2573
rect 703 2539 1271 2573
rect 1361 2539 1929 2573
rect 2019 2539 2587 2573
rect 2677 2539 3245 2573
rect 3335 2539 3903 2573
rect -3965 -2480 -3931 2480
rect -3307 -2480 -3273 2480
rect -2649 -2480 -2615 2480
rect -1991 -2480 -1957 2480
rect -1333 -2480 -1299 2480
rect -675 -2480 -641 2480
rect -17 -2480 17 2480
rect 641 -2480 675 2480
rect 1299 -2480 1333 2480
rect 1957 -2480 1991 2480
rect 2615 -2480 2649 2480
rect 3273 -2480 3307 2480
rect 3931 -2480 3965 2480
rect -3903 -2573 -3335 -2539
rect -3245 -2573 -2677 -2539
rect -2587 -2573 -2019 -2539
rect -1929 -2573 -1361 -2539
rect -1271 -2573 -703 -2539
rect -613 -2573 -45 -2539
rect 45 -2573 613 -2539
rect 703 -2573 1271 -2539
rect 1361 -2573 1929 -2539
rect 2019 -2573 2587 -2539
rect 2677 -2573 3245 -2539
rect 3335 -2573 3903 -2539
<< metal1 >>
rect -3915 2573 -3323 2579
rect -3915 2539 -3903 2573
rect -3335 2539 -3323 2573
rect -3915 2533 -3323 2539
rect -3257 2573 -2665 2579
rect -3257 2539 -3245 2573
rect -2677 2539 -2665 2573
rect -3257 2533 -2665 2539
rect -2599 2573 -2007 2579
rect -2599 2539 -2587 2573
rect -2019 2539 -2007 2573
rect -2599 2533 -2007 2539
rect -1941 2573 -1349 2579
rect -1941 2539 -1929 2573
rect -1361 2539 -1349 2573
rect -1941 2533 -1349 2539
rect -1283 2573 -691 2579
rect -1283 2539 -1271 2573
rect -703 2539 -691 2573
rect -1283 2533 -691 2539
rect -625 2573 -33 2579
rect -625 2539 -613 2573
rect -45 2539 -33 2573
rect -625 2533 -33 2539
rect 33 2573 625 2579
rect 33 2539 45 2573
rect 613 2539 625 2573
rect 33 2533 625 2539
rect 691 2573 1283 2579
rect 691 2539 703 2573
rect 1271 2539 1283 2573
rect 691 2533 1283 2539
rect 1349 2573 1941 2579
rect 1349 2539 1361 2573
rect 1929 2539 1941 2573
rect 1349 2533 1941 2539
rect 2007 2573 2599 2579
rect 2007 2539 2019 2573
rect 2587 2539 2599 2573
rect 2007 2533 2599 2539
rect 2665 2573 3257 2579
rect 2665 2539 2677 2573
rect 3245 2539 3257 2573
rect 2665 2533 3257 2539
rect 3323 2573 3915 2579
rect 3323 2539 3335 2573
rect 3903 2539 3915 2573
rect 3323 2533 3915 2539
rect -3971 2480 -3925 2492
rect -3971 -2480 -3965 2480
rect -3931 -2480 -3925 2480
rect -3971 -2492 -3925 -2480
rect -3313 2480 -3267 2492
rect -3313 -2480 -3307 2480
rect -3273 -2480 -3267 2480
rect -3313 -2492 -3267 -2480
rect -2655 2480 -2609 2492
rect -2655 -2480 -2649 2480
rect -2615 -2480 -2609 2480
rect -2655 -2492 -2609 -2480
rect -1997 2480 -1951 2492
rect -1997 -2480 -1991 2480
rect -1957 -2480 -1951 2480
rect -1997 -2492 -1951 -2480
rect -1339 2480 -1293 2492
rect -1339 -2480 -1333 2480
rect -1299 -2480 -1293 2480
rect -1339 -2492 -1293 -2480
rect -681 2480 -635 2492
rect -681 -2480 -675 2480
rect -641 -2480 -635 2480
rect -681 -2492 -635 -2480
rect -23 2480 23 2492
rect -23 -2480 -17 2480
rect 17 -2480 23 2480
rect -23 -2492 23 -2480
rect 635 2480 681 2492
rect 635 -2480 641 2480
rect 675 -2480 681 2480
rect 635 -2492 681 -2480
rect 1293 2480 1339 2492
rect 1293 -2480 1299 2480
rect 1333 -2480 1339 2480
rect 1293 -2492 1339 -2480
rect 1951 2480 1997 2492
rect 1951 -2480 1957 2480
rect 1991 -2480 1997 2480
rect 1951 -2492 1997 -2480
rect 2609 2480 2655 2492
rect 2609 -2480 2615 2480
rect 2649 -2480 2655 2480
rect 2609 -2492 2655 -2480
rect 3267 2480 3313 2492
rect 3267 -2480 3273 2480
rect 3307 -2480 3313 2480
rect 3267 -2492 3313 -2480
rect 3925 2480 3971 2492
rect 3925 -2480 3931 2480
rect 3965 -2480 3971 2480
rect 3925 -2492 3971 -2480
rect -3915 -2539 -3323 -2533
rect -3915 -2573 -3903 -2539
rect -3335 -2573 -3323 -2539
rect -3915 -2579 -3323 -2573
rect -3257 -2539 -2665 -2533
rect -3257 -2573 -3245 -2539
rect -2677 -2573 -2665 -2539
rect -3257 -2579 -2665 -2573
rect -2599 -2539 -2007 -2533
rect -2599 -2573 -2587 -2539
rect -2019 -2573 -2007 -2539
rect -2599 -2579 -2007 -2573
rect -1941 -2539 -1349 -2533
rect -1941 -2573 -1929 -2539
rect -1361 -2573 -1349 -2539
rect -1941 -2579 -1349 -2573
rect -1283 -2539 -691 -2533
rect -1283 -2573 -1271 -2539
rect -703 -2573 -691 -2539
rect -1283 -2579 -691 -2573
rect -625 -2539 -33 -2533
rect -625 -2573 -613 -2539
rect -45 -2573 -33 -2539
rect -625 -2579 -33 -2573
rect 33 -2539 625 -2533
rect 33 -2573 45 -2539
rect 613 -2573 625 -2539
rect 33 -2579 625 -2573
rect 691 -2539 1283 -2533
rect 691 -2573 703 -2539
rect 1271 -2573 1283 -2539
rect 691 -2579 1283 -2573
rect 1349 -2539 1941 -2533
rect 1349 -2573 1361 -2539
rect 1929 -2573 1941 -2539
rect 1349 -2579 1941 -2573
rect 2007 -2539 2599 -2533
rect 2007 -2573 2019 -2539
rect 2587 -2573 2599 -2539
rect 2007 -2579 2599 -2573
rect 2665 -2539 3257 -2533
rect 2665 -2573 2677 -2539
rect 3245 -2573 3257 -2539
rect 2665 -2579 3257 -2573
rect 3323 -2539 3915 -2533
rect 3323 -2573 3335 -2539
rect 3903 -2573 3915 -2539
rect 3323 -2579 3915 -2573
<< properties >>
string FIXED_BBOX -4062 -2658 4062 2658
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 24.916666666666668 l 3.0 m 1 nf 12 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
