magic
tech sky130A
magscale 1 2
timestamp 1698935188
<< locali >>
rect 3416 8344 3884 8346
rect 3416 7934 4444 8344
rect 3416 7762 4214 7934
rect 4388 7762 4444 7934
rect 3416 7238 4444 7762
rect 3416 7226 3884 7238
rect 3547 7216 3884 7226
rect 5014 168 8602 662
rect 5014 -552 5960 168
rect 7596 -552 8602 168
rect 5014 -748 8602 -552
<< viali >>
rect 4214 7762 4388 7934
rect 5960 -552 7596 168
<< metal1 >>
rect -40 9086 8604 10274
rect 3594 8810 3772 8820
rect 2718 8734 3772 8810
rect 2656 7862 2772 8090
rect 2656 7630 2672 7862
rect 2764 7630 2772 7862
rect 2656 7432 2772 7630
rect 2918 7854 3034 8088
rect 2918 7622 2926 7854
rect 3018 7622 3034 7854
rect 2918 7430 3034 7622
rect 3168 7854 3284 8076
rect 3168 7622 3182 7854
rect 3274 7622 3284 7854
rect 3168 7418 3284 7622
rect 3594 4686 3772 8734
rect 4202 7934 4402 7948
rect 4202 7762 4214 7934
rect 4388 7762 4402 7934
rect 4202 7748 4402 7762
rect 4802 5398 4940 9086
rect 5300 4928 5748 8890
rect 5782 7838 5918 8204
rect 5782 7380 5800 7838
rect 5892 7380 5918 7838
rect 5782 7100 5918 7380
rect 2788 1862 2902 2104
rect 2788 1634 2796 1862
rect 2896 1634 2902 1862
rect 2788 1422 2902 1634
rect 3048 1858 3162 2088
rect 3048 1630 3052 1858
rect 3152 1630 3162 1858
rect 3048 1406 3162 1630
rect 3306 1846 3420 2072
rect 3306 1618 3316 1846
rect 3416 1618 3420 1846
rect 3306 1390 3420 1618
rect 3596 662 3754 4686
rect 5300 4480 5412 4928
rect 5624 4480 5748 4928
rect 4228 3404 4428 3444
rect 4228 3282 4284 3404
rect 4402 3282 4428 3404
rect 4228 3244 4428 3282
rect 4238 1818 4438 1844
rect 4238 1664 4264 1818
rect 4418 1664 4438 1818
rect 4238 1644 4438 1664
rect 2714 606 3754 662
rect 3596 602 3754 606
rect 4804 430 4942 4464
rect 5132 2164 5240 2478
rect 5132 1510 5152 2164
rect 5226 1510 5240 2164
rect 5132 1076 5240 1510
rect 5300 696 5748 4480
rect 5952 4924 6400 8894
rect 5952 4476 6078 4924
rect 6290 4476 6400 4924
rect 5952 994 6400 4476
rect 6610 4928 7058 8890
rect 7102 7810 7238 8186
rect 7102 7352 7118 7810
rect 7210 7352 7238 7810
rect 7102 7082 7238 7352
rect 6610 4480 6726 4928
rect 6938 4480 7058 4928
rect 6442 2136 6550 2484
rect 6442 1482 6466 2136
rect 6540 1482 6550 2136
rect 6442 1082 6550 1482
rect 5952 708 6402 994
rect 6610 696 7058 4480
rect 7274 4922 7722 8878
rect 7274 4474 7394 4922
rect 7606 4474 7722 4922
rect 7274 684 7722 4474
rect 7926 4910 8374 8884
rect 8410 7798 8546 8188
rect 8410 7340 8434 7798
rect 8526 7340 8546 7798
rect 8410 7084 8546 7340
rect 7926 4462 8038 4910
rect 8250 4462 8374 4910
rect 7764 2128 7872 2448
rect 7764 1474 7782 2128
rect 7856 1474 7872 2128
rect 7764 1046 7872 1474
rect 7926 690 8374 4462
rect -30 168 8632 430
rect -30 -552 5960 168
rect 7596 -552 8632 168
rect -30 -918 8632 -552
<< via1 >>
rect 2672 7630 2764 7862
rect 2926 7622 3018 7854
rect 3182 7622 3274 7854
rect 4238 7784 4374 7920
rect 5800 7380 5892 7838
rect 2796 1634 2896 1862
rect 3052 1630 3152 1858
rect 3316 1618 3416 1846
rect 5412 4480 5624 4928
rect 4284 3282 4402 3404
rect 4264 1664 4418 1818
rect 5152 1510 5226 2164
rect 6078 4476 6290 4924
rect 7118 7352 7210 7810
rect 6726 4480 6938 4928
rect 6466 1482 6540 2136
rect 7394 4474 7606 4922
rect 8434 7340 8526 7798
rect 8038 4462 8250 4910
rect 7782 1474 7856 2128
<< metal2 >>
rect 5116 8352 8552 8740
rect 3844 8350 8552 8352
rect 2532 7920 8552 8350
rect 2532 7862 4238 7920
rect 2532 7630 2672 7862
rect 2764 7854 4238 7862
rect 2764 7630 2926 7854
rect 2532 7622 2926 7630
rect 3018 7622 3182 7854
rect 3274 7784 4238 7854
rect 4374 7838 8552 7920
rect 4374 7784 5800 7838
rect 3274 7622 5800 7784
rect 2532 7380 5800 7622
rect 5892 7810 8552 7838
rect 5892 7380 7118 7810
rect 2532 7352 7118 7380
rect 7210 7798 8552 7810
rect 7210 7352 8434 7798
rect 2532 7340 8434 7352
rect 8526 7340 8552 7798
rect 2532 7226 8552 7340
rect 2532 7224 4188 7226
rect 3547 7218 4188 7224
rect 3688 7216 3752 7218
rect 5116 6794 8552 7226
rect 5126 4928 8544 5168
rect 5126 4914 5412 4928
rect 4744 4684 5412 4914
rect 5126 4480 5412 4684
rect 5624 4924 6726 4928
rect 5624 4480 6078 4924
rect 5126 4476 6078 4480
rect 6290 4480 6726 4924
rect 6938 4922 8544 4928
rect 6938 4480 7394 4922
rect 6290 4476 7394 4480
rect 5126 4474 7394 4476
rect 7606 4910 8544 4922
rect 7606 4474 8038 4910
rect 5126 4462 8038 4474
rect 8250 4462 8544 4910
rect 5126 4254 8544 4462
rect 5126 3474 5310 4254
rect 4218 3404 5310 3474
rect 4218 3282 4284 3404
rect 4402 3282 5310 3404
rect 4218 3220 5310 3282
rect 4218 3216 5270 3220
rect 5112 2336 8548 2746
rect 3844 2332 8548 2336
rect 2574 2164 8548 2332
rect 2574 1862 5152 2164
rect 2574 1634 2796 1862
rect 2896 1858 5152 1862
rect 2896 1634 3052 1858
rect 2574 1630 3052 1634
rect 3152 1846 5152 1858
rect 3152 1630 3316 1846
rect 2574 1618 3316 1630
rect 3416 1818 5152 1846
rect 3416 1664 4264 1818
rect 4418 1664 5152 1818
rect 3416 1618 5152 1664
rect 2574 1510 5152 1618
rect 5226 2136 8548 2164
rect 5226 1510 6466 2136
rect 2574 1482 6466 1510
rect 6540 2128 8548 2136
rect 6540 1482 7782 2128
rect 2574 1474 7782 1482
rect 7856 1474 8548 2128
rect 2574 1210 8548 1474
rect 2574 1206 4066 1210
rect 3547 1202 4066 1206
rect 3688 1200 3752 1202
rect 5112 808 8548 1210
rect 5112 800 5802 808
rect 6520 800 8548 808
use not  x1
timestamp 1696661316
transform -1 0 5462 0 1 4624
box 472 -578 1868 1036
use sky130_fd_pr__nfet_01v8_lvt_4833E6  XM1
timestamp 1696133064
transform 1 0 6830 0 1 4780
box -1812 -4210 1812 4210
use sky130_fd_pr__pfet_01v8_lvt_ER7S26  XM26
timestamp 1698123815
transform 1 0 3037 0 1 4695
box -487 -4219 487 4219
<< labels >>
flabel metal2 4202 7748 4402 7948 0 FreeSans 256 0 0 0 out
port 1 nsew
rlabel via1 4284 3282 4402 3404 1 toggle
port 6 nsew
rlabel metal1 -40 9086 8604 10274 1 VDD
port 4 nsew
flabel metal2 4238 1644 4438 1844 0 FreeSans 256 0 0 0 in
port 2 nsew
rlabel metal1 -30 -918 8632 430 1 VSS
port 7 nsew
<< end >>
