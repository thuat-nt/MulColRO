magic
tech sky130A
magscale 1 2
timestamp 1695461589
<< checkpaint >>
rect 12333 -543 234983 59941
<< error_p >>
rect 115397 52856 115431 53230
rect 118143 49942 118177 53230
rect 118915 52856 118949 53230
rect 120468 52856 120502 53230
rect 123986 52856 124020 53230
rect 115397 49635 115431 49942
rect 115511 49731 115545 49765
rect 116169 49731 116203 49765
rect 116827 49731 116861 49765
rect 117485 49731 117519 49765
rect 118143 49731 118177 49765
rect 118801 49731 118855 49765
rect 115461 49697 115465 49731
rect 115477 49697 118855 49731
rect 46574 46520 46576 46570
rect 46602 46520 46604 46598
rect 46022 46280 46660 46520
rect 51788 46476 51790 46554
rect 51816 46476 51818 46526
rect 51732 46236 52370 46476
rect 46556 45974 46576 46094
rect 46584 45968 46604 46122
rect 51788 45924 51808 46078
rect 51816 45930 51836 46050
rect 42488 45306 43970 45418
rect 41048 45272 47214 45306
rect 42488 44648 43970 45272
rect 41048 44614 47214 44648
rect 42488 43990 43970 44614
rect 41048 43956 47214 43990
rect 42488 43842 43970 43956
rect 47264 43344 47298 43362
rect 47230 43310 47332 43328
rect 57706 42722 57762 42744
rect 68795 42667 68829 49031
rect 70225 45418 70259 48932
rect 70883 45418 70917 48932
rect 69888 45126 71370 45418
rect 69804 44678 71370 45126
rect 69888 44484 71370 44678
rect 71541 44484 71575 48932
rect 69888 44112 71942 44484
rect 69888 43842 71370 44112
rect 68909 42763 68943 42797
rect 69567 42763 69601 42797
rect 70225 42763 70259 43842
rect 70883 42763 70917 43842
rect 71541 42763 71575 44112
rect 72199 42763 72253 42797
rect 68859 42729 68863 42763
rect 68875 42729 72253 42763
rect 70225 42708 70259 42729
rect 70883 42708 70917 42729
rect 71541 42708 71575 42729
rect 51178 42596 59154 42630
rect 57706 42496 57762 42518
rect 50992 41824 59340 41844
rect 68763 41826 68829 42667
rect 68897 42661 71798 42708
rect 72139 42661 72186 42708
rect 68909 42627 69554 42661
rect 69567 42627 70212 42661
rect 70225 42627 70870 42661
rect 70883 42627 71528 42661
rect 71541 42627 72186 42661
rect 68909 42580 68955 42627
rect 68865 42568 68883 42580
rect 68909 42568 68954 42580
rect 68865 41826 68954 42568
rect 68966 41826 68984 42621
rect 68994 41826 69012 42621
rect 69567 42580 69613 42627
rect 70156 42621 70177 42627
rect 70184 42593 70205 42627
rect 70225 42580 70271 42627
rect 69524 42568 69555 42579
rect 69567 42568 69612 42580
rect 70182 42568 70213 42579
rect 70225 42568 70270 42580
rect 69464 42012 69474 42302
rect 69436 41826 69474 42012
rect 69492 41826 69502 42274
rect 69535 41826 69612 42568
rect 70193 41826 70270 42568
rect 70286 41956 70292 42621
rect 70314 41956 70320 42621
rect 70883 42580 70929 42627
rect 71476 42621 71493 42627
rect 71504 42593 71521 42627
rect 71541 42580 71587 42627
rect 70840 42568 70871 42579
rect 70883 42568 70928 42580
rect 71498 42568 71529 42579
rect 71541 42568 71586 42580
rect 70774 41956 70794 42308
rect 70802 41956 70822 42280
rect 70851 41826 70928 42568
rect 71509 41826 71586 42568
rect 71608 41956 71612 42621
rect 71636 41956 71640 42621
rect 72156 42568 72187 42579
rect 72199 42568 72233 42729
rect 54398 41752 54684 41772
rect 54432 41718 54650 41738
rect 54188 41654 54856 41688
rect 55704 41654 56372 41688
rect 44996 41618 45098 41644
rect 45754 41618 45856 41644
rect 46512 41618 46614 41644
rect 47270 41618 47372 41644
rect 45024 41590 45070 41616
rect 45782 41590 45828 41616
rect 46540 41590 46586 41616
rect 47298 41590 47344 41616
rect 54758 41354 54784 41532
rect 54786 41354 54812 41532
rect 55070 41514 55152 41530
rect 55260 41514 55300 41530
rect 55608 41408 55622 41570
rect 55636 41408 55650 41570
rect 54610 41320 55158 41354
rect 54610 41038 54644 41320
rect 54758 41246 54784 41320
rect 54786 41246 54812 41320
rect 54884 41240 54918 41320
rect 54972 41240 54983 41251
rect 54674 41196 54746 41234
rect 54796 41206 54983 41240
rect 54712 41162 54746 41196
rect 54871 41194 54872 41195
rect 54872 41193 54873 41194
rect 54872 41164 54873 41165
rect 54871 41163 54872 41164
rect 54884 41152 54918 41206
rect 54984 41196 55056 41234
rect 54930 41194 54931 41195
rect 54929 41193 54930 41194
rect 54929 41164 54930 41165
rect 54930 41163 54931 41164
rect 54972 41152 54983 41163
rect 55022 41162 55056 41196
rect 54796 41118 54983 41152
rect 54766 41038 54784 41112
rect 54794 41038 54812 41112
rect 54884 41038 54918 41118
rect 55124 41038 55158 41320
rect 54610 41004 55158 41038
rect 54766 40950 54784 41004
rect 54764 40796 54784 40950
rect 54794 40922 54812 41004
rect 55208 40946 55846 41408
rect 54792 40824 54812 40922
rect 55608 40824 55616 40946
rect 55636 40796 55644 40946
rect 44880 36893 47459 40385
rect 50933 36893 59371 40341
rect 60948 37056 60982 41604
rect 68308 40988 68366 41008
rect 68328 40569 68329 40988
rect 68366 40569 68386 40988
rect 68328 40568 68386 40569
rect 68727 40897 71744 41826
rect 72096 40903 72116 42278
rect 72124 41956 72144 42250
rect 72167 41956 72233 42568
rect 72124 40956 72233 41956
rect 72281 42667 72299 42729
rect 72313 42667 72347 49031
rect 73866 42672 73900 49036
rect 73980 42768 74014 42802
rect 74638 42768 74672 42802
rect 75296 42768 75330 42802
rect 75954 42768 75988 42802
rect 76612 42768 76646 42802
rect 77270 42768 77324 42802
rect 73930 42734 73934 42768
rect 73946 42734 77324 42768
rect 72281 41826 72347 42667
rect 72124 40944 72201 40956
rect 72124 40903 72213 40944
rect 72155 40897 72213 40903
rect 68727 40863 72213 40897
rect 68727 40795 71744 40863
rect 72155 40847 72201 40863
rect 72161 40795 72172 40847
rect 68727 40761 72213 40795
rect 44880 36870 59371 36893
rect 44880 36834 47459 36870
rect 50933 36834 59371 36870
rect 68727 36834 71744 40761
rect 72280 40725 72383 41826
rect 73834 41790 73900 42672
rect 73976 42666 74616 42704
rect 74634 42666 75274 42704
rect 75292 42666 75932 42704
rect 75950 42666 76590 42704
rect 76608 42666 77248 42704
rect 73980 42632 74616 42666
rect 74638 42662 75274 42666
rect 74638 42632 75276 42662
rect 73980 42594 74026 42632
rect 74638 42594 74684 42632
rect 75226 42626 75248 42632
rect 75254 42598 75276 42632
rect 75296 42632 75932 42666
rect 75954 42632 76590 42666
rect 76612 42632 77248 42666
rect 75296 42594 75342 42632
rect 75954 42594 76000 42632
rect 76548 42626 76564 42632
rect 76576 42598 76592 42626
rect 76612 42594 76658 42632
rect 73936 42582 73954 42594
rect 73980 42582 74025 42594
rect 74595 42582 74626 42593
rect 74638 42582 74683 42594
rect 75253 42582 75284 42593
rect 75296 42582 75341 42594
rect 75911 42582 75942 42593
rect 75954 42582 75999 42594
rect 76569 42582 76600 42593
rect 76612 42582 76657 42594
rect 73936 41790 74025 42582
rect 74534 41790 74560 42046
rect 74562 41790 74588 42018
rect 74606 41790 74683 42582
rect 75264 41790 75341 42582
rect 75854 41790 75870 42028
rect 75882 41790 75898 42000
rect 75922 41790 75999 42582
rect 76580 41790 76657 42582
rect 76678 41790 76684 42626
rect 76706 41790 76712 42626
rect 77227 42582 77258 42593
rect 77270 42582 77304 42734
rect 77162 41790 77186 42030
rect 77190 41790 77214 42002
rect 77238 41790 77304 42582
rect 77352 42672 77370 42734
rect 77384 42672 77418 49036
rect 115365 47825 115431 49635
rect 115507 49645 115511 49663
rect 115507 49629 115557 49645
rect 115568 49635 115586 49650
rect 115596 49635 115614 49648
rect 116109 49629 116156 49676
rect 116165 49645 116169 49663
rect 116165 49629 116215 49645
rect 116767 49635 116814 49676
rect 116758 49629 116814 49635
rect 116823 49645 116827 49663
rect 116823 49629 116873 49645
rect 116888 49635 116894 49638
rect 116916 49635 116922 49648
rect 117425 49629 117472 49676
rect 117481 49645 117485 49663
rect 117481 49629 117531 49645
rect 118083 49635 118130 49676
rect 118078 49629 118130 49635
rect 118139 49645 118143 49663
rect 118139 49629 118189 49645
rect 118741 49629 118788 49676
rect 115511 49595 116156 49629
rect 116169 49595 116814 49629
rect 116827 49595 117472 49629
rect 117485 49595 118130 49629
rect 118143 49595 118788 49629
rect 115511 49548 115557 49595
rect 115467 49536 115485 49548
rect 115511 49536 115545 49548
rect 115467 47924 115545 49536
rect 115568 48248 115586 49589
rect 115596 48220 115614 49589
rect 116169 49548 116215 49595
rect 116758 49589 116779 49595
rect 116786 49561 116807 49595
rect 116827 49548 116873 49595
rect 116126 49536 116157 49547
rect 116169 49536 116203 49548
rect 116784 49536 116815 49547
rect 116827 49536 116861 49548
rect 115365 46016 115399 47825
rect 115467 47763 115513 47924
rect 116066 47871 116076 49270
rect 116094 47899 116104 49242
rect 116137 47924 116203 49536
rect 116795 47924 116861 49536
rect 116888 48236 116894 49589
rect 116916 48208 116922 49589
rect 117485 49548 117531 49595
rect 118078 49589 118095 49595
rect 118106 49561 118123 49595
rect 118143 49548 118189 49595
rect 117442 49536 117473 49547
rect 117485 49536 117519 49548
rect 118100 49536 118131 49547
rect 118143 49536 118177 49548
rect 116137 47912 116171 47924
rect 116795 47912 116829 47924
rect 116125 47899 116184 47912
rect 116094 47890 116184 47899
rect 116191 47890 116222 47899
rect 116125 47871 116184 47890
rect 116066 47865 116184 47871
rect 115573 47831 116184 47865
rect 116219 47865 116250 47871
rect 116783 47865 116842 47912
rect 117376 47871 117396 49276
rect 117404 47899 117424 49248
rect 117453 47924 117519 49536
rect 118111 47924 118177 49536
rect 118210 48214 118214 49589
rect 118238 48186 118242 49589
rect 118758 49536 118789 49547
rect 118801 49536 118835 49697
rect 117453 47912 117487 47924
rect 118111 47912 118145 47924
rect 117441 47899 117500 47912
rect 117404 47896 117500 47899
rect 117507 47896 117532 47899
rect 117441 47871 117500 47896
rect 117376 47868 117500 47871
rect 117535 47868 117560 47871
rect 117441 47865 117500 47868
rect 118099 47865 118158 47912
rect 118698 47871 118718 49246
rect 118726 47871 118746 49218
rect 118769 47924 118835 49536
rect 118883 49635 118901 49697
rect 118915 49635 118949 49942
rect 120468 49640 120502 49942
rect 120582 49736 120616 49770
rect 121240 49736 121274 49770
rect 121898 49736 121932 49770
rect 122556 49736 122590 49770
rect 123214 49736 123248 49770
rect 123872 49736 123926 49770
rect 120532 49702 120536 49736
rect 120548 49702 123926 49736
rect 118769 47912 118803 47924
rect 118757 47865 118815 47912
rect 116219 47862 116842 47865
rect 116231 47831 116842 47862
rect 116889 47831 117500 47865
rect 117547 47831 118158 47865
rect 118205 47831 118815 47865
rect 116125 47815 116171 47831
rect 116783 47815 116829 47831
rect 117441 47815 117487 47831
rect 118099 47815 118145 47831
rect 118757 47815 118803 47831
rect 118883 47825 118949 49635
rect 120436 47848 120502 49640
rect 120578 49650 120582 49668
rect 120578 49634 120628 49650
rect 121180 49634 121218 49672
rect 121236 49650 121240 49668
rect 121236 49634 121286 49650
rect 121838 49640 121876 49672
rect 121828 49634 121876 49640
rect 121894 49650 121898 49668
rect 121894 49634 121944 49650
rect 122496 49634 122534 49672
rect 122552 49650 122556 49668
rect 122552 49634 122602 49650
rect 123154 49634 123192 49672
rect 123210 49650 123214 49668
rect 123210 49634 123260 49650
rect 123812 49634 123850 49672
rect 120582 49600 121218 49634
rect 121240 49630 121876 49634
rect 121240 49600 121878 49630
rect 120582 49562 120628 49600
rect 121240 49562 121286 49600
rect 121828 49594 121850 49600
rect 121856 49566 121878 49600
rect 121898 49600 122534 49634
rect 122556 49600 123192 49634
rect 123214 49600 123850 49634
rect 121898 49562 121944 49600
rect 122556 49562 122602 49600
rect 123150 49594 123166 49600
rect 123178 49566 123194 49594
rect 123214 49562 123260 49600
rect 120538 49550 120556 49562
rect 120582 49550 120616 49562
rect 121197 49550 121228 49561
rect 121240 49550 121274 49562
rect 121855 49550 121886 49561
rect 121898 49550 121932 49562
rect 122513 49550 122544 49561
rect 122556 49550 122590 49562
rect 123171 49550 123202 49561
rect 123214 49550 123248 49562
rect 120538 47938 120616 49550
rect 118111 47763 118145 47815
rect 115467 47729 118815 47763
rect 118111 46016 118145 47729
rect 118883 46016 118917 47825
rect 115365 45978 118917 46016
rect 93198 45118 93204 45130
rect 93390 45118 93398 45130
rect 93170 45090 93204 45102
rect 93390 45090 93426 45102
rect 92660 44666 93226 44700
rect 92660 44571 92694 44666
rect 93031 44586 93042 44597
rect 92855 44583 93042 44586
rect 92855 44571 93031 44583
rect 93192 44571 93226 44666
rect 92626 44537 93226 44571
rect 92660 44344 92694 44537
rect 92715 44525 92843 44537
rect 93043 44525 93140 44537
rect 92715 44524 92796 44525
rect 93043 44524 93124 44525
rect 92762 44486 92796 44524
rect 93090 44486 93124 44524
rect 92752 44460 92804 44472
rect 93031 44458 93042 44469
rect 92724 44432 92832 44444
rect 92855 44424 93042 44458
rect 93176 44444 93178 44531
rect 93192 44344 93226 44537
rect 92660 44310 93226 44344
rect 93276 44509 93896 44714
rect 98034 44512 98164 44533
rect 93276 44292 93923 44509
rect 97848 44487 98164 44512
rect 98350 44487 98756 44533
rect 97876 44459 98164 44484
rect 98350 44459 98700 44484
rect 93889 44238 93923 44292
rect 92660 44190 93226 44224
rect 92660 43902 92694 44190
rect 93031 44110 93042 44121
rect 92715 44048 92796 44095
rect 92855 44076 93042 44110
rect 93043 44048 93124 44095
rect 92762 44010 92796 44048
rect 93090 44010 93124 44048
rect 93192 43996 93226 44190
rect 93031 43982 93042 43993
rect 93158 43982 93178 43996
rect 92855 43948 93042 43982
rect 93082 43968 93178 43982
rect 93186 43982 93226 43996
rect 93276 44086 93923 44238
rect 93276 44000 93978 44086
rect 93276 43982 93923 44000
rect 93186 43962 93923 43982
rect 93192 43954 93226 43962
rect 93276 43954 93923 43962
rect 93054 43941 93923 43954
rect 93054 43940 93896 43941
rect 93158 43934 93896 43940
rect 92817 43910 93069 43913
rect 93192 43902 93226 43934
rect 92660 43879 93226 43902
rect 92660 43868 92694 43879
rect 93192 43868 93226 43879
rect 92660 43867 93226 43868
rect 92694 43853 93192 43867
rect 92660 43834 93226 43853
rect 93276 43816 93896 43934
rect 97658 43918 98278 44340
rect 98328 44292 98894 44326
rect 98328 43970 98362 44292
rect 98699 44212 98710 44223
rect 98383 44150 98464 44197
rect 98523 44178 98710 44212
rect 98711 44150 98792 44197
rect 98430 44112 98464 44150
rect 98758 44112 98792 44150
rect 98699 44084 98710 44095
rect 98523 44050 98710 44084
rect 98860 43970 98894 44292
rect 98328 43936 98894 43970
rect 97716 43864 97734 43903
rect 98034 43875 98064 43910
rect 98090 43875 98092 43910
rect 97750 43864 97768 43869
rect 97658 43818 98278 43864
rect 98390 43850 98832 43884
rect 98328 43823 98894 43850
rect 97658 43816 98338 43818
rect 97658 43802 98396 43816
rect 97658 43790 98278 43802
rect 97658 43788 98310 43790
rect 97658 43755 98368 43788
rect 97658 43721 101528 43755
rect 97658 43685 98278 43721
rect 98328 43588 98368 43721
rect 98376 43594 98396 43714
rect 98430 43687 98464 43690
rect 98758 43687 98792 43690
rect 98328 43556 98362 43588
rect 98860 43556 98894 43721
rect 77352 41790 77418 42672
rect 78278 41826 78518 42162
rect 77802 41790 78264 41826
rect 72412 41756 78264 41790
rect 73834 40818 73900 41756
rect 73936 41752 74025 41756
rect 73914 41688 73930 41694
rect 73936 41688 74014 41752
rect 74534 41694 74560 41756
rect 74562 41694 74588 41756
rect 74606 41752 74683 41756
rect 74606 41704 74672 41752
rect 74594 41688 74672 41704
rect 74676 41688 74714 41726
rect 73910 41654 73934 41688
rect 73936 41654 74714 41688
rect 73914 41648 73930 41654
rect 73936 41616 74014 41654
rect 73948 41604 74014 41616
rect 73946 40970 74014 41604
rect 74024 41254 74052 41648
rect 74594 41616 74672 41654
rect 74676 41616 74698 41654
rect 74606 40970 74672 41616
rect 74704 41615 74706 41620
rect 74732 41616 74754 41750
rect 75264 41726 75341 41756
rect 75854 41726 75870 41756
rect 75882 41726 75898 41756
rect 75922 41726 75999 41756
rect 76580 41752 76657 41756
rect 75264 41704 75472 41726
rect 75252 41688 75472 41704
rect 75486 41688 76230 41726
rect 76580 41704 76646 41752
rect 76568 41688 76646 41704
rect 76678 41694 76684 41756
rect 76706 41694 76712 41756
rect 76950 41688 76988 41726
rect 77162 41694 77186 41756
rect 77190 41694 77214 41756
rect 77238 41719 77304 41756
rect 77238 41704 77316 41719
rect 77226 41688 77316 41704
rect 74766 41654 75472 41688
rect 75524 41654 76230 41688
rect 76282 41654 76988 41688
rect 77040 41654 77316 41688
rect 75252 41648 75341 41654
rect 75252 41616 75370 41648
rect 74693 41604 74738 41615
rect 73946 40818 73982 40970
rect 73992 40818 73993 40970
rect 74606 40954 74651 40970
rect 74670 40954 74672 40970
rect 74704 40958 74738 41604
rect 75264 40970 75370 41616
rect 74606 40920 74644 40954
rect 74704 40920 74742 40958
rect 75264 40920 75309 40970
rect 75334 40958 75370 40970
rect 75390 40958 75426 41648
rect 75910 41616 75999 41654
rect 76568 41616 76646 41654
rect 77226 41616 77316 41654
rect 75451 41604 75507 41615
rect 75462 40958 75507 41604
rect 75922 40970 75999 41616
rect 76209 41604 76265 41615
rect 75922 40958 75967 40970
rect 76220 40958 76265 41604
rect 76580 40970 76646 41616
rect 76967 41604 77012 41615
rect 75320 40920 75967 40958
rect 75978 40920 76276 40958
rect 76580 40954 76625 40970
rect 76978 40958 77012 41604
rect 77238 40970 77304 41616
rect 76580 40920 76618 40954
rect 76978 40920 77016 40958
rect 77238 40954 77283 40970
rect 77238 40920 77276 40954
rect 74042 40914 74644 40920
rect 74042 40886 74646 40914
rect 74604 40822 74646 40886
rect 74604 40818 74651 40822
rect 74660 40818 74674 40914
rect 74700 40897 75309 40920
rect 74693 40886 75309 40897
rect 75358 40886 75967 40920
rect 76016 40886 76618 40920
rect 76674 40886 77276 40920
rect 74704 40822 74738 40886
rect 74704 40818 74749 40822
rect 75264 40818 75309 40886
rect 75334 40818 75370 40880
rect 75390 40818 75426 40880
rect 75462 40818 75507 40886
rect 75922 40818 75967 40886
rect 76220 40818 76265 40886
rect 76580 40822 76614 40886
rect 76978 40822 77012 40886
rect 77238 40822 77272 40886
rect 76580 40818 76625 40822
rect 76978 40818 77023 40822
rect 77238 40818 77283 40822
rect 77352 40818 77418 41756
rect 77454 41742 77684 41750
rect 77628 41648 77684 41656
rect 77802 41524 78264 41756
rect 78278 41524 78740 41826
rect 85654 41790 85688 43318
rect 93968 41790 94002 43318
rect 115365 42963 115399 45978
rect 118111 45960 118145 45978
rect 115434 45922 118852 45960
rect 115479 43059 115513 43093
rect 116137 43059 116171 43093
rect 116795 43059 116829 43093
rect 117453 43059 117487 43093
rect 118111 43059 118145 45922
rect 118769 43059 118803 43093
rect 115447 43025 118837 43059
rect 97552 41790 97586 42944
rect 81368 41756 99108 41790
rect 85654 41688 85688 41756
rect 85756 41688 85790 41756
rect 86046 41688 86084 41726
rect 86804 41688 86842 41726
rect 87562 41688 87600 41726
rect 88320 41688 88358 41726
rect 89078 41688 89116 41726
rect 89836 41688 89874 41726
rect 90594 41688 90632 41726
rect 91352 41688 91390 41726
rect 92110 41688 92148 41726
rect 92868 41688 92906 41726
rect 93626 41688 93664 41726
rect 93866 41688 93900 41756
rect 93968 41688 94002 41756
rect 85654 41654 86084 41688
rect 86136 41654 86842 41688
rect 86894 41654 87600 41688
rect 87652 41654 88358 41688
rect 88410 41654 89116 41688
rect 89168 41654 89874 41688
rect 89926 41654 90632 41688
rect 90684 41654 91390 41688
rect 91442 41654 92148 41688
rect 92200 41654 92906 41688
rect 92958 41654 93664 41688
rect 93716 41654 94002 41688
rect 96644 41654 96674 41688
rect 77856 41440 78206 41474
rect 77666 41400 77690 41426
rect 77694 41372 77718 41398
rect 77628 41326 77654 41352
rect 73834 40784 77418 40818
rect 72280 38046 72351 40725
rect 72548 38694 72574 38700
rect 72576 38694 72602 38728
rect 72956 38636 73418 39274
rect 73014 38552 73364 38586
rect 73014 38072 73048 38552
rect 73134 38518 73226 38522
rect 73134 38484 73240 38518
rect 73172 38450 73240 38484
rect 73176 38412 73222 38450
rect 73117 38400 73173 38411
rect 73128 38224 73173 38400
rect 73188 38400 73222 38412
rect 73234 38400 73261 38411
rect 73188 38224 73261 38400
rect 73188 38212 73222 38224
rect 73134 38208 73226 38212
rect 73134 38174 73240 38208
rect 73172 38140 73240 38174
rect 73176 38124 73222 38140
rect 73330 38072 73364 38552
rect 73014 38046 73364 38072
rect 73834 38046 73868 40784
rect 73946 38046 73982 40784
rect 73986 38568 73988 38694
rect 73992 38568 73993 40784
rect 74604 40416 74651 40784
rect 74660 40416 74674 40784
rect 74606 39722 74651 40416
rect 74704 39722 74749 40784
rect 74606 39584 74640 39722
rect 74704 39584 74738 39722
rect 73986 38560 74026 38568
rect 74042 38560 74054 38596
rect 73992 38046 73993 38560
rect 74606 38046 74651 39584
rect 74698 38560 74702 38694
rect 74704 38046 74749 39584
rect 75264 38046 75309 40784
rect 75334 40416 75370 40784
rect 75390 40416 75426 40784
rect 75334 38560 75370 39228
rect 75390 38560 75426 39228
rect 75462 38046 75507 40784
rect 75922 38046 75967 40784
rect 76220 38046 76265 40784
rect 76580 39910 76625 40784
rect 76978 39910 77023 40784
rect 76580 39584 76614 39910
rect 76978 39584 77012 39910
rect 77038 39894 77046 39910
rect 77238 39884 77283 40784
rect 77238 39584 77272 39884
rect 76580 38046 76625 39584
rect 76978 38046 77023 39584
rect 77238 38046 77283 39584
rect 77352 38046 77386 40784
rect 77666 40748 77678 41102
rect 77694 40748 77706 41102
rect 77856 40960 77890 41440
rect 78048 41372 78086 41410
rect 78014 41338 78086 41372
rect 77959 41288 78004 41299
rect 78047 41288 78092 41299
rect 77970 41112 78004 41288
rect 78058 41112 78092 41288
rect 78048 41062 78086 41100
rect 78014 41028 78086 41062
rect 78172 40960 78206 41440
rect 77856 40926 78206 40960
rect 78332 41440 78682 41474
rect 78332 40960 78366 41440
rect 78494 41406 78532 41410
rect 78494 41388 78558 41406
rect 78482 41338 78558 41388
rect 78482 41322 78540 41338
rect 78460 41300 78480 41304
rect 78460 41299 78486 41300
rect 78435 41288 78486 41299
rect 78446 41112 78486 41288
rect 78460 41100 78486 41112
rect 78488 41100 78528 41322
rect 78534 41299 78562 41304
rect 78534 41112 78568 41299
rect 78460 41096 78480 41100
rect 78488 41096 78532 41100
rect 78534 41096 78562 41112
rect 78488 41078 78558 41096
rect 78482 41028 78558 41078
rect 78482 41012 78540 41028
rect 78648 40960 78682 41440
rect 78332 40926 78682 40960
rect 77694 40692 77734 40748
rect 84558 38046 84592 41604
rect 85654 39896 85688 41654
rect 85756 41354 85790 41654
rect 85828 41616 85829 41617
rect 93827 41616 93828 41617
rect 85827 41615 85828 41616
rect 93828 41615 93829 41616
rect 86063 41604 86108 41615
rect 86821 41604 86866 41615
rect 87579 41604 87624 41615
rect 88337 41604 88382 41615
rect 89095 41604 89140 41615
rect 89853 41604 89898 41615
rect 90611 41604 90656 41615
rect 91369 41604 91414 41615
rect 92127 41604 92172 41615
rect 92885 41604 92930 41615
rect 93643 41604 93688 41615
rect 86062 41338 86063 41339
rect 86061 41337 86062 41338
rect 86074 41326 86108 41604
rect 86119 41338 86120 41339
rect 86820 41338 86821 41339
rect 86120 41337 86121 41338
rect 86819 41337 86820 41338
rect 86832 41326 86866 41604
rect 86877 41338 86878 41339
rect 87578 41338 87579 41339
rect 86878 41337 86879 41338
rect 87577 41337 87578 41338
rect 87590 41326 87624 41604
rect 87635 41338 87636 41339
rect 88336 41338 88337 41339
rect 87636 41337 87637 41338
rect 88335 41337 88336 41338
rect 88348 41326 88382 41604
rect 88393 41338 88394 41339
rect 89094 41338 89095 41339
rect 88394 41337 88395 41338
rect 89093 41337 89094 41338
rect 89106 41326 89140 41604
rect 89790 41418 89858 41426
rect 89818 41390 89858 41398
rect 89151 41338 89152 41339
rect 89852 41338 89853 41339
rect 89152 41337 89153 41338
rect 89851 41337 89852 41338
rect 89864 41326 89898 41604
rect 89904 41418 89970 41426
rect 89904 41390 89942 41398
rect 89909 41338 89910 41339
rect 90610 41338 90611 41339
rect 89910 41337 89911 41338
rect 90609 41337 90610 41338
rect 90622 41326 90656 41604
rect 91304 41418 91374 41438
rect 91332 41390 91374 41410
rect 90667 41338 90668 41339
rect 91368 41338 91369 41339
rect 90668 41337 90669 41338
rect 91367 41337 91368 41338
rect 91380 41326 91414 41604
rect 91420 41418 91484 41438
rect 91420 41390 91456 41410
rect 91425 41338 91426 41339
rect 92126 41338 92127 41339
rect 91426 41337 91427 41338
rect 92125 41337 92126 41338
rect 92138 41326 92172 41604
rect 92183 41338 92184 41339
rect 92884 41338 92885 41339
rect 92184 41337 92185 41338
rect 92883 41337 92884 41338
rect 92896 41326 92930 41604
rect 92941 41338 92942 41339
rect 93642 41338 93643 41339
rect 92942 41337 92943 41338
rect 93641 41337 93642 41338
rect 93654 41326 93688 41604
rect 93866 41354 93900 41654
rect 93699 41338 93700 41339
rect 93700 41337 93701 41338
rect 93816 41326 93827 41337
rect 85718 41264 85790 41302
rect 85840 41292 93827 41326
rect 86061 41280 86062 41281
rect 86062 41279 86063 41280
rect 85756 40696 85790 41264
rect 86062 40680 86063 40681
rect 86061 40679 86062 40680
rect 86074 40668 86108 41292
rect 86120 41280 86121 41281
rect 86819 41280 86820 41281
rect 86119 41279 86120 41280
rect 86820 41279 86821 41280
rect 86832 40712 86866 41292
rect 86878 41280 86879 41281
rect 87577 41280 87578 41281
rect 86877 41279 86878 41280
rect 87578 41279 87579 41280
rect 86788 40706 86908 40712
rect 86119 40680 86120 40681
rect 86820 40680 86821 40681
rect 86120 40679 86121 40680
rect 86819 40679 86820 40680
rect 86832 40668 86866 40706
rect 86877 40680 86878 40681
rect 87578 40680 87579 40681
rect 86878 40679 86879 40680
rect 87577 40679 87578 40680
rect 87590 40668 87624 41292
rect 87636 41280 87637 41281
rect 88335 41280 88336 41281
rect 87635 41279 87636 41280
rect 88336 41279 88337 41280
rect 87635 40680 87636 40681
rect 88336 40680 88337 40681
rect 87636 40679 87637 40680
rect 88335 40679 88336 40680
rect 88348 40668 88382 41292
rect 88394 41280 88395 41281
rect 89093 41280 89094 41281
rect 88393 41279 88394 41280
rect 89094 41279 89095 41280
rect 88393 40680 88394 40681
rect 89094 40680 89095 40681
rect 88394 40679 88395 40680
rect 89093 40679 89094 40680
rect 89106 40668 89140 41292
rect 89152 41280 89153 41281
rect 89851 41280 89852 41281
rect 89151 41279 89152 41280
rect 89852 41279 89853 41280
rect 89151 40680 89152 40681
rect 89852 40680 89853 40681
rect 89152 40679 89153 40680
rect 89851 40679 89852 40680
rect 89864 40668 89898 41292
rect 89910 41280 89911 41281
rect 90609 41280 90610 41281
rect 89909 41279 89910 41280
rect 90610 41279 90611 41280
rect 89909 40680 89910 40681
rect 90610 40680 90611 40681
rect 89910 40679 89911 40680
rect 90609 40679 90610 40680
rect 90622 40668 90656 41292
rect 90668 41280 90669 41281
rect 91367 41280 91368 41281
rect 90667 41279 90668 41280
rect 91368 41279 91369 41280
rect 90667 40680 90668 40681
rect 91368 40680 91369 40681
rect 90668 40679 90669 40680
rect 91367 40679 91368 40680
rect 91380 40668 91414 41292
rect 91426 41280 91427 41281
rect 92125 41280 92126 41281
rect 91425 41279 91426 41280
rect 92126 41279 92127 41280
rect 91425 40680 91426 40681
rect 92126 40680 92127 40681
rect 91426 40679 91427 40680
rect 92125 40679 92126 40680
rect 92138 40668 92172 41292
rect 92184 41280 92185 41281
rect 92883 41280 92884 41281
rect 92183 41279 92184 41280
rect 92884 41279 92885 41280
rect 92183 40680 92184 40681
rect 92884 40680 92885 40681
rect 92184 40679 92185 40680
rect 92883 40679 92884 40680
rect 92896 40668 92930 41292
rect 92942 41280 92943 41281
rect 93641 41280 93642 41281
rect 92941 41279 92942 41280
rect 93642 41279 93643 41280
rect 92941 40680 92942 40681
rect 93642 40680 93643 40681
rect 92942 40679 92943 40680
rect 93641 40679 93642 40680
rect 93654 40668 93688 41292
rect 93700 41280 93701 41281
rect 93699 41279 93700 41280
rect 93828 41264 93900 41302
rect 93866 40696 93900 41264
rect 93699 40680 93700 40681
rect 93700 40679 93701 40680
rect 93816 40668 93827 40679
rect 85718 40606 85790 40644
rect 85840 40634 93827 40668
rect 86061 40622 86062 40623
rect 86062 40621 86063 40622
rect 85756 40038 85790 40606
rect 86062 40022 86063 40023
rect 86061 40021 86062 40022
rect 86074 40010 86108 40634
rect 86120 40622 86121 40623
rect 86819 40622 86820 40623
rect 86119 40621 86120 40622
rect 86820 40621 86821 40622
rect 86119 40022 86120 40023
rect 86820 40022 86821 40023
rect 86120 40021 86121 40022
rect 86819 40021 86820 40022
rect 86832 40010 86866 40634
rect 86878 40622 86879 40623
rect 87577 40622 87578 40623
rect 86877 40621 86878 40622
rect 87578 40621 87579 40622
rect 86877 40022 86878 40023
rect 87578 40022 87579 40023
rect 86878 40021 86879 40022
rect 87577 40021 87578 40022
rect 87590 40010 87624 40634
rect 87636 40622 87637 40623
rect 88335 40622 88336 40623
rect 87635 40621 87636 40622
rect 88336 40621 88337 40622
rect 87635 40022 87636 40023
rect 88336 40022 88337 40023
rect 87636 40021 87637 40022
rect 88335 40021 88336 40022
rect 88348 40010 88382 40634
rect 88394 40622 88395 40623
rect 89093 40622 89094 40623
rect 88393 40621 88394 40622
rect 89094 40621 89095 40622
rect 88393 40022 88394 40023
rect 89094 40022 89095 40023
rect 88394 40021 88395 40022
rect 89093 40021 89094 40022
rect 89106 40010 89140 40634
rect 89152 40622 89153 40623
rect 89851 40622 89852 40623
rect 89151 40621 89152 40622
rect 89852 40621 89853 40622
rect 89756 40042 89766 40108
rect 89784 40070 89794 40108
rect 89151 40022 89152 40023
rect 89852 40022 89853 40023
rect 89152 40021 89153 40022
rect 89851 40021 89852 40022
rect 89864 40010 89898 40634
rect 89910 40622 89911 40623
rect 90609 40622 90610 40623
rect 89909 40621 89910 40622
rect 90610 40621 90611 40622
rect 89909 40022 89910 40023
rect 90610 40022 90611 40023
rect 89910 40021 89911 40022
rect 90609 40021 90610 40022
rect 90622 40010 90656 40634
rect 90668 40622 90669 40623
rect 91367 40622 91368 40623
rect 90667 40621 90668 40622
rect 91368 40621 91369 40622
rect 90667 40022 90668 40023
rect 90668 40021 90669 40022
rect 91332 40020 91374 40044
rect 91304 40010 91374 40016
rect 91380 40010 91414 40634
rect 91426 40622 91427 40623
rect 92125 40622 92126 40623
rect 91425 40621 91426 40622
rect 92126 40621 92127 40622
rect 91420 40020 91456 40044
rect 92126 40022 92127 40023
rect 92125 40021 92126 40022
rect 91420 40010 91484 40016
rect 92138 40010 92172 40634
rect 92184 40622 92185 40623
rect 92883 40622 92884 40623
rect 92183 40621 92184 40622
rect 92884 40621 92885 40622
rect 92183 40022 92184 40023
rect 92884 40022 92885 40023
rect 92184 40021 92185 40022
rect 92883 40021 92884 40022
rect 92896 40010 92930 40634
rect 92942 40622 92943 40623
rect 93641 40622 93642 40623
rect 92941 40621 92942 40622
rect 93642 40621 93643 40622
rect 92941 40022 92942 40023
rect 93642 40022 93643 40023
rect 92942 40021 92943 40022
rect 93641 40021 93642 40022
rect 93654 40010 93688 40634
rect 93700 40622 93701 40623
rect 93699 40621 93700 40622
rect 93828 40606 93900 40644
rect 93866 40038 93900 40606
rect 93699 40022 93700 40023
rect 93700 40021 93701 40022
rect 93816 40010 93827 40021
rect 85840 39976 93827 40010
rect 86074 39896 86108 39976
rect 86832 39896 86866 39976
rect 87590 39896 87624 39976
rect 88348 39896 88382 39976
rect 89106 39896 89140 39976
rect 89864 39896 89898 39976
rect 90622 39896 90656 39976
rect 91380 39896 91414 39976
rect 92138 39896 92172 39976
rect 92896 39896 92930 39976
rect 93654 39896 93688 39976
rect 93968 39896 94002 41654
rect 96678 41620 96708 41722
rect 97552 41688 97586 41756
rect 97630 41708 97648 41722
rect 97602 41688 97648 41694
rect 97654 41688 97688 41756
rect 98174 41722 98212 41726
rect 98932 41722 98970 41726
rect 97694 41708 98214 41722
rect 98224 41708 98972 41722
rect 98174 41694 98212 41708
rect 98932 41694 98970 41708
rect 97694 41688 98212 41694
rect 97552 41654 98212 41688
rect 98252 41680 98970 41694
rect 98264 41654 98970 41680
rect 96704 40154 96720 40672
rect 96742 40192 96758 40634
rect 85654 39862 94002 39896
rect 89106 38379 89140 39862
rect 89740 39528 89766 39558
rect 89768 39556 89794 39558
rect 89830 39556 89854 39558
rect 89858 39528 89882 39558
rect 97552 39522 97586 41654
rect 97654 41638 97688 41654
rect 97726 41616 98190 41622
rect 98248 41616 98948 41622
rect 99074 41610 99108 41756
rect 97616 41548 97688 41586
rect 97738 41576 99108 41610
rect 98189 41564 98190 41565
rect 98190 41563 98191 41564
rect 97654 40980 97688 41548
rect 98190 40964 98191 40965
rect 98189 40963 98190 40964
rect 98202 40952 98236 41576
rect 98248 41564 98249 41565
rect 98947 41564 98948 41565
rect 98247 41563 98248 41564
rect 98948 41563 98949 41564
rect 98247 40964 98248 40965
rect 98948 40964 98949 40965
rect 98248 40963 98249 40964
rect 98947 40963 98948 40964
rect 98960 40952 98994 41576
rect 99074 40952 99108 41576
rect 97616 40890 97688 40928
rect 97738 40918 99108 40952
rect 98189 40906 98190 40907
rect 98190 40905 98191 40906
rect 97654 40322 97688 40890
rect 98190 40306 98191 40307
rect 98189 40305 98190 40306
rect 98202 40294 98236 40918
rect 98248 40906 98249 40907
rect 98947 40906 98948 40907
rect 98247 40905 98248 40906
rect 98948 40905 98949 40906
rect 98247 40306 98248 40307
rect 98948 40306 98949 40307
rect 98248 40305 98249 40306
rect 98947 40305 98948 40306
rect 98960 40294 98994 40918
rect 99074 40294 99108 40918
rect 97616 40232 97688 40270
rect 97738 40260 99108 40294
rect 98189 40248 98190 40249
rect 98190 40247 98191 40248
rect 97654 39664 97688 40232
rect 98190 39648 98191 39649
rect 98189 39647 98190 39648
rect 98202 39636 98236 40260
rect 98248 40248 98249 40249
rect 98947 40248 98948 40249
rect 98247 40247 98248 40248
rect 98948 40247 98949 40248
rect 98247 39648 98248 39649
rect 98948 39648 98949 39649
rect 98248 39647 98249 39648
rect 98947 39647 98948 39648
rect 98960 39636 98994 40260
rect 99074 39636 99108 40260
rect 97738 39618 99108 39636
rect 115351 41461 115399 42963
rect 115479 42973 115513 43025
rect 116137 43004 116171 43025
rect 116795 43004 116829 43025
rect 117453 43004 117487 43025
rect 118111 43004 118145 43025
rect 118769 43004 118803 43025
rect 116095 42973 116171 43004
rect 116753 42973 116829 43004
rect 117411 42973 117487 43004
rect 118069 42973 118145 43004
rect 115479 42876 115525 42973
rect 116095 42957 116183 42973
rect 116753 42957 116841 42973
rect 117411 42957 117499 42973
rect 118069 42957 118157 42973
rect 118727 42957 118803 43004
rect 118883 42963 118917 45978
rect 120436 46006 120470 47848
rect 120538 47786 120584 47938
rect 121136 47894 121162 49014
rect 121164 47894 121190 48986
rect 121208 47938 121274 49550
rect 121866 47938 121932 49550
rect 121208 47926 121242 47938
rect 121866 47926 121900 47938
rect 121196 47888 121246 47926
rect 121300 47894 121318 47910
rect 121854 47888 121904 47926
rect 122456 47894 122472 48996
rect 122484 47894 122500 48968
rect 122524 47938 122590 49550
rect 123182 47938 123248 49550
rect 123280 48192 123286 49594
rect 123308 48164 123314 49594
rect 123829 49550 123860 49561
rect 123872 49550 123906 49702
rect 122524 47926 122558 47938
rect 123182 47926 123216 47938
rect 122512 47888 122562 47926
rect 123170 47888 123220 47926
rect 123764 47894 123788 48998
rect 123792 47894 123816 48970
rect 123840 47938 123906 49550
rect 123954 49640 123972 49702
rect 123986 49640 124020 49942
rect 123840 47926 123874 47938
rect 123828 47888 123878 47926
rect 120644 47854 121246 47888
rect 121302 47854 121904 47888
rect 121960 47854 122562 47888
rect 122618 47854 123220 47888
rect 123276 47854 123878 47888
rect 121196 47838 121242 47854
rect 121854 47838 121900 47854
rect 122512 47838 122558 47854
rect 123170 47838 123216 47854
rect 123828 47838 123874 47854
rect 123954 47848 124020 49640
rect 124574 48576 124694 48596
rect 124880 48578 125120 49130
rect 124880 48576 125170 48578
rect 124568 48548 124722 48568
rect 124880 48550 125120 48576
rect 124880 48548 125198 48550
rect 124880 48492 125120 48548
rect 121208 47786 121242 47838
rect 120538 47752 123886 47786
rect 121208 46006 121242 47752
rect 123176 46006 123198 46196
rect 123954 46006 123988 47848
rect 131942 46520 131944 46570
rect 131970 46520 131972 46598
rect 131390 46280 132028 46520
rect 137156 46476 137158 46554
rect 137184 46476 137186 46526
rect 137100 46236 137738 46476
rect 120436 45978 123988 46006
rect 120130 45536 120132 45584
rect 120102 45508 120132 45528
rect 120436 42968 120470 45978
rect 121208 45950 121242 45978
rect 123176 45950 123198 45978
rect 120508 45922 123926 45950
rect 120550 43064 120584 43098
rect 121208 43064 121242 45922
rect 123176 45528 123198 45922
rect 121900 43266 121906 44340
rect 121900 43098 121932 43266
rect 121866 43064 121932 43098
rect 121956 43064 121960 43294
rect 122524 43064 122558 43098
rect 123118 43064 123144 43258
rect 123176 43230 123200 44340
rect 123146 43098 123200 43230
rect 123146 43064 123216 43098
rect 123840 43064 123874 43098
rect 120518 43030 123908 43064
rect 115527 42923 116183 42957
rect 116185 42923 116841 42957
rect 116843 42923 117499 42957
rect 117501 42923 118157 42957
rect 118159 42923 118803 42957
rect 116103 42917 116107 42923
rect 116131 42889 116135 42923
rect 116137 42876 116183 42923
rect 116795 42876 116841 42923
rect 117419 42917 117423 42923
rect 117447 42889 117451 42923
rect 117453 42876 117499 42923
rect 118111 42876 118157 42923
rect 118735 42917 118739 42923
rect 118763 42889 118767 42923
rect 115479 42864 115513 42876
rect 116112 42864 116125 42875
rect 116137 42864 116171 42876
rect 116770 42864 116783 42875
rect 116795 42864 116829 42876
rect 117428 42864 117441 42875
rect 117453 42864 117487 42876
rect 118086 42864 118099 42875
rect 118111 42864 118145 42876
rect 118744 42864 118757 42875
rect 118769 42864 118803 42923
rect 115465 41560 115513 42864
rect 116123 41560 116171 42864
rect 116781 41560 116829 42864
rect 97722 39602 99232 39618
rect 98202 39584 98236 39602
rect 98960 39584 98994 39602
rect 99074 39584 99108 39602
rect 97688 39568 99198 39584
rect 98202 39522 98236 39568
rect 98960 39522 98994 39568
rect 99074 39522 99108 39568
rect 89346 39446 89668 39518
rect 97552 39488 101528 39522
rect 89148 38984 89786 39446
rect 89836 39358 90384 39392
rect 89836 39076 89870 39358
rect 90011 39278 90209 39289
rect 89900 39234 90010 39272
rect 90022 39244 90209 39278
rect 90210 39234 90320 39272
rect 89938 39200 90010 39234
rect 90011 39190 90209 39201
rect 90248 39200 90320 39234
rect 90022 39156 90209 39190
rect 90350 39076 90384 39358
rect 89836 39042 90384 39076
rect 91346 39036 91364 39236
rect 91374 39008 91392 39264
rect 85623 38046 94061 38379
rect 72280 38012 72369 38046
rect 72418 38023 99006 38046
rect 99074 38023 99108 39488
rect 72418 38012 99108 38023
rect 72280 36904 72351 38012
rect 72430 37044 72464 38012
rect 73188 37982 73222 38012
rect 73010 37944 73748 37982
rect 73834 37944 73868 38012
rect 73946 37982 73982 38012
rect 73918 37944 73982 37982
rect 72476 37910 73222 37944
rect 73250 37910 73982 37944
rect 73188 37044 73222 37910
rect 72430 37006 72504 37044
rect 73160 37006 73222 37044
rect 73834 37006 73868 37910
rect 73946 37044 73982 37910
rect 73918 37040 73982 37044
rect 73992 37944 73993 38012
rect 74606 38008 74651 38012
rect 74704 38008 74749 38012
rect 74606 37982 74640 38008
rect 74704 37982 74738 38008
rect 75264 37982 75309 38012
rect 75462 37982 75507 38012
rect 75922 37982 75967 38012
rect 76220 37982 76265 38012
rect 74606 37944 74644 37982
rect 74676 37944 74738 37982
rect 75260 37944 76265 37982
rect 76580 38008 76625 38012
rect 76978 38008 77023 38012
rect 77238 38008 77283 38012
rect 76580 37982 76614 38008
rect 76978 37982 77012 38008
rect 76580 37944 76618 37982
rect 76950 37944 77012 37982
rect 77238 37982 77272 38008
rect 77238 37944 77276 37982
rect 77352 37944 77386 38012
rect 77736 37982 77770 38012
rect 78494 37982 78528 38012
rect 79252 37982 79286 38012
rect 80010 37982 80044 38012
rect 80768 37982 80802 38012
rect 81526 37982 81560 38012
rect 82284 37982 82318 38012
rect 83042 37982 83076 38012
rect 83800 37982 83834 38012
rect 83844 37982 83868 38008
rect 84558 37982 84592 38012
rect 85316 37982 85350 38012
rect 85623 37982 94061 38012
rect 94412 37982 94446 38012
rect 95170 37982 95204 38012
rect 95928 37982 95962 38012
rect 96686 37982 96720 38012
rect 97444 37982 97478 38012
rect 99074 38005 99108 38012
rect 77708 37944 77770 37982
rect 78466 37944 78528 37982
rect 79224 37944 79286 37982
rect 79982 37944 80044 37982
rect 80740 37944 80802 37982
rect 81498 37944 81560 37982
rect 82256 37944 82318 37982
rect 83014 37944 83076 37982
rect 83772 37944 94061 37982
rect 94384 37944 94446 37982
rect 95142 37944 95204 37982
rect 95900 37944 95962 37982
rect 96658 37944 96720 37982
rect 97416 37978 97478 37982
rect 97416 37950 97484 37978
rect 97410 37944 97484 37950
rect 97493 37944 99144 38005
rect 73992 37910 74738 37944
rect 74750 37910 75507 37944
rect 75524 37910 76265 37944
rect 76282 37910 77012 37944
rect 77024 37910 77770 37944
rect 77782 37910 78528 37944
rect 78540 37910 79286 37944
rect 79298 37910 80044 37944
rect 80056 37910 80802 37944
rect 80814 37910 81560 37944
rect 81572 37910 82318 37944
rect 82330 37910 83076 37944
rect 83088 37910 83834 37944
rect 73918 37012 73988 37040
rect 73912 37006 73988 37012
rect 72430 36938 72470 37006
rect 72480 36972 73222 37006
rect 73234 36972 73988 37006
rect 72480 36966 72498 36972
rect 72430 36904 72464 36938
rect 73188 36904 73222 36972
rect 73834 36904 73868 36972
rect 73912 36966 73930 36972
rect 73940 36938 73988 36972
rect 73992 37006 73993 37910
rect 74606 37372 74640 37910
rect 74604 37012 74646 37372
rect 74660 37012 74674 37372
rect 74704 37044 74738 37910
rect 75264 37044 75309 37910
rect 75334 37044 75370 37372
rect 75390 37044 75426 37372
rect 75462 37044 75507 37910
rect 75922 37044 75967 37910
rect 76220 37044 76265 37910
rect 73996 37006 74016 37012
rect 74606 37006 74644 37012
rect 74676 37006 74738 37044
rect 75260 37006 76265 37044
rect 76580 37044 76614 37910
rect 76978 37044 77012 37910
rect 76580 37006 76618 37044
rect 76950 37006 77012 37044
rect 77238 37044 77272 37910
rect 77238 37006 77276 37044
rect 77352 37006 77386 37910
rect 77736 37906 77770 37910
rect 78494 37906 78528 37910
rect 79252 37906 79286 37910
rect 80010 37906 80044 37910
rect 80768 37906 80802 37910
rect 77524 37876 81202 37906
rect 77736 37044 77770 37876
rect 78494 37044 78528 37876
rect 79252 37044 79286 37876
rect 80010 37044 80044 37876
rect 80768 37044 80802 37876
rect 81526 37044 81560 37910
rect 82284 37044 82318 37910
rect 83042 37044 83076 37910
rect 83800 37044 83834 37910
rect 83844 37910 84592 37944
rect 84620 37910 85350 37944
rect 85378 37910 94446 37944
rect 94458 37910 95204 37944
rect 95216 37910 95962 37944
rect 95974 37910 96720 37944
rect 96732 37910 97484 37944
rect 97490 37910 99144 37944
rect 83844 37044 83868 37910
rect 84558 37044 84592 37910
rect 85316 37044 85350 37910
rect 85623 37044 94061 37910
rect 94412 37044 94446 37910
rect 95170 37044 95204 37910
rect 95928 37044 95962 37910
rect 96686 37044 96720 37910
rect 97410 37904 97428 37910
rect 97438 37876 97484 37910
rect 97444 37044 97478 37876
rect 77500 37006 81260 37044
rect 81498 37040 81560 37044
rect 81498 37012 81566 37040
rect 81492 37006 81566 37012
rect 81576 37006 81594 37012
rect 82256 37006 82318 37044
rect 83014 37040 83076 37044
rect 83014 37012 83082 37040
rect 83008 37006 83082 37012
rect 83092 37006 83110 37012
rect 83772 37006 94061 37044
rect 94384 37006 94446 37044
rect 95142 37006 95204 37044
rect 95900 37006 95962 37044
rect 96658 37006 96720 37044
rect 97416 37006 97478 37044
rect 97493 37006 99144 37910
rect 73992 36972 74738 37006
rect 74750 36972 75507 37006
rect 75524 36972 76265 37006
rect 76282 36972 77012 37006
rect 77024 36972 77770 37006
rect 77798 36972 78534 37006
rect 73946 36904 73982 36938
rect 73992 36904 73993 36972
rect 73996 36966 74016 36972
rect 74606 36966 74640 36972
rect 74604 36904 74646 36966
rect 74660 36904 74674 36966
rect 74704 36904 74738 36972
rect 75264 36904 75309 36972
rect 75334 36904 75370 36966
rect 75390 36904 75426 36966
rect 75462 36904 75507 36972
rect 75922 36904 75967 36972
rect 76220 36904 76265 36972
rect 76580 36904 76614 36972
rect 76978 36904 77012 36972
rect 77238 36904 77272 36972
rect 77352 36904 77386 36972
rect 77736 36904 77770 36972
rect 78460 36966 78478 36972
rect 78488 36938 78534 36972
rect 78544 36972 79286 37006
rect 79314 36972 80050 37006
rect 78544 36966 78562 36972
rect 78494 36904 78528 36938
rect 79252 36904 79286 36972
rect 79976 36966 79994 36972
rect 80004 36938 80050 36972
rect 80060 36972 80802 37006
rect 80830 36972 81566 37006
rect 81572 36972 82318 37006
rect 82330 36972 83082 37006
rect 83088 36972 83834 37006
rect 80060 36966 80078 36972
rect 80010 36904 80044 36938
rect 80768 36904 80802 36972
rect 81492 36966 81510 36972
rect 81520 36938 81566 36972
rect 81576 36966 81594 36972
rect 81526 36904 81560 36938
rect 82284 36904 82318 36972
rect 83008 36966 83026 36972
rect 83036 36938 83082 36972
rect 83092 36966 83110 36972
rect 83042 36904 83076 36938
rect 83800 36904 83834 36972
rect 83844 36972 84598 37006
rect 83844 36904 83868 36972
rect 84524 36966 84542 36972
rect 84552 36938 84598 36972
rect 84608 36972 85350 37006
rect 85378 36972 94446 37006
rect 94458 36972 95204 37006
rect 95216 36972 95962 37006
rect 95974 36972 96720 37006
rect 96732 36972 97478 37006
rect 97490 36972 99144 37006
rect 84608 36966 84626 36972
rect 84558 36904 84592 36938
rect 85316 36904 85350 36972
rect 85623 36904 94061 36972
rect 94412 36904 94446 36972
rect 95170 36904 95204 36972
rect 95928 36904 95962 36972
rect 96686 36904 96720 36972
rect 97444 36904 97478 36972
rect 97493 36904 99144 36972
rect 72280 36870 72369 36904
rect 72412 36870 99144 36904
rect 51056 36822 51676 36834
rect 51056 36820 51708 36822
rect 51056 36787 51766 36820
rect 51056 36753 59239 36787
rect 51056 36717 51676 36753
rect 51726 36620 51766 36753
rect 51774 36626 51794 36746
rect 51828 36719 51862 36722
rect 52156 36719 52190 36722
rect 51726 36588 51760 36620
rect 52258 36588 52292 36753
rect 44324 36298 44788 36310
rect 44324 36264 44788 36276
rect 68763 35995 68797 36834
rect 72280 36626 72351 36870
rect 72212 36384 72250 36570
rect 72268 36384 72351 36626
rect 68877 36091 68911 36125
rect 69535 36091 69569 36125
rect 70193 36091 70227 36125
rect 70851 36091 70885 36125
rect 71509 36091 71543 36125
rect 72167 36091 72201 36125
rect 68845 36057 72235 36091
rect 46030 35604 46960 35618
rect 45494 34364 45518 34418
rect 45522 34364 45574 34390
rect 45494 34254 45518 34318
rect 45522 34282 45574 34318
rect 45642 33700 47436 35446
rect 41048 33666 47436 33700
rect 45642 32858 47436 33666
rect 50914 33756 55150 35446
rect 68749 34493 68797 35995
rect 68877 36005 68911 36057
rect 69535 36036 69569 36057
rect 69493 36005 69569 36036
rect 69592 36036 69603 36054
rect 70193 36036 70227 36057
rect 70851 36036 70885 36057
rect 71509 36036 71543 36057
rect 72167 36036 72201 36057
rect 68877 35908 68923 36005
rect 69493 35989 69581 36005
rect 69592 35989 72201 36036
rect 72280 35995 72351 36384
rect 68925 35955 69581 35989
rect 69583 35955 70239 35989
rect 70241 35955 70897 35989
rect 70899 35955 71555 35989
rect 71557 35955 72201 35989
rect 69501 35949 69505 35955
rect 69529 35921 69533 35955
rect 69535 35908 69581 35955
rect 68877 35896 68911 35908
rect 69510 35896 69523 35907
rect 69535 35896 69569 35908
rect 68863 34592 68911 35896
rect 69521 34592 69569 35896
rect 50914 33544 55268 33756
rect 45678 31375 45712 32858
rect 50914 32484 55150 33544
rect 54932 32358 54938 32436
rect 54960 32358 54966 32464
rect 54912 32104 55150 32358
rect 54932 32086 54938 32104
rect 54960 32086 54966 32104
rect 55166 32086 55404 32104
rect 52182 31704 52188 31904
rect 54532 31664 55150 32086
rect 68749 31840 68783 34493
rect 68863 34431 68897 34592
rect 69521 34580 69555 34592
rect 69558 34580 69569 34592
rect 69592 34580 69603 35955
rect 70193 35908 70239 35955
rect 70817 35949 70821 35955
rect 70845 35921 70849 35955
rect 70851 35908 70897 35955
rect 71509 35908 71555 35955
rect 72133 35949 72137 35955
rect 72161 35921 72165 35955
rect 70168 35896 70181 35907
rect 70193 35896 70238 35908
rect 70826 35896 70839 35907
rect 70851 35896 70896 35908
rect 71484 35896 71497 35907
rect 71509 35896 71554 35908
rect 72142 35896 72155 35907
rect 72167 35896 72201 35955
rect 70179 34592 70238 35896
rect 70179 34580 70213 34592
rect 70760 34580 70762 35314
rect 70788 34580 70790 35314
rect 70837 34592 70896 35896
rect 71495 34592 71554 35896
rect 70837 34580 70871 34592
rect 71495 34580 71529 34592
rect 72082 34580 72084 35606
rect 72110 34580 72112 35578
rect 72153 34592 72201 35896
rect 72153 34580 72187 34592
rect 68899 34465 68903 34567
rect 68927 34533 68931 34539
rect 69507 34533 72187 34580
rect 68923 34499 68931 34533
rect 68939 34499 69555 34533
rect 69581 34499 69589 34533
rect 69597 34499 70213 34533
rect 68927 34493 68931 34499
rect 69509 34483 69555 34499
rect 70167 34483 70213 34499
rect 69521 34431 69555 34483
rect 70179 34431 70213 34483
rect 70215 34465 70219 34533
rect 70243 34493 70247 34533
rect 70255 34499 70871 34533
rect 70913 34499 71529 34533
rect 70760 34486 70762 34493
rect 70788 34458 70790 34493
rect 70825 34483 70871 34499
rect 71483 34483 71529 34499
rect 70837 34431 70871 34483
rect 71495 34431 71529 34483
rect 71531 34465 71535 34533
rect 71559 34493 71563 34533
rect 71571 34499 72187 34533
rect 72082 34486 72084 34493
rect 72110 34458 72112 34493
rect 72141 34483 72187 34499
rect 72153 34431 72187 34483
rect 68851 34397 72199 34431
rect 72234 34226 72238 34638
rect 72267 34361 72351 35995
rect 72267 33160 72350 34361
rect 72430 34174 72464 36870
rect 73834 36096 73868 36870
rect 73946 36096 73982 36870
rect 73992 36096 73993 36870
rect 74604 36308 74646 36870
rect 74604 36194 74651 36308
rect 74660 36250 74674 36870
rect 74704 36308 74738 36870
rect 74606 36096 74651 36194
rect 74704 36096 74749 36308
rect 75264 36096 75309 36870
rect 75334 36096 75370 36870
rect 75390 36096 75426 36870
rect 75462 36096 75507 36870
rect 75922 36096 75967 36870
rect 76220 36096 76265 36870
rect 76580 36308 76614 36870
rect 76978 36308 77012 36870
rect 77238 36308 77272 36870
rect 76580 36096 76625 36308
rect 76978 36096 77023 36308
rect 77238 36096 77283 36308
rect 77352 36096 77386 36870
rect 80010 36127 80044 36870
rect 73820 36062 77386 36096
rect 73820 35446 73868 36062
rect 73946 36032 73982 36062
rect 73992 36032 73993 36062
rect 74606 36032 74651 36062
rect 74704 36032 74749 36062
rect 75264 36032 75309 36062
rect 75320 36032 75370 36062
rect 75390 36032 75426 36062
rect 75462 36032 75507 36062
rect 75922 36032 75967 36062
rect 76220 36032 76265 36062
rect 76580 36032 76625 36062
rect 76978 36032 77023 36062
rect 73946 35994 74602 36032
rect 73923 35910 73934 35921
rect 73946 35910 73993 35994
rect 73996 35960 74602 35994
rect 74606 35994 75260 36032
rect 74606 35921 74651 35994
rect 74654 35960 75260 35994
rect 75264 35994 75918 36032
rect 74692 35922 74750 35960
rect 75264 35950 75309 35994
rect 75312 35960 75918 35994
rect 75922 35994 76576 36032
rect 75320 35950 75370 35954
rect 74581 35910 74651 35921
rect 73934 35446 73993 35910
rect 74592 35446 74651 35910
rect 74704 35446 74749 35922
rect 75246 35921 75370 35950
rect 75239 35910 75370 35921
rect 75246 35808 75370 35910
rect 74960 35446 75370 35808
rect 75376 35446 75426 35954
rect 75450 35922 75508 35960
rect 75462 35446 75507 35922
rect 75922 35921 75967 35994
rect 75970 35960 76576 35994
rect 76580 35994 77234 36032
rect 76208 35922 76266 35960
rect 76580 35942 76625 35994
rect 76628 35960 77234 35994
rect 75897 35910 75967 35921
rect 75908 35446 75967 35910
rect 76220 35446 76265 35922
rect 76562 35921 76636 35942
rect 76966 35922 77024 35960
rect 76555 35910 76636 35921
rect 76562 35842 76636 35910
rect 76432 35446 76754 35842
rect 76978 35446 77023 35922
rect 77238 35921 77283 36062
rect 77213 35910 77283 35921
rect 77224 35446 77283 35910
rect 77338 35446 77386 36062
rect 77469 35446 81093 36127
rect 82542 35446 82570 36130
rect 83810 36096 83834 36870
rect 83844 36096 83868 36870
rect 85623 36096 94061 36870
rect 73042 35376 82570 35446
rect 82576 36062 94061 36096
rect 72386 34152 72506 34174
rect 72386 34026 72798 34152
rect 72392 33622 72798 34026
rect 72430 33312 72464 33622
rect 73042 33160 82550 35376
rect 82576 33160 82610 36062
rect 83810 36032 83834 36062
rect 83844 36032 83868 36062
rect 85316 36032 85350 36062
rect 85623 36032 94061 36062
rect 83042 36010 83080 36032
rect 83030 35994 83088 36010
rect 83320 35994 83358 36032
rect 83800 36010 83838 36032
rect 83844 36010 84016 36032
rect 83788 35994 84016 36010
rect 84030 35994 84674 36032
rect 84688 35994 94061 36032
rect 82752 35960 83358 35994
rect 83410 35960 84016 35994
rect 84068 35960 84674 35994
rect 84726 35960 85356 35994
rect 83030 35922 83088 35960
rect 83788 35922 83868 35960
rect 84546 35922 84604 35960
rect 85282 35954 85356 35960
rect 85372 35960 94061 35994
rect 85372 35954 85384 35960
rect 82679 35910 82724 35921
rect 82690 33300 82724 35910
rect 83042 33312 83076 35922
rect 83337 35910 83382 35921
rect 83348 33300 83382 35910
rect 83800 33312 83834 35922
rect 83844 34810 83868 35922
rect 83995 35910 84051 35921
rect 84006 34810 84051 35910
rect 83900 33990 83922 34294
rect 83956 33990 83978 34294
rect 84006 33300 84040 34810
rect 84558 34786 84603 35922
rect 84692 35921 84704 35922
rect 84653 35910 84709 35921
rect 84624 34804 84654 35328
rect 84664 34786 84709 35910
rect 84720 35328 84732 35950
rect 85304 35926 85356 35954
rect 85304 35922 85310 35926
rect 85316 35910 85350 35926
rect 84558 33312 84592 34786
rect 84664 34224 84698 34786
rect 84630 33414 84642 34224
rect 84658 33358 84704 34224
rect 84664 33300 84704 33358
rect 84720 33929 84732 34224
rect 85316 33929 85356 35910
rect 85362 33929 85367 35921
rect 85623 34755 94061 35960
rect 85980 34226 86014 34755
rect 85946 33929 85972 34226
rect 85974 33929 86020 34226
rect 86034 33929 86048 34226
rect 86094 33929 86128 34755
rect 91264 33929 91274 34124
rect 91292 33929 91302 34096
rect 82678 33262 82736 33300
rect 83014 33262 83052 33300
rect 83336 33262 83394 33300
rect 83772 33262 83810 33300
rect 83994 33262 84052 33300
rect 84530 33262 84568 33300
rect 84652 33268 84710 33300
rect 84720 33268 93169 33929
rect 95928 33312 95962 36870
rect 97493 34668 99144 36870
rect 115351 34789 115385 41461
rect 115465 41399 115499 41560
rect 116123 41548 116157 41560
rect 116781 41548 116815 41560
rect 115501 41433 115505 41535
rect 115529 41501 115533 41507
rect 116109 41501 116157 41548
rect 116767 41501 116815 41548
rect 115525 41467 115533 41501
rect 115541 41467 116157 41501
rect 116183 41467 116191 41501
rect 116199 41467 116815 41501
rect 115529 41461 115533 41467
rect 116111 41451 116157 41467
rect 116769 41451 116815 41467
rect 116123 41399 116157 41451
rect 116781 41399 116815 41451
rect 116817 41433 116821 41535
rect 117362 41507 117364 42604
rect 117390 41507 117392 42576
rect 117439 41560 117487 42864
rect 118097 41560 118145 42864
rect 117439 41548 117473 41560
rect 118097 41548 118131 41560
rect 116845 41501 116849 41507
rect 117425 41501 117473 41548
rect 118083 41501 118131 41548
rect 116841 41467 116849 41501
rect 116857 41467 117473 41501
rect 117499 41467 117507 41501
rect 117515 41467 118131 41501
rect 116845 41461 116849 41467
rect 117362 41454 117364 41461
rect 117390 41426 117392 41461
rect 117427 41451 117473 41467
rect 118085 41451 118131 41467
rect 117439 41399 117473 41451
rect 118097 41399 118131 41451
rect 118133 41433 118137 41535
rect 118684 41507 118686 42574
rect 118712 41507 118714 42546
rect 118755 41560 118803 42864
rect 118755 41548 118789 41560
rect 118161 41501 118165 41507
rect 118741 41501 118789 41548
rect 118157 41467 118165 41501
rect 118173 41467 118789 41501
rect 118161 41461 118165 41467
rect 118684 41454 118686 41461
rect 118712 41426 118714 41461
rect 118743 41451 118789 41467
rect 118755 41399 118789 41451
rect 118869 41461 118917 42963
rect 120422 41484 120470 42968
rect 120550 42978 120584 43030
rect 121166 42996 121204 43000
rect 120550 42890 120596 42978
rect 121166 42962 121206 42996
rect 120598 42928 121206 42962
rect 121174 42922 121178 42928
rect 121202 42894 121206 42928
rect 121208 42978 121242 43030
rect 121208 42890 121254 42978
rect 121824 42962 121862 43000
rect 121256 42928 121862 42962
rect 121866 42968 121932 43030
rect 121956 42968 121960 43030
rect 121866 42922 121912 42968
rect 122482 42962 122520 43000
rect 121914 42928 122520 42962
rect 122524 42978 122558 43030
rect 123118 43000 123144 43030
rect 123146 43000 123216 43030
rect 123118 42978 123216 43000
rect 123798 42996 123836 43000
rect 120550 42878 120584 42890
rect 121183 42878 121196 42889
rect 121208 42878 121242 42890
rect 121841 42878 121854 42889
rect 121866 42878 121932 42922
rect 120536 41574 120584 42878
rect 115453 41365 118801 41399
rect 118869 36381 118903 41461
rect 118869 36132 118939 36381
rect 97493 34648 99222 34668
rect 115450 34657 118939 36132
rect 120422 36127 120456 41484
rect 120536 41422 120570 41574
rect 120572 41456 120576 41558
rect 121122 41530 121130 42342
rect 121150 41530 121158 42314
rect 121194 41574 121242 42878
rect 121852 41864 121932 42878
rect 121194 41562 121228 41574
rect 121852 41562 121906 41864
rect 121956 41836 121960 42922
rect 122524 42890 122570 42978
rect 123118 42968 123228 42978
rect 123140 42962 123178 42968
rect 122572 42928 123178 42962
rect 123182 42922 123228 42968
rect 123798 42962 123838 42996
rect 123230 42928 123838 42962
rect 123806 42922 123810 42928
rect 122499 42878 122512 42889
rect 122524 42878 122558 42890
rect 122510 41574 122558 42878
rect 123118 41800 123144 42922
rect 123146 42890 123228 42922
rect 123834 42894 123838 42928
rect 123146 41828 123216 42890
rect 123815 42878 123828 42889
rect 123840 42878 123874 43030
rect 123954 42968 123988 45978
rect 131924 45974 131944 46094
rect 131952 45968 131972 46122
rect 137156 45924 137176 46078
rect 137184 45930 137204 46050
rect 124606 44614 132582 44648
rect 125188 44032 126292 44052
rect 123134 41754 123144 41800
rect 123162 41754 123216 41828
rect 123750 41754 123756 42326
rect 123778 41754 123784 42298
rect 123168 41616 123216 41754
rect 122510 41562 122544 41574
rect 120600 41524 120604 41530
rect 121180 41524 121228 41562
rect 121838 41530 121892 41562
rect 121838 41524 121886 41530
rect 120596 41490 120604 41524
rect 120612 41490 121228 41524
rect 121254 41490 121262 41524
rect 121270 41490 121886 41524
rect 120600 41484 120604 41490
rect 121122 41478 121130 41484
rect 121150 41450 121158 41484
rect 121182 41474 121228 41490
rect 121840 41484 121886 41490
rect 121888 41484 121892 41530
rect 121916 41524 121920 41530
rect 122496 41524 122544 41562
rect 123134 41530 123144 41616
rect 123162 41574 123216 41616
rect 123162 41562 123202 41574
rect 123154 41524 123202 41562
rect 121912 41490 121920 41524
rect 121928 41490 122544 41524
rect 122570 41490 122578 41524
rect 122586 41490 123202 41524
rect 121916 41484 121920 41490
rect 121840 41474 121892 41484
rect 122498 41474 122544 41490
rect 121194 41422 121228 41474
rect 121852 41428 121892 41474
rect 121852 41422 121886 41428
rect 122510 41422 122544 41474
rect 123134 41422 123144 41484
rect 123156 41474 123202 41490
rect 123162 41422 123202 41474
rect 123204 41456 123208 41558
rect 123750 41530 123756 41616
rect 123778 41530 123784 41616
rect 123826 41574 123874 42878
rect 123826 41562 123860 41574
rect 123232 41524 123236 41530
rect 123812 41524 123860 41562
rect 123228 41490 123236 41524
rect 123244 41490 123860 41524
rect 123232 41484 123236 41490
rect 123750 41472 123756 41484
rect 123778 41450 123784 41484
rect 123814 41474 123860 41490
rect 123826 41422 123860 41474
rect 123940 41484 123988 42968
rect 124384 42954 127695 43095
rect 132666 43064 132668 43098
rect 124267 42923 127695 42954
rect 124384 42920 127695 42923
rect 124187 42542 124210 42904
rect 124233 42889 127695 42920
rect 124215 42542 124238 42876
rect 124384 41902 127695 42889
rect 129178 43030 132713 43064
rect 129178 42674 129212 43030
rect 129922 42962 129960 43000
rect 130580 42962 130618 43000
rect 131238 42962 131276 43000
rect 131896 42962 131934 43000
rect 132554 42962 132592 43000
rect 129354 42928 129960 42962
rect 130012 42928 130618 42962
rect 130670 42928 131276 42962
rect 131328 42928 131934 42962
rect 131986 42928 132592 42962
rect 132632 42918 132650 42928
rect 129281 42878 129326 42889
rect 129939 42878 129984 42889
rect 130597 42878 130642 42889
rect 131255 42878 131300 42889
rect 131913 42878 131958 42889
rect 129292 42674 129326 42878
rect 129337 42686 129338 42687
rect 129938 42686 129939 42687
rect 129338 42685 129339 42686
rect 129937 42685 129938 42686
rect 129950 42674 129984 42878
rect 129995 42686 129996 42687
rect 130596 42686 130597 42687
rect 129996 42685 129997 42686
rect 130595 42685 130596 42686
rect 130608 42674 130642 42878
rect 130653 42686 130654 42687
rect 131254 42686 131255 42687
rect 130654 42685 130655 42686
rect 131253 42685 131254 42686
rect 131266 42674 131300 42878
rect 131311 42686 131312 42687
rect 131912 42686 131913 42687
rect 131312 42685 131313 42686
rect 131911 42685 131912 42686
rect 131924 42674 131958 42878
rect 132548 42766 132566 42918
rect 132626 42916 132650 42918
rect 132598 42890 132616 42894
rect 132626 42890 132654 42916
rect 132576 42889 132654 42890
rect 132571 42878 132654 42889
rect 132576 42738 132654 42878
rect 132582 42702 132654 42738
rect 132582 42690 132650 42702
rect 131969 42686 131970 42687
rect 132570 42686 132571 42687
rect 131970 42685 131971 42686
rect 132569 42685 132570 42686
rect 132582 42674 132628 42690
rect 132632 42686 132650 42690
rect 132662 42686 132666 43030
rect 132696 42702 132713 43030
rect 129144 42671 132628 42674
rect 129144 42662 132622 42671
rect 129144 42652 132616 42662
rect 132696 42659 132700 42702
rect 129144 42650 132622 42652
rect 129144 42640 132628 42650
rect 129178 42016 129212 42640
rect 129292 42016 129326 42640
rect 129338 42628 129339 42629
rect 129937 42628 129938 42629
rect 129337 42627 129338 42628
rect 129938 42627 129939 42628
rect 129337 42028 129338 42029
rect 129938 42028 129939 42029
rect 129338 42027 129339 42028
rect 129937 42027 129938 42028
rect 129950 42016 129984 42640
rect 129996 42628 129997 42629
rect 130595 42628 130596 42629
rect 129995 42627 129996 42628
rect 130596 42627 130597 42628
rect 129995 42028 129996 42029
rect 130596 42028 130597 42029
rect 129996 42027 129997 42028
rect 130595 42027 130596 42028
rect 130608 42016 130642 42640
rect 130654 42628 130655 42629
rect 131253 42628 131254 42629
rect 130653 42627 130654 42628
rect 131254 42627 131255 42628
rect 130653 42028 130654 42029
rect 131254 42028 131255 42029
rect 130654 42027 130655 42028
rect 131253 42027 131254 42028
rect 131266 42016 131300 42640
rect 131312 42628 131313 42629
rect 131911 42628 131912 42629
rect 131311 42627 131312 42628
rect 131912 42627 131913 42628
rect 131311 42028 131312 42029
rect 131912 42028 131913 42029
rect 131312 42027 131313 42028
rect 131911 42027 131912 42028
rect 131924 42016 131958 42640
rect 131970 42628 131971 42629
rect 132569 42628 132570 42629
rect 131969 42627 131970 42628
rect 132570 42627 132571 42628
rect 132582 42624 132628 42640
rect 132632 42624 132650 42628
rect 132582 42612 132650 42624
rect 132582 42562 132654 42612
rect 131969 42028 131970 42029
rect 132570 42028 132571 42029
rect 131970 42027 131971 42028
rect 132569 42027 132570 42028
rect 132582 42016 132628 42562
rect 132632 42044 132654 42562
rect 132632 42028 132650 42044
rect 132662 42028 132666 42628
rect 132696 42044 132713 42659
rect 129144 42013 132628 42016
rect 129144 41982 132616 42013
rect 132696 41994 132700 42044
rect 129178 41902 129212 41982
rect 129292 41902 129326 41982
rect 129950 41902 129984 41982
rect 130608 41902 130642 41982
rect 131266 41902 131300 41982
rect 131924 41902 131958 41982
rect 132582 41902 132616 41982
rect 124384 41868 132628 41902
rect 132696 41868 132706 41936
rect 132734 41902 132768 43118
rect 154163 42667 154197 49031
rect 156909 45584 156943 48932
rect 156909 45232 156949 45584
rect 154277 42763 154311 42797
rect 154935 42763 154969 42797
rect 155593 42763 155627 42797
rect 156251 42763 156285 42797
rect 156909 42763 156943 45232
rect 157567 43059 157601 43093
rect 157681 43059 157715 49031
rect 160006 43095 160040 48946
rect 159198 43059 160605 43095
rect 162638 43064 162672 43098
rect 162752 43064 162786 49036
rect 157017 43025 160605 43059
rect 157017 42763 157051 43025
rect 157146 42957 157613 43004
rect 157193 42923 157613 42957
rect 157555 42876 157613 42923
rect 157120 42864 157176 42875
rect 157131 42763 157176 42864
rect 157567 42797 157612 42876
rect 157567 42763 157621 42797
rect 157681 42763 157715 43025
rect 159198 42804 160605 43025
rect 154227 42729 154231 42763
rect 154243 42729 157715 42763
rect 124384 41832 127695 41868
rect 120524 41388 123872 41422
rect 121194 36127 121228 41388
rect 121852 36127 121886 41388
rect 123134 41020 123144 41388
rect 123162 41020 123200 41388
rect 122576 40514 123168 40528
rect 123202 40514 123356 40528
rect 122610 40480 123168 40494
rect 123202 40480 123356 40494
rect 123134 38560 123144 39832
rect 123162 38560 123200 39832
rect 123134 37060 123144 37372
rect 123162 37060 123200 37372
rect 121894 36134 121918 36594
rect 121900 36127 121918 36134
rect 120386 34680 122759 36127
rect 123134 34862 123144 35156
rect 123162 34914 123200 35156
rect 123294 35100 123296 36614
rect 123162 34902 123202 34914
rect 123162 34890 123208 34902
rect 123940 34812 123974 41484
rect 124183 41412 124184 41498
rect 124221 41374 124222 41536
rect 124390 41494 124812 41832
rect 124866 41494 125288 41832
rect 127625 40349 127659 41832
rect 127660 41452 127695 41706
rect 127914 40990 127949 41452
rect 128370 41280 128472 41292
rect 129178 40385 129212 41868
rect 129254 41640 129268 41726
rect 129292 41602 129306 41764
rect 154131 40857 154197 42667
rect 154273 42677 154277 42695
rect 154273 42661 154323 42677
rect 154334 42667 154352 42682
rect 154362 42667 154380 42680
rect 154875 42661 154922 42708
rect 154931 42677 154935 42695
rect 154931 42661 154981 42677
rect 155533 42667 155580 42708
rect 155524 42661 155580 42667
rect 155589 42677 155593 42695
rect 155589 42661 155639 42677
rect 155654 42667 155660 42670
rect 155682 42667 155688 42680
rect 156191 42661 156238 42708
rect 156247 42677 156251 42695
rect 156247 42661 156297 42677
rect 156849 42667 156896 42708
rect 156909 42695 156943 42729
rect 156844 42661 156896 42667
rect 156905 42677 156943 42695
rect 156948 42677 156949 42729
rect 157017 42708 157051 42729
rect 157131 42726 157176 42729
rect 157567 42726 157612 42729
rect 157131 42708 157165 42726
rect 156905 42661 156955 42677
rect 157017 42661 157064 42708
rect 157131 42677 157178 42708
rect 157119 42661 157178 42677
rect 157507 42661 157554 42708
rect 154277 42627 154922 42661
rect 154935 42627 155580 42661
rect 155593 42627 156238 42661
rect 156251 42627 156896 42661
rect 156909 42627 157554 42661
rect 154277 42580 154323 42627
rect 154233 42568 154251 42580
rect 154277 42568 154311 42580
rect 154233 40944 154311 42568
rect 154334 41280 154352 42621
rect 154362 41252 154380 42621
rect 154935 42580 154981 42627
rect 155524 42621 155545 42627
rect 155552 42593 155573 42627
rect 155593 42580 155639 42627
rect 154892 42568 154923 42579
rect 154935 42568 154969 42580
rect 155550 42568 155581 42579
rect 155593 42568 155627 42580
rect 154832 40944 154842 42302
rect 154860 40944 154870 42274
rect 154903 40944 154969 42568
rect 155561 40944 155627 42568
rect 155654 41268 155660 42621
rect 155682 41240 155688 42621
rect 156251 42580 156297 42627
rect 156844 42621 156861 42627
rect 156872 42593 156889 42627
rect 156909 42621 156955 42627
rect 156909 42580 156980 42621
rect 156208 42568 156239 42579
rect 156251 42568 156285 42580
rect 156866 42568 156897 42579
rect 156909 42568 156943 42580
rect 156142 40944 156162 42308
rect 156170 40944 156190 42280
rect 156219 40944 156285 42568
rect 156877 40959 156943 42568
rect 156948 41246 156980 42580
rect 156948 40959 156949 41246
rect 157004 41218 157008 42621
rect 156877 40944 156949 40959
rect 157017 40944 157051 42627
rect 157119 42580 157177 42627
rect 157131 40944 157165 42580
rect 157567 42579 157601 42726
rect 157524 42568 157601 42579
rect 157535 40956 157601 42568
rect 157535 40944 157580 40956
rect 154233 40940 156598 40944
rect 154233 40930 154279 40940
rect 154292 40930 156598 40940
rect 154233 40906 156598 40930
rect 154131 40454 154165 40857
rect 154233 40795 154279 40906
rect 154292 40897 156598 40906
rect 156865 40897 156924 40944
rect 157017 40897 157064 40944
rect 157131 40897 157178 40944
rect 157535 40897 157582 40944
rect 154339 40863 154950 40897
rect 154985 40894 155608 40897
rect 154997 40863 155608 40894
rect 155655 40863 156266 40897
rect 156313 40863 156924 40897
rect 156971 40863 157582 40897
rect 154891 40847 154937 40863
rect 155549 40847 155595 40863
rect 156207 40847 156253 40863
rect 156865 40857 156911 40863
rect 156865 40847 156917 40857
rect 156877 40801 156917 40847
rect 156877 40795 156911 40801
rect 157017 40795 157051 40863
rect 157131 40795 157165 40863
rect 157535 40795 157569 40863
rect 157649 40795 157715 42729
rect 159166 42768 160605 42804
rect 162088 43030 165544 43064
rect 160664 42768 160698 42802
rect 161322 42768 161356 42802
rect 161980 42768 162014 42802
rect 162088 42768 162122 43030
rect 162638 42993 162676 43000
rect 162638 42978 162684 42993
rect 162626 42962 162684 42978
rect 162264 42928 162684 42962
rect 162626 42890 162684 42928
rect 162191 42878 162236 42889
rect 162202 42768 162236 42878
rect 162638 42802 162672 42890
rect 162638 42768 162692 42802
rect 162752 42768 162786 43030
rect 159166 42734 162786 42768
rect 159166 42704 160605 42734
rect 159166 42662 160642 42704
rect 160658 42682 160672 42728
rect 160658 42672 160710 42682
rect 160660 42666 160710 42672
rect 161262 42666 161300 42704
rect 161318 42682 161322 42700
rect 161318 42666 161368 42682
rect 161920 42666 161958 42704
rect 161976 42682 161980 42700
rect 162018 42682 162020 42734
rect 162088 42704 162122 42734
rect 162202 42704 162236 42734
rect 161976 42666 162026 42682
rect 162088 42666 162126 42704
rect 162202 42682 162240 42704
rect 162190 42666 162248 42682
rect 162578 42666 162616 42704
rect 159166 42632 160644 42662
rect 159166 42626 160616 42632
rect 157746 41218 157752 42570
rect 158512 41562 158550 41762
rect 158568 41534 158578 41790
rect 154233 40761 157715 40795
rect 159166 40920 160605 42626
rect 160622 42598 160644 42632
rect 160664 42632 161300 42666
rect 161322 42632 161958 42666
rect 161980 42632 162616 42666
rect 160622 42593 160636 42598
rect 160664 42594 160710 42632
rect 161322 42594 161368 42632
rect 161980 42626 162026 42632
rect 162088 42626 162122 42632
rect 161980 42594 162052 42626
rect 160621 42582 160652 42593
rect 160664 42582 160698 42594
rect 161279 42582 161310 42593
rect 161322 42582 161356 42594
rect 161937 42582 161968 42593
rect 161980 42582 162014 42594
rect 160622 41260 160698 42582
rect 160626 40970 160698 41260
rect 160626 40958 160666 40970
rect 160620 40920 160670 40958
rect 161222 40926 161238 41858
rect 161250 40926 161266 41858
rect 161290 40970 161356 42582
rect 161366 41168 161386 41858
rect 161948 40982 162014 42582
rect 162018 41224 162052 42594
rect 162018 40982 162020 41224
rect 162074 41168 162122 42626
rect 162190 42594 162248 42632
rect 161290 40958 161324 40970
rect 161948 40958 162020 40982
rect 162088 40958 162122 41168
rect 162202 40958 162236 42594
rect 162638 42593 162672 42734
rect 162595 42582 162672 42593
rect 162606 40970 162672 42582
rect 161278 40920 161328 40958
rect 161936 40926 161988 40958
rect 161936 40920 161986 40926
rect 162088 40920 162126 40958
rect 162202 40920 162240 40958
rect 162606 40954 162651 40970
rect 162606 40920 162644 40954
rect 159166 40886 160670 40920
rect 160726 40886 161328 40920
rect 161384 40886 161986 40920
rect 162042 40886 162644 40920
rect 159166 40818 160605 40886
rect 160620 40870 160666 40886
rect 161278 40870 161324 40886
rect 161936 40880 161982 40886
rect 161936 40870 161988 40880
rect 161948 40824 161988 40870
rect 161948 40818 161982 40824
rect 162088 40818 162122 40886
rect 162202 40822 162236 40886
rect 162606 40822 162640 40886
rect 162202 40818 162247 40822
rect 162606 40818 162651 40822
rect 162720 40818 162786 42734
rect 162822 42314 162838 42316
rect 162816 41210 162838 42314
rect 162860 42218 162894 42878
rect 162860 42136 162960 42218
rect 162822 40926 162838 41126
rect 159166 40784 162786 40818
rect 154245 40454 154279 40488
rect 154903 40454 154937 40488
rect 155561 40454 155595 40488
rect 156219 40454 156253 40488
rect 152946 40420 156402 40454
rect 129142 40349 132766 40385
rect 124425 40315 132766 40349
rect 124425 36831 124459 40315
rect 124879 40314 124913 40315
rect 124879 40241 124919 40314
rect 124938 40241 124947 40286
rect 124879 40235 124913 40241
rect 125537 40235 125571 40315
rect 126195 40235 126229 40315
rect 126853 40235 126887 40315
rect 127511 40235 127545 40315
rect 127625 40235 127659 40315
rect 124480 40173 124561 40220
rect 124620 40201 127659 40235
rect 124879 40195 124913 40201
rect 124866 40189 124867 40190
rect 124867 40188 124868 40189
rect 124527 39605 124561 40173
rect 124879 40130 124919 40195
rect 124925 40189 124926 40190
rect 124924 40188 124925 40189
rect 124938 40158 124947 40195
rect 125524 40189 125525 40190
rect 125525 40188 125526 40189
rect 124867 39589 124868 39590
rect 124866 39588 124867 39589
rect 124879 39577 124913 40130
rect 124924 39589 124925 39590
rect 125525 39589 125526 39590
rect 124925 39588 124926 39589
rect 125524 39588 125525 39589
rect 125537 39577 125571 40201
rect 125583 40189 125584 40190
rect 126182 40189 126183 40190
rect 125582 40188 125583 40189
rect 126183 40188 126184 40189
rect 125582 39589 125583 39590
rect 126183 39589 126184 39590
rect 125583 39588 125584 39589
rect 126182 39588 126183 39589
rect 126195 39577 126229 40201
rect 126241 40189 126242 40190
rect 126840 40189 126841 40190
rect 126240 40188 126241 40189
rect 126841 40188 126842 40189
rect 126240 39589 126241 39590
rect 126841 39589 126842 39590
rect 126241 39588 126242 39589
rect 126840 39588 126841 39589
rect 126853 39577 126887 40201
rect 126899 40189 126900 40190
rect 127498 40189 127499 40190
rect 126898 40188 126899 40189
rect 127499 40188 127500 40189
rect 126898 39589 126899 39590
rect 127499 39589 127500 39590
rect 126899 39588 126900 39589
rect 127498 39588 127499 39589
rect 127511 39577 127545 40201
rect 127625 39577 127659 40201
rect 129142 39577 132784 40315
rect 145984 40290 145988 40295
rect 145914 40262 145960 40267
rect 145914 40255 145982 40262
rect 145920 40252 145982 40255
rect 124480 39515 124561 39562
rect 124620 39543 132784 39577
rect 124866 39531 124867 39532
rect 124867 39530 124868 39531
rect 124527 38947 124561 39515
rect 124867 38931 124868 38932
rect 124866 38930 124867 38931
rect 124879 38919 124913 39543
rect 124925 39531 124926 39532
rect 125524 39531 125525 39532
rect 124924 39530 124925 39531
rect 125525 39530 125526 39531
rect 125537 38934 125571 39543
rect 125583 39531 125584 39532
rect 126182 39531 126183 39532
rect 125582 39530 125583 39531
rect 126183 39530 126184 39531
rect 125762 38934 125974 39066
rect 124924 38931 124925 38932
rect 124925 38930 124926 38931
rect 125452 38919 125974 38934
rect 126183 38931 126184 38932
rect 126182 38930 126183 38931
rect 126195 38919 126229 39543
rect 126241 39531 126242 39532
rect 126840 39531 126841 39532
rect 126240 39530 126241 39531
rect 126841 39530 126842 39531
rect 126240 38931 126241 38932
rect 126841 38931 126842 38932
rect 126241 38930 126242 38931
rect 126840 38930 126841 38931
rect 126853 38919 126887 39543
rect 126899 39531 126900 39532
rect 127498 39531 127499 39532
rect 126898 39530 126899 39531
rect 127499 39530 127500 39531
rect 126898 38931 126899 38932
rect 127499 38931 127500 38932
rect 126899 38930 126900 38931
rect 127498 38930 127499 38931
rect 127511 38919 127545 39543
rect 127625 38919 127659 39543
rect 128336 39500 128726 39534
rect 127690 39018 127946 39024
rect 128336 39002 128370 39500
rect 128550 39432 128597 39479
rect 128512 39398 128597 39432
rect 128439 39339 128484 39350
rect 128567 39339 128612 39350
rect 128450 39163 128484 39339
rect 128578 39163 128612 39339
rect 128550 39104 128597 39151
rect 128512 39070 128597 39104
rect 128692 39002 128726 39500
rect 128846 39018 129102 39036
rect 127718 38990 127918 38996
rect 128336 38968 128726 39002
rect 128874 38990 129074 39008
rect 124480 38857 124561 38904
rect 124620 38885 127659 38919
rect 124866 38873 124867 38874
rect 124867 38872 124868 38873
rect 124527 38289 124561 38857
rect 124867 38273 124868 38274
rect 124866 38272 124867 38273
rect 124879 38261 124913 38885
rect 124925 38873 124926 38874
rect 124924 38872 124925 38873
rect 125452 38864 125974 38885
rect 126182 38873 126183 38874
rect 126183 38872 126184 38873
rect 124919 38836 124996 38852
rect 125444 38836 125531 38852
rect 124924 38273 124925 38274
rect 125525 38273 125526 38274
rect 124925 38272 124926 38273
rect 125524 38272 125525 38273
rect 125537 38261 125571 38864
rect 125577 38836 125658 38852
rect 125762 38618 125974 38864
rect 126106 38836 126189 38852
rect 125582 38273 125583 38274
rect 126183 38273 126184 38274
rect 125583 38272 125584 38273
rect 126182 38272 126183 38273
rect 126195 38261 126229 38885
rect 126241 38873 126242 38874
rect 126840 38873 126841 38874
rect 126240 38872 126241 38873
rect 126841 38872 126842 38873
rect 126235 38836 126260 38852
rect 126240 38273 126241 38274
rect 126841 38273 126842 38274
rect 126241 38272 126242 38273
rect 126840 38272 126841 38273
rect 126853 38261 126887 38885
rect 126899 38873 126900 38874
rect 127498 38873 127499 38874
rect 126898 38872 126899 38873
rect 127499 38872 127500 38873
rect 126898 38273 126899 38274
rect 127499 38273 127500 38274
rect 126899 38272 126900 38273
rect 127498 38272 127499 38273
rect 127511 38261 127545 38885
rect 127625 38261 127659 38885
rect 127918 38804 128178 38824
rect 127918 38776 128178 38796
rect 128322 38298 128744 38918
rect 128874 38808 129074 38824
rect 128846 38780 129102 38796
rect 129142 38261 132784 39543
rect 143762 38841 144198 38864
rect 143796 38807 144164 38830
rect 144669 38742 144703 40209
rect 145928 40070 145982 40252
rect 145928 39782 145960 40070
rect 145920 39779 145960 39782
rect 145914 39767 145960 39779
rect 145984 40042 146010 40290
rect 147230 40264 147276 40267
rect 147212 40255 147276 40264
rect 153658 40266 153662 40271
rect 147212 40252 147270 40255
rect 147212 40078 147228 40252
rect 153658 40080 153686 40266
rect 145984 39739 145988 40042
rect 147230 39779 147270 39782
rect 147230 39767 147276 39779
rect 145982 39686 146550 39720
rect 148754 39420 148978 39440
rect 150946 39424 151166 39444
rect 148774 39268 148775 39420
rect 148958 39268 148978 39420
rect 150966 39268 150967 39424
rect 151146 39268 151166 39424
rect 153658 39228 153662 40080
rect 144126 38708 146266 38742
rect 137936 38304 137992 38306
rect 124480 38199 124561 38246
rect 124620 38227 132784 38261
rect 124866 38215 124867 38216
rect 124867 38214 124868 38215
rect 124527 37631 124561 38199
rect 124867 37615 124868 37616
rect 124866 37614 124867 37615
rect 124879 37603 124913 38227
rect 124925 38215 124926 38216
rect 125524 38215 125525 38216
rect 124924 38214 124925 38215
rect 125525 38214 125526 38215
rect 124924 37615 124925 37616
rect 125525 37615 125526 37616
rect 124925 37614 124926 37615
rect 125524 37614 125525 37615
rect 125537 37603 125571 38227
rect 125583 38215 125584 38216
rect 126182 38215 126183 38216
rect 125582 38214 125583 38215
rect 126183 38214 126184 38215
rect 125582 37615 125583 37616
rect 126183 37615 126184 37616
rect 125583 37614 125584 37615
rect 126182 37614 126183 37615
rect 126195 37603 126229 38227
rect 126241 38215 126242 38216
rect 126840 38215 126841 38216
rect 126240 38214 126241 38215
rect 126841 38214 126842 38215
rect 126240 37615 126241 37616
rect 126841 37615 126842 37616
rect 126241 37614 126242 37615
rect 126840 37614 126841 37615
rect 126853 37603 126887 38227
rect 126899 38215 126900 38216
rect 127498 38215 127499 38216
rect 126898 38214 126899 38215
rect 127499 38214 127500 38215
rect 126898 37615 126899 37616
rect 127499 37615 127500 37616
rect 126899 37614 126900 37615
rect 127498 37614 127499 37615
rect 127511 37603 127545 38227
rect 127625 37603 127659 38227
rect 128886 38156 128928 38162
rect 129066 38156 129094 38162
rect 128858 38128 128928 38134
rect 129066 38128 129122 38134
rect 129142 37603 132784 38227
rect 144126 38217 144160 38708
rect 144567 38640 144601 38708
rect 144669 38640 144703 38708
rect 144302 38606 144703 38640
rect 144519 38559 144520 38560
rect 144520 38558 144521 38559
rect 144229 38547 144274 38558
rect 144240 38217 144274 38547
rect 144567 38245 144601 38606
rect 144285 38229 144286 38230
rect 144286 38228 144287 38229
rect 144508 38217 144519 38228
rect 144092 38183 144519 38217
rect 137936 38142 137992 38146
rect 137936 38086 137992 38090
rect 124480 37541 124561 37588
rect 124620 37569 132784 37603
rect 124866 37557 124867 37558
rect 124867 37556 124868 37557
rect 124527 36973 124561 37541
rect 124867 36957 124868 36958
rect 124866 36956 124867 36957
rect 124879 36945 124913 37569
rect 124925 37557 124926 37558
rect 125524 37557 125525 37558
rect 124924 37556 124925 37557
rect 125525 37556 125526 37557
rect 124924 36957 124925 36958
rect 125525 36957 125526 36958
rect 124925 36956 124926 36957
rect 125524 36956 125525 36957
rect 125537 36945 125571 37569
rect 125583 37557 125584 37558
rect 126182 37557 126183 37558
rect 125582 37556 125583 37557
rect 126183 37556 126184 37557
rect 125582 36957 125583 36958
rect 126183 36957 126184 36958
rect 125583 36956 125584 36957
rect 126182 36956 126183 36957
rect 126195 36945 126229 37569
rect 126241 37557 126242 37558
rect 126840 37557 126841 37558
rect 126240 37556 126241 37557
rect 126841 37556 126842 37557
rect 126240 36957 126241 36958
rect 126841 36957 126842 36958
rect 126241 36956 126242 36957
rect 126840 36956 126841 36957
rect 126853 36945 126887 37569
rect 126899 37557 126900 37558
rect 127498 37557 127499 37558
rect 126898 37556 126899 37557
rect 127499 37556 127500 37557
rect 126898 36957 126899 36958
rect 127499 36957 127500 36958
rect 126899 36956 126900 36957
rect 127498 36956 127499 36957
rect 127511 36945 127545 37569
rect 127625 36945 127659 37569
rect 128324 37563 128580 37569
rect 128352 37535 128552 37554
rect 124620 36911 127659 36945
rect 124879 36831 124913 36911
rect 125537 36831 125571 36911
rect 126195 36831 126229 36911
rect 126853 36831 126887 36911
rect 127511 36831 127545 36911
rect 127625 36831 127659 36911
rect 129142 36831 132784 37569
rect 144126 37559 144160 38183
rect 144240 37571 144274 38183
rect 144286 38171 144287 38172
rect 144285 38170 144286 38171
rect 144520 38155 144601 38202
rect 144285 37571 144286 37572
rect 144286 37570 144287 37571
rect 144304 37570 144306 37593
rect 144567 37587 144601 38155
rect 144304 37559 144334 37565
rect 144508 37559 144519 37570
rect 144092 37525 144194 37559
rect 144202 37546 144520 37559
rect 144202 37533 144524 37546
rect 144252 37525 144524 37533
rect 144126 37410 144160 37525
rect 144262 37519 144520 37525
rect 144286 37513 144520 37519
rect 144290 37512 144342 37513
rect 144669 37512 144703 38606
rect 147444 38350 147468 38560
rect 145598 37834 145622 37842
rect 145598 37582 145624 37834
rect 145598 37570 145622 37582
rect 144286 37491 144703 37512
rect 144302 37478 144703 37491
rect 144567 37410 144601 37478
rect 144669 37410 144703 37478
rect 124425 36797 132766 36831
rect 127625 36482 127659 36797
rect 129142 36761 132766 36797
rect 124384 36446 127695 36482
rect 129178 36446 129212 36761
rect 131296 36496 131300 36658
rect 131334 36534 131338 36620
rect 124384 36412 132628 36446
rect 132696 36412 132706 36480
rect 124282 36132 124296 36270
rect 124384 36132 127695 36412
rect 129178 36332 129212 36412
rect 129292 36332 129326 36412
rect 129338 36332 129938 36343
rect 129950 36332 129984 36412
rect 129996 36332 130596 36343
rect 130608 36332 130642 36412
rect 130654 36332 131254 36343
rect 131266 36332 131300 36412
rect 131312 36332 131912 36343
rect 131924 36332 131958 36412
rect 131970 36332 132570 36343
rect 132582 36332 132616 36412
rect 132700 36350 132730 36384
rect 129144 36310 132616 36332
rect 129144 36308 132622 36310
rect 129144 36298 132628 36308
rect 124206 36096 127695 36132
rect 124206 36062 127794 36096
rect 124206 35674 127695 36062
rect 127760 35674 127794 36062
rect 128464 35928 128912 36090
rect 128388 35878 128912 35928
rect 128388 35774 128542 35878
rect 129178 35674 129212 36298
rect 129292 36286 129326 36298
rect 129338 36286 129339 36287
rect 129937 36286 129938 36287
rect 129950 36286 129984 36298
rect 129996 36286 129997 36287
rect 130595 36286 130596 36287
rect 130608 36286 130642 36298
rect 130654 36286 130655 36287
rect 131253 36286 131254 36287
rect 131266 36286 131300 36298
rect 131312 36286 131313 36287
rect 131911 36286 131912 36287
rect 131924 36286 131958 36298
rect 131970 36286 131971 36287
rect 132569 36286 132570 36287
rect 129292 36285 129338 36286
rect 129938 36285 129939 36286
rect 129950 36285 129996 36286
rect 130596 36285 130597 36286
rect 130608 36285 130654 36286
rect 131254 36285 131255 36286
rect 131266 36285 131312 36286
rect 131912 36285 131913 36286
rect 131924 36285 131970 36286
rect 132570 36285 132571 36286
rect 129292 36127 129337 36285
rect 129950 36127 129995 36285
rect 130608 36127 130653 36285
rect 131266 36127 131311 36285
rect 131924 36127 131969 36285
rect 132582 36282 132628 36298
rect 132582 36270 132650 36282
rect 132582 36214 132654 36270
rect 132582 36127 132628 36214
rect 132632 36127 132654 36214
rect 132696 36127 132713 36317
rect 132734 36127 132768 36412
rect 129283 35674 132804 36127
rect 132860 36094 132907 36127
rect 124206 35640 127794 35674
rect 129144 35640 132804 35674
rect 124206 35016 127695 35640
rect 127760 35016 127794 35640
rect 129178 35016 129212 35640
rect 129283 35016 132804 35640
rect 133114 35456 133161 36094
rect 133340 36058 133374 37384
rect 144126 37376 146266 37410
rect 136424 36950 137044 37372
rect 137094 37324 137660 37358
rect 137094 37002 137128 37324
rect 137465 37244 137476 37255
rect 137149 37182 137230 37229
rect 137289 37210 137476 37244
rect 137477 37182 137558 37229
rect 137196 37144 137230 37182
rect 137524 37144 137558 37182
rect 137465 37116 137476 37127
rect 137289 37082 137476 37116
rect 137626 37002 137660 37324
rect 144669 37192 144703 37376
rect 137094 36968 137660 37002
rect 136482 36896 136500 36935
rect 136800 36907 136830 36942
rect 136856 36907 136858 36942
rect 137472 36928 137992 36942
rect 136516 36896 136534 36901
rect 136830 36896 136856 36907
rect 136424 36850 137044 36896
rect 137156 36882 137598 36916
rect 137094 36855 137660 36882
rect 136424 36848 137104 36850
rect 136424 36834 137162 36848
rect 136424 36822 137044 36834
rect 136424 36820 137076 36822
rect 136424 36787 137134 36820
rect 136424 36753 141848 36787
rect 136424 36717 137044 36753
rect 137094 36620 137134 36753
rect 137142 36626 137162 36746
rect 137196 36719 137230 36722
rect 137524 36719 137558 36722
rect 137094 36588 137128 36620
rect 137626 36588 137660 36753
rect 144114 36717 144739 37192
rect 134354 36096 135696 36132
rect 136282 36126 136500 36130
rect 136936 36096 136970 36212
rect 137112 36172 141848 36206
rect 137060 36144 137118 36162
rect 137050 36134 137084 36138
rect 137000 36108 137044 36118
rect 137050 36116 137090 36134
rect 137050 36096 137084 36116
rect 137628 36108 137850 36130
rect 133454 36058 133478 36092
rect 134354 36072 137942 36096
rect 142222 36072 142256 36212
rect 144150 36072 144184 36717
rect 145494 36696 145514 36978
rect 134354 36062 144666 36072
rect 133246 36024 133540 36058
rect 133340 35990 133374 36024
rect 133340 35922 133398 35990
rect 133472 35962 133488 35996
rect 133340 35662 133374 35922
rect 133392 35687 133408 35863
rect 133416 35687 133426 35863
rect 133442 35700 133492 35929
rect 133442 35675 133500 35700
rect 133340 35594 133398 35662
rect 133340 35526 133374 35594
rect 133444 35526 133500 35675
rect 133506 35526 133540 36024
rect 133246 35492 133540 35526
rect 133626 36024 134016 36058
rect 133626 35526 133660 36024
rect 133840 35956 133887 36003
rect 133802 35922 133887 35956
rect 133729 35863 133774 35874
rect 133857 35863 133902 35874
rect 133740 35687 133774 35863
rect 133868 35687 133902 35863
rect 133840 35628 133887 35675
rect 133802 35594 133887 35628
rect 133982 35526 134016 36024
rect 133626 35492 134016 35526
rect 133340 35442 133374 35492
rect 133444 35490 133500 35492
rect 133380 35442 133500 35490
rect 133304 35078 133554 35442
rect 133608 35078 134030 35442
rect 134354 35078 135696 36062
rect 136414 36041 144666 36062
rect 136318 36038 144666 36041
rect 136318 36010 136352 36038
rect 136284 35994 136386 36010
rect 136936 35994 136970 36038
rect 137050 36025 137088 36032
rect 137038 36010 137088 36025
rect 137038 35994 137096 36010
rect 137108 35994 137146 36032
rect 137766 35994 137804 36032
rect 124206 34982 127794 35016
rect 129144 34982 132804 35016
rect 133610 35004 133642 35078
rect 133644 35004 133676 35078
rect 133758 35028 133792 35038
rect 133846 35028 133880 35038
rect 133724 34994 133914 35004
rect 97493 34640 99144 34648
rect 97493 34620 99194 34640
rect 97493 34565 99144 34620
rect 97493 34531 101528 34565
rect 97493 34381 99144 34531
rect 97804 34380 98352 34381
rect 98402 34326 99040 34381
rect 98334 34214 98338 34216
rect 98976 33996 98994 34154
rect 99014 34030 99032 34116
rect 99074 33996 99108 34381
rect 98976 33992 99194 33996
rect 98994 33978 99194 33992
rect 99074 33962 99108 33978
rect 98994 33944 99228 33962
rect 99074 33942 99108 33944
rect 97662 33908 101528 33942
rect 82678 33228 83052 33262
rect 83104 33228 83810 33262
rect 83862 33228 84568 33262
rect 84608 33262 84710 33268
rect 84731 33262 93169 33268
rect 84608 33228 93169 33262
rect 94350 33244 94396 33268
rect 82678 33212 82736 33228
rect 83336 33212 83394 33228
rect 83994 33212 84052 33228
rect 84608 33222 84636 33228
rect 84652 33212 84710 33228
rect 82678 33197 82693 33212
rect 82690 33160 82724 33194
rect 83348 33160 83382 33194
rect 84006 33160 84040 33194
rect 84664 33160 84698 33194
rect 84731 33160 93169 33228
rect 94358 33222 94396 33244
rect 94414 33194 94424 33296
rect 97662 33262 97696 33908
rect 98202 33828 98236 33908
rect 98364 33828 98948 33839
rect 98960 33828 98994 33908
rect 99074 33828 99108 33908
rect 105836 33834 105852 33940
rect 97726 33766 97798 33804
rect 97848 33794 99142 33828
rect 98189 33782 98190 33783
rect 98190 33781 98191 33782
rect 97764 33262 97798 33766
rect 98202 33312 98236 33794
rect 98248 33782 98249 33783
rect 98947 33782 98948 33783
rect 98960 33782 98994 33794
rect 98247 33781 98248 33782
rect 98948 33781 98949 33782
rect 98960 33518 99005 33782
rect 99074 33518 99108 33794
rect 105826 33788 105852 33834
rect 105836 33710 105852 33788
rect 105854 33760 105864 33862
rect 105854 33716 105868 33738
rect 105826 33688 105868 33710
rect 97835 33300 97836 33301
rect 97836 33299 97837 33300
rect 98174 33262 98212 33300
rect 98510 33262 101476 33518
rect 97662 33228 98212 33262
rect 98264 33236 101476 33262
rect 97662 33160 97696 33228
rect 97764 33198 97798 33228
rect 98074 33222 98186 33228
rect 98252 33222 101476 33236
rect 98510 33208 101476 33222
rect 98102 33194 98214 33208
rect 98224 33194 101476 33208
rect 97764 33182 97798 33194
rect 97848 33160 101476 33194
rect 72267 33126 72355 33160
rect 73042 33126 101476 33160
rect 72267 33090 72337 33126
rect 73042 33090 82550 33126
rect 41048 31341 47423 31375
rect 45678 31261 45712 31341
rect 45792 31261 45826 31341
rect 47228 31261 47239 31272
rect 45644 31227 47239 31261
rect 45678 30814 45712 31227
rect 45792 30814 45826 31227
rect 45838 31215 45839 31216
rect 45837 31214 45838 31215
rect 47240 31199 47321 31246
rect 45678 30622 45950 30814
rect 47287 30631 47321 31199
rect 45678 30603 46532 30622
rect 47228 30603 47239 30614
rect 45644 30569 47239 30603
rect 45678 30548 46532 30569
rect 45678 30370 45950 30548
rect 46030 30532 46086 30548
rect 47240 30541 47321 30588
rect 46030 30476 46086 30492
rect 45678 29945 45712 30370
rect 45792 29945 45826 30370
rect 47287 29973 47321 30541
rect 45837 29957 45838 29958
rect 45838 29956 45839 29957
rect 47228 29945 47239 29956
rect 45644 29911 47239 29945
rect 45678 29287 45712 29911
rect 45792 29287 45826 29911
rect 45838 29899 45839 29900
rect 45837 29898 45838 29899
rect 47240 29883 47321 29930
rect 46030 29374 46086 29376
rect 46030 29318 46086 29320
rect 47287 29315 47321 29883
rect 45837 29299 45838 29300
rect 45838 29298 45839 29299
rect 47228 29287 47239 29298
rect 45644 29253 47239 29287
rect 45678 29078 45712 29253
rect 45792 29239 45826 29253
rect 45838 29241 45839 29242
rect 45837 29240 45838 29241
rect 47240 29227 47368 29272
rect 47239 29226 47240 29227
rect 45814 29212 46086 29214
rect 45842 29184 46086 29186
rect 46030 29180 46086 29184
rect 47287 29180 47321 29225
rect 47389 29180 47423 31341
rect 55002 31032 55006 31288
rect 55030 31060 55034 31260
rect 55080 31001 55114 31664
rect 55166 31642 55404 31664
rect 45854 29146 47423 29180
rect 47287 29078 47321 29146
rect 47389 29078 47423 29146
rect 50927 30994 59197 31001
rect 50927 30967 59293 30994
rect 50927 29180 50961 30967
rect 51908 30887 51942 30967
rect 54966 30887 55000 30967
rect 55080 30887 55114 30967
rect 57752 30887 57786 30967
rect 57935 30949 58836 30967
rect 57935 30942 59166 30949
rect 57854 30933 57888 30936
rect 57854 30920 57888 30921
rect 57907 30914 58780 30938
rect 50982 30825 51063 30872
rect 51122 30853 55114 30887
rect 57718 30853 57786 30887
rect 57807 30887 57935 30899
rect 59098 30887 59109 30898
rect 57807 30853 59109 30887
rect 51895 30841 51896 30842
rect 51896 30840 51897 30841
rect 51029 30257 51063 30825
rect 51908 30260 51942 30853
rect 51954 30841 51955 30842
rect 54953 30841 54954 30842
rect 51953 30840 51954 30841
rect 54954 30840 54955 30841
rect 51806 30254 52082 30260
rect 51896 30241 51897 30242
rect 51895 30240 51896 30241
rect 51908 30229 51942 30254
rect 51953 30241 51954 30242
rect 54954 30241 54955 30242
rect 51954 30240 51955 30241
rect 54953 30240 54954 30241
rect 54966 30229 55000 30853
rect 55080 30229 55114 30853
rect 57752 30229 57786 30853
rect 57838 30841 57935 30853
rect 57854 30352 57888 30841
rect 59110 30825 59191 30872
rect 59157 30337 59191 30825
rect 59110 30336 59191 30337
rect 59110 30324 59207 30336
rect 59259 30324 59293 30967
rect 60518 30374 60574 30386
rect 61762 30374 61818 30386
rect 60518 30324 60574 30330
rect 57807 30274 57888 30309
rect 57947 30291 61208 30324
rect 61762 30318 61818 30330
rect 57935 30290 61208 30291
rect 57935 30284 59207 30290
rect 58866 30278 59207 30284
rect 58866 30274 59191 30278
rect 57807 30262 57894 30274
rect 57854 30242 57894 30262
rect 59151 30257 59191 30274
rect 59151 30248 59166 30257
rect 59151 30245 59197 30248
rect 50982 30167 51063 30214
rect 51122 30195 55114 30229
rect 57718 30195 57786 30229
rect 57807 30241 57894 30242
rect 57807 30235 57935 30241
rect 57807 30229 58866 30235
rect 59098 30229 59109 30240
rect 57807 30195 59109 30229
rect 59123 30217 59225 30220
rect 51895 30183 51896 30184
rect 51896 30182 51897 30183
rect 51029 29599 51063 30167
rect 51556 30158 51612 30174
rect 51556 30102 51612 30118
rect 51896 29583 51897 29584
rect 51895 29582 51896 29583
rect 51908 29571 51942 30195
rect 51954 30183 51955 30184
rect 54953 30183 54954 30184
rect 51953 30182 51954 30183
rect 54954 30182 54955 30183
rect 52182 30158 52238 30174
rect 52182 30102 52238 30118
rect 51953 29583 51954 29584
rect 54954 29583 54955 29584
rect 51954 29582 51955 29583
rect 54953 29582 54954 29583
rect 54966 29571 55000 30195
rect 55080 29571 55114 30195
rect 57752 29571 57786 30195
rect 57838 30183 57935 30195
rect 57854 29694 57888 30183
rect 59110 30167 59191 30214
rect 59157 29679 59191 30167
rect 59110 29678 59191 29679
rect 57792 29670 58866 29672
rect 57935 29666 58866 29670
rect 59110 29666 59207 29678
rect 57807 29616 57888 29651
rect 57935 29626 59207 29666
rect 59110 29620 59207 29626
rect 57807 29604 58810 29616
rect 57854 29584 58810 29604
rect 59151 29599 59191 29620
rect 59151 29588 59166 29599
rect 59151 29587 59197 29588
rect 50982 29509 51063 29556
rect 51122 29537 55114 29571
rect 57718 29537 57786 29571
rect 57807 29577 58810 29584
rect 59098 29577 59109 29582
rect 57807 29570 59110 29577
rect 57807 29537 59109 29570
rect 59123 29559 59225 29560
rect 51895 29525 51896 29526
rect 51896 29524 51897 29525
rect 51029 29180 51063 29509
rect 51908 29239 51942 29537
rect 51954 29525 51955 29526
rect 54953 29525 54954 29526
rect 51953 29524 51954 29525
rect 54954 29524 54955 29525
rect 54966 29239 55000 29537
rect 51109 29227 51110 29228
rect 51110 29226 51111 29227
rect 51880 29180 51927 29227
rect 54938 29180 54985 29227
rect 50927 29146 51927 29180
rect 51970 29146 54985 29180
rect 50927 29078 50961 29146
rect 51029 29078 51063 29146
rect 55080 29078 55114 29537
rect 45678 29044 55114 29078
rect 47389 28424 47423 29044
rect 50927 28424 50961 29044
rect 52182 28944 52836 28946
rect 57752 28894 57786 29537
rect 57838 29525 57935 29537
rect 57854 29036 57888 29525
rect 59110 29509 59191 29556
rect 59157 29021 59191 29509
rect 59110 29020 59191 29021
rect 59110 29008 59207 29020
rect 57947 28977 59207 29008
rect 57947 28974 59222 28977
rect 59110 28962 59222 28974
rect 57814 28894 59098 28928
rect 59157 28925 59191 28928
rect 59259 28894 59293 30290
rect 60518 29714 60574 29728
rect 61762 29714 61818 29728
rect 60518 29658 60574 29672
rect 61762 29658 61818 29672
rect 60518 29054 60574 29070
rect 61762 29054 61818 29070
rect 60518 28998 60574 29014
rect 61762 28998 61818 29014
rect 57752 28860 61208 28894
rect 59259 28466 59293 28860
rect 57752 28432 61208 28466
rect 45714 28390 55150 28424
rect 45714 27971 45748 28390
rect 47287 28322 47321 28390
rect 47389 28322 47423 28390
rect 45890 28288 47423 28322
rect 47239 28241 47240 28242
rect 47240 28240 47241 28241
rect 45817 28229 45862 28240
rect 45828 27971 45862 28229
rect 46108 28054 46164 28068
rect 47287 27999 47321 28288
rect 45873 27983 45874 27984
rect 45874 27982 45875 27983
rect 47228 27971 47239 27982
rect 45680 27937 47239 27971
rect 45714 27857 45748 27937
rect 45828 27857 45862 27937
rect 47389 27857 47423 28288
rect 50927 28322 50961 28390
rect 51000 28338 51023 28384
rect 50972 28322 51023 28328
rect 51029 28322 51063 28390
rect 51069 28338 51384 28384
rect 51069 28322 51384 28328
rect 51916 28322 51963 28369
rect 52242 28356 54774 28384
rect 54974 28356 55021 28369
rect 52208 28338 55021 28356
rect 54974 28328 55021 28338
rect 52208 28322 55021 28328
rect 50927 28289 51963 28322
rect 52006 28294 55021 28322
rect 51990 28289 55021 28294
rect 50927 28288 55021 28289
rect 41048 27823 47423 27857
rect 45714 26925 45748 27823
rect 48888 27516 48920 27938
rect 48926 27554 48958 27900
rect 50927 27483 50961 28288
rect 51029 28283 51063 28288
rect 51650 28282 51664 28288
rect 51864 28282 51928 28288
rect 51029 28267 51063 28276
rect 51636 28274 51650 28282
rect 51664 28274 51706 28282
rect 51166 28267 51786 28274
rect 51932 28267 52306 28288
rect 54718 28282 54986 28288
rect 51110 28261 54990 28267
rect 51110 28255 55014 28261
rect 55116 28255 55150 28390
rect 57752 28255 57786 28432
rect 57792 28352 58860 28362
rect 59110 28352 59222 28364
rect 57792 28349 59222 28352
rect 57792 28338 59207 28349
rect 57807 28290 57888 28337
rect 57935 28318 59207 28338
rect 57935 28317 58860 28318
rect 59110 28317 59207 28318
rect 57935 28316 59207 28317
rect 59259 28316 59293 28432
rect 57935 28312 59293 28316
rect 60518 28312 60574 28316
rect 61762 28312 61818 28316
rect 59110 28306 59207 28312
rect 57854 28268 57888 28290
rect 57907 28284 58804 28306
rect 59151 28271 59197 28306
rect 51106 28254 55150 28255
rect 51024 28240 51097 28242
rect 51110 28241 55150 28254
rect 50982 28193 51110 28240
rect 51122 28221 55150 28241
rect 57718 28221 57786 28255
rect 57807 28267 57888 28268
rect 57807 28255 57935 28267
rect 59098 28255 59109 28266
rect 57807 28221 59109 28255
rect 59123 28243 59225 28260
rect 51029 27625 51110 28193
rect 51166 27852 51786 28221
rect 51836 27904 51870 28221
rect 51931 28209 51932 28210
rect 51932 28208 51933 28209
rect 51944 28131 51978 28221
rect 51990 28209 51991 28210
rect 51989 28208 51990 28209
rect 52207 28146 52218 28157
rect 51891 28118 51991 28131
rect 51891 28084 52006 28118
rect 52031 28112 52218 28146
rect 52219 28084 52300 28131
rect 51932 28046 52006 28084
rect 52266 28046 52300 28084
rect 51932 28030 51990 28046
rect 51944 27904 51978 28030
rect 52207 28018 52218 28029
rect 52031 27984 52218 28018
rect 52368 27904 52402 28221
rect 54989 28209 54990 28210
rect 54990 28208 54991 28209
rect 51836 27870 52402 27904
rect 51084 27597 51101 27625
rect 51166 27608 51786 27798
rect 51944 27784 51978 27870
rect 51836 27750 52402 27784
rect 51836 27676 51870 27750
rect 51836 27638 51876 27676
rect 51944 27655 51978 27750
rect 52242 27704 52298 27728
rect 52214 27681 52298 27704
rect 52207 27680 52298 27681
rect 52207 27676 52218 27680
rect 52207 27672 52219 27676
rect 52207 27670 52298 27672
rect 52031 27655 52298 27670
rect 51891 27648 51991 27655
rect 51884 27642 51991 27648
rect 52031 27652 52300 27655
rect 51884 27638 52006 27642
rect 51826 27624 51834 27630
rect 51111 27597 51786 27608
rect 51836 27618 51870 27638
rect 51891 27618 52006 27638
rect 52031 27636 52218 27652
rect 52219 27618 52300 27652
rect 52368 27618 52402 27750
rect 51836 27608 52492 27618
rect 54990 27609 54991 27610
rect 54989 27608 54990 27609
rect 51836 27597 52592 27608
rect 55002 27597 55036 28221
rect 55116 27597 55150 28221
rect 57752 27597 57786 28221
rect 57838 28209 57935 28221
rect 57854 27722 57888 28209
rect 59110 28193 59191 28240
rect 59157 27707 59191 28193
rect 59110 27706 59191 27707
rect 59110 27694 59207 27706
rect 57807 27644 57888 27679
rect 57947 27660 59207 27694
rect 59110 27648 59207 27660
rect 57807 27632 57894 27644
rect 57848 27624 57894 27632
rect 59157 27625 59191 27648
rect 57854 27610 57894 27624
rect 59151 27613 59197 27624
rect 57807 27609 57894 27610
rect 57807 27603 57935 27609
rect 57807 27598 58764 27603
rect 57807 27597 57935 27598
rect 59098 27597 59109 27608
rect 51084 27563 59109 27597
rect 59123 27585 59225 27596
rect 51166 27483 51786 27563
rect 51836 27544 52492 27563
rect 51836 27530 51870 27544
rect 51836 27522 51876 27530
rect 51884 27528 51904 27530
rect 51836 27483 51870 27522
rect 51944 27483 51978 27544
rect 52207 27542 52218 27544
rect 52015 27529 52223 27542
rect 52031 27517 52218 27529
rect 52015 27508 52223 27517
rect 52368 27483 52402 27544
rect 55002 27483 55036 27563
rect 55116 27483 55150 27563
rect 57752 27483 57786 27563
rect 57823 27551 57935 27563
rect 59259 27483 59293 28312
rect 60518 28256 60574 28260
rect 61762 28256 61818 28260
rect 60518 27754 60574 27756
rect 61762 27754 61818 27756
rect 60518 27698 60574 27700
rect 61762 27698 61818 27700
rect 68713 27689 70426 31840
rect 72267 29782 72301 33090
rect 73078 32566 73112 33090
rect 73074 32532 73368 32566
rect 73078 32405 73112 32532
rect 73192 32511 73226 32532
rect 73058 32371 73112 32405
rect 73180 32383 73226 32511
rect 73192 32371 73226 32383
rect 73238 32371 73265 32382
rect 73080 32195 73146 32371
rect 73192 32195 73265 32371
rect 73078 32034 73112 32195
rect 73192 32183 73226 32195
rect 73180 32071 73226 32183
rect 73192 32034 73226 32071
rect 73334 32034 73368 32532
rect 73074 32000 73368 32034
rect 73784 32512 77408 33090
rect 77505 32512 77539 33090
rect 77619 32564 77653 33090
rect 78277 32564 78311 33090
rect 77619 32512 77664 32564
rect 73784 32454 78130 32512
rect 78277 32454 78322 32564
rect 73078 31950 73112 32000
rect 73042 31666 73386 31950
rect 73784 31666 78582 32454
rect 78820 31666 79661 33090
rect 80251 31666 80296 33090
rect 80909 32564 80943 33090
rect 80909 32502 80954 32564
rect 81023 32502 81057 33090
rect 82366 32658 82400 33090
rect 82366 32576 82456 32658
rect 81734 32532 82124 32566
rect 80468 31952 81292 32502
rect 81734 32034 81768 32532
rect 81863 32464 81995 32511
rect 81910 32430 81995 32464
rect 81837 32371 81893 32382
rect 81965 32371 82021 32382
rect 81848 32195 81893 32371
rect 81976 32195 82021 32371
rect 81863 32136 81995 32183
rect 81910 32102 81995 32136
rect 82090 32034 82124 32532
rect 81734 32000 82124 32034
rect 80502 31666 80714 31952
rect 80909 31666 80954 31952
rect 81023 31666 81057 31952
rect 81158 31866 81276 31952
rect 81720 31666 82142 31950
rect 82366 31666 82400 32576
rect 73042 31632 82412 31666
rect 73042 31611 73386 31632
rect 73784 31611 78582 31632
rect 78820 31611 79661 31632
rect 80251 31611 80296 31632
rect 80909 31611 80943 31632
rect 73042 31564 80534 31611
rect 80909 31564 80956 31611
rect 81023 31564 81057 31632
rect 81720 31564 82142 31632
rect 82366 31611 82400 31632
rect 82338 31564 82400 31611
rect 73042 31530 82400 31564
rect 73042 31330 73386 31530
rect 73108 30546 73350 30814
rect 73050 30424 73350 30546
rect 73108 30370 73350 30424
rect 50927 27449 59293 27483
rect 51166 27376 51786 27449
rect 51836 27428 51870 27449
rect 51944 27428 51978 27449
rect 52368 27428 52402 27449
rect 51836 27394 52402 27428
rect 51648 27210 51650 27274
rect 51676 27210 51706 27246
rect 55116 27010 55150 27449
rect 57752 27010 57786 27449
rect 60620 27090 60676 27098
rect 61760 27090 61816 27098
rect 60518 27034 60676 27042
rect 61760 27034 61818 27042
rect 41048 26891 46531 26925
rect 45714 26811 45748 26891
rect 45828 26811 45862 26891
rect 46336 26811 46347 26822
rect 45680 26777 46347 26811
rect 23298 25242 23972 25255
rect 22667 25221 23972 25242
rect 22682 25079 23302 25221
rect 23352 25187 23886 25206
rect 23386 25172 23884 25187
rect 23352 25147 23918 25153
rect 23352 25144 23386 25147
rect 23884 25144 23918 25147
rect 23318 25141 23420 25144
rect 23850 25141 23952 25144
rect 23318 25138 23952 25141
rect 23318 25107 23386 25138
rect 23509 25126 23761 25130
rect 23497 25107 23773 25126
rect 23850 25107 23952 25138
rect 22673 25040 23302 25079
rect 22600 24954 23302 25040
rect 22673 24802 23302 24954
rect 23352 25066 23386 25107
rect 23723 25092 23734 25095
rect 23531 25077 23739 25092
rect 23407 25066 23488 25077
rect 23531 25073 23816 25077
rect 23352 25024 23392 25066
rect 23400 25030 23488 25066
rect 23547 25058 23734 25073
rect 23735 25030 23816 25073
rect 23400 25024 23420 25030
rect 23352 24850 23386 25024
rect 23454 24992 23488 25030
rect 23782 24992 23816 25030
rect 23723 24964 23734 24975
rect 23547 24930 23734 24964
rect 23884 24850 23918 25107
rect 23352 24816 23918 24850
rect 22673 24748 22707 24802
rect 22673 24511 23302 24748
rect 22682 24326 23302 24511
rect 23352 24696 23918 24730
rect 23352 24483 23386 24696
rect 23723 24616 23734 24627
rect 23400 24489 23402 24576
rect 23407 24554 23488 24601
rect 23547 24582 23734 24616
rect 23735 24554 23816 24601
rect 23454 24500 23488 24554
rect 23782 24517 23816 24554
rect 23774 24508 23826 24517
rect 23776 24504 23822 24508
rect 23782 24500 23816 24504
rect 23536 24495 23734 24499
rect 23547 24483 23723 24488
rect 23746 24483 23854 24489
rect 23884 24483 23918 24696
rect 23318 24449 23952 24483
rect 23352 24374 23386 24449
rect 23884 24374 23918 24449
rect 23352 24340 23918 24374
rect 23180 23722 23380 23732
rect 23152 23694 23408 23704
rect 30760 21667 30973 25291
rect 31106 20312 31136 20320
rect 30942 20298 31014 20312
rect 31106 20298 31798 20312
rect 31106 20284 31108 20292
rect 30970 20270 31014 20284
rect 31106 20270 31770 20284
rect 22978 17516 24492 17530
rect 22712 17478 22736 17500
rect 22690 17454 22736 17478
rect 17612 16302 18792 16674
rect 29588 16596 30978 18890
rect 32368 16696 32402 26672
rect 45714 26153 45748 26777
rect 45828 26153 45862 26777
rect 45874 26765 45875 26766
rect 45873 26764 45874 26765
rect 46348 26749 46429 26796
rect 46395 26181 46429 26749
rect 45873 26165 45874 26166
rect 45874 26164 45875 26165
rect 46336 26153 46347 26164
rect 45680 26119 46347 26153
rect 45714 25495 45748 26119
rect 45828 25495 45862 26119
rect 45874 26107 45875 26108
rect 45873 26106 45874 26107
rect 46348 26091 46429 26138
rect 46395 25523 46429 26091
rect 45873 25507 45874 25508
rect 45874 25506 45875 25507
rect 46336 25495 46347 25506
rect 45680 25461 46347 25495
rect 45714 24837 45748 25461
rect 45828 24837 45862 25461
rect 45874 25449 45875 25450
rect 45873 25448 45874 25449
rect 46348 25433 46429 25480
rect 46395 24865 46429 25433
rect 45873 24849 45874 24850
rect 45874 24848 45875 24849
rect 46336 24837 46347 24848
rect 45680 24803 46347 24837
rect 45714 24179 45748 24803
rect 45828 24179 45862 24803
rect 45874 24791 45875 24792
rect 45873 24790 45874 24791
rect 46348 24775 46429 24822
rect 46395 24207 46429 24775
rect 45873 24191 45874 24192
rect 45874 24190 45875 24191
rect 46336 24179 46347 24190
rect 45680 24145 46347 24179
rect 45106 23536 45512 23914
rect 45026 23521 45512 23536
rect 45714 23521 45748 24145
rect 45828 23521 45862 24145
rect 45874 24133 45875 24134
rect 45873 24132 45874 24133
rect 46348 24117 46429 24164
rect 46395 23549 46429 24117
rect 45873 23533 45874 23534
rect 45874 23532 45875 23533
rect 46336 23521 46347 23532
rect 41048 23487 46347 23521
rect 45026 23466 45512 23487
rect 45106 23407 45512 23466
rect 45714 23407 45748 23487
rect 45828 23407 45862 23487
rect 46497 23407 46531 26891
rect 41048 23373 46531 23407
rect 51024 26208 55186 27010
rect 51024 26188 55204 26208
rect 57716 26194 59444 27010
rect 60628 26996 60676 27004
rect 61760 26996 61928 27024
rect 60620 26940 60676 26948
rect 61760 26940 61816 26968
rect 60676 26412 60684 26440
rect 60620 26356 60684 26384
rect 51024 23386 55186 26188
rect 59272 25572 59306 26140
rect 73078 25396 73112 29782
rect 73192 29227 73226 29782
rect 73784 29227 78582 31530
rect 78820 31524 79638 31530
rect 78820 29227 79661 31524
rect 80251 29227 80296 31530
rect 80909 29227 80943 31530
rect 73192 29180 80534 29227
rect 80909 29180 80956 29227
rect 81023 29180 81057 31530
rect 81720 31330 82142 31530
rect 82366 29227 82400 31530
rect 82338 29180 82400 29227
rect 73192 29112 73232 29180
rect 73242 29146 82400 29180
rect 73242 29140 73260 29146
rect 73192 29078 73226 29112
rect 73784 29090 78582 29146
rect 78820 29140 79638 29146
rect 73784 29078 78658 29090
rect 78820 29078 79661 29140
rect 80251 29078 80296 29146
rect 80909 29078 80943 29146
rect 81023 29078 81057 29146
rect 82366 29078 82400 29146
rect 73174 29044 82412 29078
rect 82418 29044 82434 29078
rect 73784 28558 78582 29044
rect 78624 28558 78658 29044
rect 73784 28524 78658 28558
rect 73784 28474 78582 28524
rect 73176 28424 73226 28458
rect 73784 28424 78672 28474
rect 78820 28424 79661 29044
rect 80251 28424 80296 29044
rect 80909 28424 80943 29044
rect 81023 28424 81057 29044
rect 82366 28424 82400 28458
rect 73114 28390 73166 28424
rect 73180 28390 82412 28424
rect 64946 24178 65342 24198
rect 64966 23869 64967 24178
rect 65322 23869 65342 24178
rect 64966 23868 65342 23869
rect 42158 22526 42184 22560
rect 42158 22438 42184 22472
rect 42192 22404 42218 22594
rect 45714 22154 45748 23373
rect 55022 23006 55186 23260
rect 54642 22566 55186 22988
rect 55192 22806 55206 23112
rect 55220 22806 55262 23112
rect 55276 22988 55440 23006
rect 55192 22636 55204 22806
rect 55276 22544 55440 22566
rect 47756 22152 47812 22162
rect 46108 22096 47812 22106
rect 50747 22022 55186 22193
rect 44964 20428 46384 20458
rect 46400 20436 46434 20475
rect 46502 20428 46536 21758
rect 51182 21160 55206 21165
rect 51216 21126 55240 21131
rect 73114 20464 73148 28390
rect 73180 28267 73202 28390
rect 73784 28369 78672 28390
rect 78820 28369 79661 28390
rect 80251 28369 80296 28390
rect 80909 28369 80943 28390
rect 73243 28322 80534 28369
rect 80909 28322 80956 28369
rect 81023 28322 81057 28390
rect 82366 28338 82412 28369
rect 82354 28322 82412 28338
rect 73290 28288 82412 28322
rect 73180 25495 73226 28267
rect 73238 28229 73273 28240
rect 73180 25483 73202 25495
rect 73228 25483 73273 28229
rect 73784 27908 78672 28288
rect 78820 28282 79638 28288
rect 78820 27920 79661 28282
rect 80251 27920 80296 28288
rect 80909 27920 80943 28288
rect 78820 27908 79633 27920
rect 79638 27908 79661 27920
rect 73784 27861 80534 27908
rect 80881 27861 80928 27908
rect 73784 27827 79612 27861
rect 79655 27827 80270 27861
rect 80313 27827 80928 27861
rect 73784 27759 78582 27827
rect 78820 27759 79612 27827
rect 81023 27759 81057 28288
rect 82354 28279 82390 28288
rect 82354 28241 82400 28279
rect 73784 27725 81057 27759
rect 81632 27776 82022 27810
rect 73784 27712 78582 27725
rect 76250 25822 76284 27712
rect 76286 26874 76331 27712
rect 77362 27062 78582 27712
rect 76286 25822 76320 26874
rect 76226 25788 78592 25822
rect 76226 25693 76284 25788
rect 76286 25693 76320 25788
rect 78397 25708 78408 25719
rect 76226 25646 76362 25693
rect 76421 25674 78408 25708
rect 78409 25646 78490 25693
rect 76226 25495 76284 25646
rect 76226 25483 76260 25495
rect 76286 25483 76320 25646
rect 76328 25483 76362 25646
rect 73216 25436 74728 25483
rect 75286 25436 76269 25483
rect 76286 25470 76362 25483
rect 76278 25436 76362 25470
rect 76536 25442 76630 25446
rect 76368 25436 76630 25442
rect 78456 25436 78490 25646
rect 78558 25436 78592 25788
rect 78820 25483 79612 27725
rect 81632 27278 81666 27776
rect 81846 27708 81893 27755
rect 81808 27674 81893 27708
rect 81735 27615 81780 27626
rect 81863 27615 81908 27626
rect 81746 27439 81780 27615
rect 81874 27439 81908 27615
rect 81846 27380 81893 27427
rect 81808 27346 81893 27380
rect 81988 27278 82022 27776
rect 81632 27244 82022 27278
rect 81614 26574 82036 27194
rect 82366 27186 82400 28241
rect 82402 28229 82434 28245
rect 82402 27186 82436 28229
rect 82480 27246 82514 33090
rect 82540 32564 82550 33090
rect 82540 31632 82570 32564
rect 82540 28460 82550 31632
rect 82576 29782 82610 33126
rect 84731 33090 93169 33126
rect 82728 31966 82730 32022
rect 82728 31710 82730 31766
rect 82728 31566 82730 31622
rect 82728 31310 82730 31366
rect 84731 31130 86164 33090
rect 97662 31810 97696 33126
rect 97764 33092 97798 33124
rect 98510 32580 101476 33126
rect 102022 32084 103672 33522
rect 104108 32082 105758 33520
rect 105836 33384 105852 33688
rect 105874 33198 105908 33766
rect 105914 33716 105968 33738
rect 105914 33688 105940 33710
rect 107056 33298 107060 33303
rect 107056 33112 107084 33298
rect 105836 33078 105852 33082
rect 97488 31804 99796 31810
rect 95538 31774 99796 31804
rect 95588 31622 95602 31724
rect 95616 31650 95658 31696
rect 97262 31656 97484 31676
rect 97300 31618 97446 31638
rect 84731 31113 91456 31130
rect 84731 31096 86164 31113
rect 84731 31062 91518 31096
rect 84731 30982 86164 31062
rect 86642 30982 91334 30993
rect 84731 30948 91334 30982
rect 84731 30489 86164 30948
rect 91335 30920 91463 30967
rect 87932 30662 88378 30768
rect 87796 30586 88378 30662
rect 87932 30526 88378 30586
rect 86738 30500 89058 30512
rect 91382 30502 91463 30920
rect 91335 30500 91463 30502
rect 86642 30489 91463 30500
rect 91484 30489 91518 31062
rect 84731 30455 91552 30489
rect 84731 30375 86164 30455
rect 86738 30375 86772 30455
rect 88882 30410 88929 30455
rect 86914 30409 88929 30410
rect 86898 30376 88929 30409
rect 87076 30375 87132 30376
rect 88626 30375 88682 30376
rect 89024 30375 89058 30455
rect 91335 30448 91463 30455
rect 91335 30443 91447 30448
rect 91264 30375 91376 30380
rect 91422 30375 91424 30380
rect 91484 30375 91518 30455
rect 97488 30408 99796 31774
rect 100066 30408 102374 31816
rect 102536 31288 102792 31290
rect 102564 31260 102764 31262
rect 97488 30390 102374 30408
rect 84731 30341 93037 30375
rect 97488 30372 99796 30390
rect 100066 30378 102374 30390
rect 84731 30330 86164 30341
rect 86738 30340 86772 30341
rect 86266 30336 86900 30340
rect 86266 30330 88898 30336
rect 88910 30330 88944 30333
rect 89024 30330 89058 30341
rect 91292 30330 91376 30341
rect 84731 30329 91376 30330
rect 84731 30324 87132 30329
rect 88626 30324 91376 30329
rect 84731 30318 91376 30324
rect 91422 30318 91480 30341
rect 84731 30307 91339 30318
rect 84731 30305 86164 30307
rect 82576 28460 82604 28478
rect 82540 28390 82604 28460
rect 82516 27748 82604 28390
rect 84006 27934 84040 29782
rect 85116 28894 86164 30305
rect 86738 30290 89098 30307
rect 86738 29666 86772 30290
rect 86852 29666 86886 30290
rect 88842 30284 88904 30290
rect 86898 30278 86899 30279
rect 86897 30277 86898 30278
rect 88870 30256 88904 30282
rect 88910 30240 88944 30290
rect 88950 30284 89098 30290
rect 89024 30282 89058 30284
rect 88950 30256 89070 30282
rect 89024 30240 89058 30256
rect 88908 30192 89058 30240
rect 88898 30122 89058 30192
rect 87942 29868 88388 30110
rect 88898 29890 88958 30122
rect 88062 29782 88302 29868
rect 87076 29714 87132 29728
rect 88772 29714 88828 29728
rect 86897 29678 86898 29679
rect 88898 29678 88899 29679
rect 88910 29678 88944 29890
rect 86898 29677 86899 29678
rect 87076 29666 87132 29672
rect 88372 29666 88992 29678
rect 89024 29666 89058 30122
rect 91484 29782 91518 30341
rect 97756 30188 97790 30372
rect 102414 30352 102666 30356
rect 102448 30318 102670 30322
rect 107056 30276 107060 33112
rect 97548 30154 98372 30188
rect 86738 29664 89058 29666
rect 86738 29632 89608 29664
rect 86738 29090 86772 29632
rect 86852 29280 86886 29632
rect 86898 29620 86899 29621
rect 86897 29619 86898 29620
rect 88372 29416 88992 29632
rect 87942 29398 88992 29416
rect 87686 29284 88992 29398
rect 86852 29090 86897 29280
rect 87942 29256 88992 29284
rect 89024 29630 89608 29632
rect 89024 29308 89076 29630
rect 89574 29616 89608 29630
rect 89414 29606 90454 29616
rect 89413 29550 89424 29561
rect 89097 29488 89178 29535
rect 89237 29516 89424 29550
rect 89425 29488 89506 29535
rect 89144 29450 89178 29488
rect 89472 29450 89506 29488
rect 89413 29422 89424 29433
rect 89237 29388 89424 29422
rect 89574 29308 89608 29606
rect 89024 29274 89608 29308
rect 90298 29340 91554 29376
rect 95442 29340 95476 29782
rect 90298 29306 95654 29340
rect 87942 29174 88388 29256
rect 86548 29056 86938 29090
rect 86548 29008 86582 29056
rect 86738 29022 86772 29056
rect 86690 29021 86772 29022
rect 86677 29008 86772 29021
rect 86852 29008 86886 29056
rect 86897 29020 86898 29021
rect 86898 29019 86899 29020
rect 86904 29008 86938 29056
rect 87024 29056 87414 29090
rect 87024 29008 87058 29056
rect 87166 29021 87272 29022
rect 87153 29008 87285 29021
rect 87380 29008 87414 29056
rect 88898 29020 88899 29021
rect 88897 29019 88898 29020
rect 88230 29008 88448 29019
rect 88778 29008 88828 29014
rect 88910 29008 88944 29256
rect 89024 29008 89058 29274
rect 90298 29008 91554 29306
rect 86548 28974 91554 29008
rect 86548 28902 86582 28974
rect 86693 28962 86796 28974
rect 86738 28954 86796 28962
rect 86852 28961 86886 28974
rect 86350 28894 86640 28902
rect 86662 28894 86696 28928
rect 86738 28894 86772 28954
rect 86840 28935 86890 28961
rect 86826 28934 86890 28935
rect 86818 28928 86826 28934
rect 86790 28907 86826 28928
rect 86790 28902 86830 28907
rect 86840 28902 86890 28934
rect 86904 28902 86938 28974
rect 87024 28902 87058 28974
rect 87076 28934 87132 28958
rect 87200 28954 87285 28974
rect 87138 28906 87172 28928
rect 87266 28906 87300 28928
rect 87127 28902 87172 28906
rect 86790 28894 86824 28902
rect 86826 28894 86890 28902
rect 86892 28895 87172 28902
rect 87255 28895 87300 28906
rect 86892 28894 87132 28895
rect 87138 28894 87172 28895
rect 87266 28894 87300 28895
rect 87380 28894 87414 28974
rect 88230 28908 88448 28928
rect 88910 28894 88944 28974
rect 89024 28894 89058 28974
rect 90298 28894 91554 28974
rect 85116 28860 91554 28894
rect 85116 28858 86164 28860
rect 86548 28858 86582 28860
rect 86738 28858 86772 28860
rect 86790 28858 86806 28860
rect 86814 28858 86824 28860
rect 86840 28858 86890 28860
rect 86904 28858 86938 28860
rect 87024 28858 87058 28860
rect 87138 28858 87172 28860
rect 87266 28858 87300 28860
rect 87380 28858 87414 28860
rect 89024 28858 89058 28860
rect 90298 28858 91554 28860
rect 85116 28824 91554 28858
rect 85322 28822 85356 28824
rect 85980 28822 86014 28824
rect 86094 28822 86128 28824
rect 86512 28822 89094 28824
rect 90334 28822 90368 28824
rect 90448 28822 90482 28824
rect 84790 28788 93138 28822
rect 83980 27884 84016 27922
rect 84790 27884 84824 28788
rect 85232 28714 85244 28772
rect 85260 28714 85272 28744
rect 85322 28708 85356 28788
rect 85980 28708 86014 28788
rect 86094 28708 86128 28788
rect 84854 28646 84926 28684
rect 84976 28674 86128 28708
rect 84892 28078 84926 28646
rect 85232 28608 85244 28668
rect 85260 28636 85272 28668
rect 85309 28662 85310 28663
rect 85310 28661 85311 28662
rect 85322 28502 85356 28674
rect 85368 28662 85369 28663
rect 85967 28662 85968 28663
rect 85367 28661 85368 28662
rect 85968 28661 85969 28662
rect 85980 28502 86014 28674
rect 86094 28502 86128 28674
rect 86512 28502 89094 28788
rect 90334 28708 90368 28788
rect 90448 28708 90482 28788
rect 92952 28708 92963 28719
rect 90334 28674 92963 28708
rect 90334 28502 90368 28674
rect 90448 28502 90482 28674
rect 90494 28662 90495 28663
rect 90493 28661 90494 28662
rect 92964 28646 93036 28684
rect 85116 28328 91554 28502
rect 92964 28366 92965 28367
rect 92963 28365 92964 28366
rect 93002 28328 93036 28646
rect 93104 28328 93138 28788
rect 85116 28294 93138 28328
rect 85116 28226 91554 28294
rect 93002 28226 93036 28294
rect 93104 28226 93138 28294
rect 95442 28226 95476 29306
rect 95478 29204 95510 29238
rect 95528 29166 95536 29296
rect 95544 29166 95578 29192
rect 95513 29154 95578 29166
rect 95506 28660 95578 29154
rect 95506 28629 95552 28660
rect 95506 28622 95540 28629
rect 95506 28608 95510 28622
rect 95506 28570 95552 28608
rect 95506 28378 95578 28570
rect 95588 28564 95602 28666
rect 95620 28638 95654 29306
rect 97548 28874 97582 30154
rect 97666 30102 97704 30144
rect 97628 30014 97654 30036
rect 97674 30018 97694 30102
rect 97708 30092 97746 30102
rect 97708 30070 97750 30092
rect 97756 30070 97790 30154
rect 102512 30138 103160 30140
rect 103170 30138 103818 30140
rect 103828 30138 104476 30140
rect 104486 30138 105134 30140
rect 105144 30138 105792 30140
rect 102512 30136 102670 30138
rect 102540 30110 103132 30112
rect 103198 30110 103790 30112
rect 103856 30110 104448 30112
rect 104514 30110 105106 30112
rect 105172 30110 105764 30112
rect 102540 30108 102698 30110
rect 97708 30046 97790 30070
rect 97686 30014 97688 30018
rect 97708 30014 97746 30046
rect 97628 30002 97726 30014
rect 97650 29064 97722 30002
rect 97650 29014 97726 29064
rect 97686 29010 97688 29014
rect 97674 28908 97694 29010
rect 97708 28982 97746 29014
rect 97756 28982 97790 30046
rect 101226 29920 101250 29974
rect 101342 29920 101364 29954
rect 101280 29886 101304 29920
rect 101318 29886 101828 29920
rect 101246 29824 101250 29858
rect 98806 29754 98892 29782
rect 98720 29738 98892 29754
rect 98720 29600 98874 29738
rect 101280 29604 101314 29886
rect 101318 29800 101368 29886
rect 101455 29806 101653 29817
rect 101318 29762 101454 29800
rect 101466 29772 101653 29806
rect 101654 29762 101764 29800
rect 101318 29712 101376 29762
rect 101382 29728 101454 29762
rect 101455 29718 101653 29729
rect 101692 29728 101764 29762
rect 101318 29604 101368 29712
rect 101466 29684 101653 29718
rect 101794 29604 101828 29886
rect 101280 29570 101304 29604
rect 101318 29570 101828 29604
rect 101878 29512 102172 29974
rect 102340 29512 102516 29974
rect 107056 29303 107060 30138
rect 108988 29516 108992 33303
rect 109512 31974 109760 31994
rect 109532 31783 109533 31974
rect 109740 31783 109760 31974
rect 109532 31782 109760 31783
rect 121259 29782 121293 34680
rect 124206 34657 127695 34982
rect 124386 32860 124390 34657
rect 124420 32928 124454 34657
rect 124522 34386 124556 34657
rect 125002 34370 125003 34371
rect 125001 34369 125002 34370
rect 125014 34358 125048 34657
rect 125059 34370 125060 34371
rect 125660 34370 125661 34371
rect 125060 34369 125061 34370
rect 125659 34369 125660 34370
rect 125672 34358 125706 34657
rect 125717 34370 125718 34371
rect 126318 34370 126319 34371
rect 125718 34369 125719 34370
rect 126317 34369 126318 34370
rect 126330 34358 126364 34657
rect 126375 34370 126376 34371
rect 126976 34370 126977 34371
rect 126376 34369 126377 34370
rect 126975 34369 126976 34370
rect 126988 34358 127022 34657
rect 127033 34370 127034 34371
rect 127634 34370 127635 34371
rect 127034 34369 127035 34370
rect 127633 34369 127634 34370
rect 127646 34358 127680 34657
rect 127760 34358 127794 34982
rect 129178 34750 129212 34982
rect 129283 34750 132804 34982
rect 133484 34892 133518 34904
rect 133262 34858 133518 34892
rect 133644 34892 133678 34904
rect 133960 34892 133994 34904
rect 133644 34858 133994 34892
rect 134390 34850 134424 35078
rect 134504 34850 134538 34884
rect 135162 34850 135196 34884
rect 135820 34850 135854 34884
rect 136318 34850 136352 35994
rect 136540 35992 137146 35994
rect 137198 35992 137804 35994
rect 136454 35960 136466 35992
rect 136524 35970 137146 35992
rect 136509 35960 137146 35970
rect 137182 35960 137804 35992
rect 136509 35958 137096 35960
rect 137908 35958 137942 36038
rect 142108 35958 142142 36038
rect 142222 35958 142256 36038
rect 144150 35958 144184 36038
rect 144264 36024 144298 36038
rect 144252 35982 144310 36024
rect 144264 35978 144298 35982
rect 144292 35970 144480 35978
rect 144292 35964 144492 35970
rect 144230 35958 144492 35964
rect 136386 35922 136394 35936
rect 136478 35926 142256 35958
rect 136478 35922 136488 35926
rect 136490 35922 136492 35926
rect 136504 35924 142256 35926
rect 144116 35924 144184 35958
rect 144226 35956 144492 35958
rect 144230 35944 144492 35956
rect 144288 35934 144492 35944
rect 144288 35924 144602 35934
rect 136524 35922 137096 35924
rect 136382 35908 136454 35922
rect 136472 35912 136488 35922
rect 136524 35912 136525 35913
rect 136382 35896 136460 35908
rect 136386 35868 136394 35896
rect 136374 35364 136394 35868
rect 136414 35840 136460 35896
rect 136402 35392 136454 35840
rect 136386 35288 136394 35364
rect 136414 35344 136460 35392
rect 136466 35344 136512 35912
rect 136523 35911 136524 35912
rect 136414 35328 136512 35344
rect 136414 35316 136454 35328
rect 136438 35312 136454 35316
rect 136466 35312 136512 35328
rect 136523 35312 136524 35313
rect 136386 35276 136394 35278
rect 136438 35276 136450 35312
rect 136478 35300 136512 35312
rect 136524 35311 136525 35312
rect 136936 35300 136970 35922
rect 137050 35346 137084 35922
rect 137125 35910 137170 35921
rect 137783 35910 137828 35921
rect 137050 35330 137084 35334
rect 137136 35330 137170 35910
rect 137794 35330 137828 35910
rect 137908 35330 137942 35924
rect 142095 35912 142096 35913
rect 142096 35911 142097 35912
rect 138120 35330 138160 35338
rect 138176 35330 138188 35366
rect 142108 35346 142142 35924
rect 142108 35330 142142 35334
rect 137078 35304 142114 35330
rect 137074 35300 142118 35304
rect 142222 35300 142256 35924
rect 144150 35842 144184 35924
rect 144310 35912 144602 35924
rect 144326 35910 144602 35912
rect 144530 35842 144564 35896
rect 144632 35842 144666 36038
rect 144150 35808 144974 35842
rect 144530 35348 144564 35808
rect 144632 35348 144666 35808
rect 147416 35602 147418 36990
rect 147392 35396 147418 35602
rect 147416 35390 147418 35396
rect 147742 36122 153662 38864
rect 154131 36122 154165 40420
rect 154245 40383 154292 40399
rect 154233 40318 154292 40383
rect 154903 40368 154950 40399
rect 155561 40368 155608 40399
rect 156219 40368 156266 40399
rect 154891 40352 154950 40368
rect 155549 40352 155608 40368
rect 156207 40352 156266 40368
rect 154342 40318 154950 40352
rect 155000 40318 155608 40352
rect 155658 40318 156266 40352
rect 154233 40309 154268 40318
rect 154891 40309 154926 40318
rect 155549 40309 155584 40318
rect 156207 40309 156242 40318
rect 154233 40271 154279 40309
rect 154184 36230 154210 36346
rect 154212 36271 154238 36318
rect 154245 36271 154279 40271
rect 154280 40270 154313 40275
rect 154891 40271 154937 40309
rect 154280 37906 154314 40270
rect 154280 36283 154325 37906
rect 154334 36274 154338 36486
rect 154362 36271 154366 36514
rect 154903 36271 154937 40271
rect 154938 40270 154971 40275
rect 155549 40271 155595 40309
rect 154938 37906 154972 40270
rect 155561 39228 155595 40271
rect 155527 38560 155538 39228
rect 155555 38560 155595 39228
rect 154938 36283 154983 37906
rect 155561 37372 155595 38560
rect 155527 36306 155538 37372
rect 155555 36306 155595 37372
rect 155561 36271 155595 36306
rect 155596 40270 155629 40275
rect 156207 40271 156253 40309
rect 155596 37906 155630 40270
rect 156185 38560 156188 39228
rect 156213 38560 156216 39228
rect 155596 36283 155641 37906
rect 155654 36276 155664 36484
rect 155682 36271 155692 36512
rect 156185 36271 156188 37372
rect 156213 36271 156216 37372
rect 156219 36271 156253 40271
rect 156254 40270 156287 40275
rect 156254 37906 156288 40270
rect 156254 36283 156299 37906
rect 154212 36230 154292 36271
rect 154233 36190 154292 36230
rect 154295 36224 154950 36271
rect 154953 36224 155608 36271
rect 155611 36224 156266 36271
rect 154233 36174 154268 36190
rect 154233 36159 154248 36174
rect 154302 36156 154320 36224
rect 154330 36190 154950 36224
rect 155000 36190 155608 36224
rect 154330 36184 154348 36190
rect 154891 36174 154926 36190
rect 155549 36174 155584 36190
rect 155618 36156 155628 36224
rect 155646 36184 155656 36224
rect 155658 36190 156266 36224
rect 156207 36174 156242 36190
rect 154245 36122 154279 36156
rect 154903 36122 154937 36156
rect 155561 36122 155595 36156
rect 156219 36122 156253 36156
rect 156368 36122 156402 40420
rect 147742 36091 156402 36122
rect 156877 36091 156911 40761
rect 157017 36091 157051 40761
rect 157131 37906 157165 40761
rect 157350 38618 157352 38774
rect 157535 37906 157569 40761
rect 157131 36091 157176 37906
rect 157535 36091 157580 37906
rect 157649 36091 157683 40761
rect 159067 39248 159082 39330
rect 158360 39204 158750 39238
rect 159105 39210 159120 39368
rect 157686 38560 157696 38756
rect 158360 38706 158394 39204
rect 158447 39043 158481 39204
rect 158574 39136 158621 39183
rect 158536 39102 158621 39136
rect 158493 39043 158508 39054
rect 158591 39043 158636 39054
rect 158447 38867 158508 39043
rect 158602 38867 158636 39043
rect 158447 38844 158481 38867
rect 158447 38706 158487 38844
rect 158496 38720 158515 38816
rect 158574 38808 158621 38855
rect 158536 38774 158621 38808
rect 158716 38706 158750 39204
rect 157742 38560 157752 38700
rect 158360 38672 158750 38706
rect 158346 38002 158768 38622
rect 159071 38560 159098 38712
rect 159099 38560 159126 38740
rect 158348 37030 158354 37286
rect 158376 37058 158382 37258
rect 147742 36088 157683 36091
rect 147742 35748 153662 36088
rect 154131 35995 154165 36088
rect 154213 36057 157683 36088
rect 147742 35528 153672 35748
rect 144452 35334 144844 35348
rect 144388 35322 144844 35334
rect 144452 35306 144844 35322
rect 145518 35312 146064 35348
rect 146614 35318 146940 35348
rect 147276 35318 147606 35348
rect 136478 35296 142176 35300
rect 136382 35238 136454 35276
rect 136478 35266 142118 35296
rect 142188 35266 142256 35300
rect 144360 35300 144844 35306
rect 144360 35294 144492 35300
rect 144632 35292 144666 35300
rect 136478 35254 136512 35266
rect 136524 35254 136525 35255
rect 136386 35216 136394 35238
rect 136368 34854 136394 35216
rect 136414 35218 136454 35238
rect 136466 35218 136512 35254
rect 136523 35253 136524 35254
rect 136414 35188 136523 35218
rect 136396 34854 136523 35188
rect 136936 35194 136970 35266
rect 137096 35262 142118 35266
rect 137096 35254 142096 35262
rect 137136 35218 137170 35254
rect 137794 35218 137828 35254
rect 137136 35194 137181 35218
rect 137794 35194 137839 35218
rect 137908 35194 137942 35254
rect 138120 35230 138160 35254
rect 138176 35240 138188 35254
rect 142222 35194 142256 35266
rect 144452 35244 144900 35292
rect 145490 35284 146092 35292
rect 146586 35290 146940 35292
rect 147276 35290 147634 35292
rect 136936 35160 142256 35194
rect 136368 34850 136523 34854
rect 137136 34850 137181 35160
rect 137794 34850 137839 35160
rect 137908 34850 137942 35160
rect 133412 34816 143664 34850
rect 129178 34716 132804 34750
rect 124484 34296 124556 34334
rect 124606 34324 127794 34358
rect 125001 34312 125002 34313
rect 125002 34311 125003 34312
rect 124522 33728 124556 34296
rect 125002 33712 125003 33713
rect 125001 33711 125002 33712
rect 125014 33700 125048 34324
rect 125060 34312 125061 34313
rect 125659 34312 125660 34313
rect 125059 34311 125060 34312
rect 125660 34311 125661 34312
rect 125059 33712 125060 33713
rect 125660 33712 125661 33713
rect 125060 33711 125061 33712
rect 125659 33711 125660 33712
rect 125672 33700 125706 34324
rect 125718 34312 125719 34313
rect 126317 34312 126318 34313
rect 125717 34311 125718 34312
rect 126318 34311 126319 34312
rect 125717 33712 125718 33713
rect 126318 33712 126319 33713
rect 125718 33711 125719 33712
rect 126317 33711 126318 33712
rect 126330 33700 126364 34324
rect 126376 34312 126377 34313
rect 126975 34312 126976 34313
rect 126375 34311 126376 34312
rect 126976 34311 126977 34312
rect 126375 33712 126376 33713
rect 126976 33712 126977 33713
rect 126376 33711 126377 33712
rect 126975 33711 126976 33712
rect 126988 33700 127022 34324
rect 127034 34312 127035 34313
rect 127633 34312 127634 34313
rect 127033 34311 127034 34312
rect 127634 34311 127635 34312
rect 127033 33712 127034 33713
rect 127634 33712 127635 33713
rect 127034 33711 127035 33712
rect 127633 33711 127634 33712
rect 127646 33700 127680 34324
rect 127760 33700 127794 34324
rect 124484 33638 124556 33676
rect 124606 33666 127794 33700
rect 125001 33654 125002 33655
rect 125002 33653 125003 33654
rect 124522 33070 124556 33638
rect 125002 33054 125003 33055
rect 125001 33053 125002 33054
rect 125014 33042 125048 33666
rect 125060 33654 125061 33655
rect 125659 33654 125660 33655
rect 125059 33653 125060 33654
rect 125660 33653 125661 33654
rect 125059 33054 125060 33055
rect 125660 33054 125661 33055
rect 125060 33053 125061 33054
rect 125659 33053 125660 33054
rect 125672 33042 125706 33666
rect 125718 33654 125719 33655
rect 126317 33654 126318 33655
rect 125717 33653 125718 33654
rect 126318 33653 126319 33654
rect 125717 33054 125718 33055
rect 126318 33054 126319 33055
rect 125718 33053 125719 33054
rect 126317 33053 126318 33054
rect 126330 33042 126364 33666
rect 126376 33654 126377 33655
rect 126975 33654 126976 33655
rect 126375 33653 126376 33654
rect 126976 33653 126977 33654
rect 126375 33054 126376 33055
rect 126976 33054 126977 33055
rect 126376 33053 126377 33054
rect 126975 33053 126976 33054
rect 126988 33042 127022 33666
rect 127034 33654 127035 33655
rect 127633 33654 127634 33655
rect 127033 33653 127034 33654
rect 127634 33653 127635 33654
rect 127033 33054 127034 33055
rect 127634 33054 127635 33055
rect 127034 33053 127035 33054
rect 127633 33053 127634 33054
rect 127646 33042 127680 33666
rect 127760 33042 127794 33666
rect 124606 33008 127794 33042
rect 125014 32928 125048 33008
rect 125672 32928 125706 33008
rect 126330 32928 126364 33008
rect 126988 32928 127022 33008
rect 127646 32928 127680 33008
rect 127760 32928 127794 33008
rect 129283 32928 132804 34716
rect 134390 34736 134424 34816
rect 134504 34736 134538 34816
rect 135162 34736 135196 34816
rect 135444 34736 135808 34747
rect 135820 34736 135854 34816
rect 136318 34747 136352 34816
rect 135866 34736 136356 34747
rect 136368 34742 136394 34816
rect 136396 34802 136523 34816
rect 137136 34802 137181 34816
rect 137794 34802 137839 34816
rect 136396 34748 136454 34802
rect 136466 34748 136512 34802
rect 136396 34742 136512 34748
rect 136404 34740 136512 34742
rect 136382 34736 136512 34740
rect 137136 34736 137170 34802
rect 137794 34736 137828 34802
rect 137908 34736 137942 34816
rect 143630 34760 143664 34816
rect 143478 34736 143489 34747
rect 143490 34740 143664 34760
rect 134390 34702 143489 34736
rect 134390 34278 134424 34702
rect 134504 34278 134538 34702
rect 134550 34690 134551 34691
rect 135149 34690 135150 34691
rect 134549 34689 134550 34690
rect 135150 34689 135151 34690
rect 134549 34290 134550 34291
rect 135150 34290 135151 34291
rect 134550 34289 134551 34290
rect 135149 34289 135150 34290
rect 135162 34278 135196 34702
rect 135208 34690 135209 34691
rect 135807 34690 135808 34691
rect 135820 34690 135854 34702
rect 135866 34690 135867 34691
rect 135207 34689 135208 34690
rect 135808 34689 135809 34690
rect 135820 34689 135866 34690
rect 135820 34291 135865 34689
rect 135207 34290 135208 34291
rect 135808 34290 135809 34291
rect 135820 34290 135866 34291
rect 135208 34289 135209 34290
rect 135807 34289 135808 34290
rect 135256 34278 135808 34289
rect 135820 34278 135854 34290
rect 135866 34289 135867 34290
rect 136318 34289 136352 34702
rect 136386 34630 136394 34696
rect 136404 34690 136512 34702
rect 136414 34658 136454 34690
rect 136438 34654 136454 34658
rect 136438 34618 136450 34654
rect 136478 34642 136512 34690
rect 137136 34642 137170 34702
rect 137794 34642 137828 34702
rect 137908 34642 137942 34702
rect 143490 34674 143562 34712
rect 143528 34654 143562 34674
rect 143490 34642 143578 34654
rect 143630 34642 143664 34740
rect 136382 34580 136454 34618
rect 136420 34362 136454 34580
rect 135866 34278 136356 34289
rect 136380 34284 136394 34362
rect 136408 34290 136454 34362
rect 136478 34608 143578 34642
rect 143596 34608 143664 34642
rect 136478 34290 136512 34608
rect 136404 34282 136512 34290
rect 136382 34278 136512 34282
rect 137136 34278 137170 34608
rect 137794 34278 137828 34608
rect 137908 34278 137942 34608
rect 143490 34596 143578 34608
rect 143528 34306 143562 34596
rect 143478 34278 143489 34289
rect 134390 34244 143489 34278
rect 134390 34164 134424 34244
rect 134504 34164 134538 34244
rect 135162 34164 135196 34244
rect 135820 34164 135854 34244
rect 136318 34164 136352 34244
rect 136380 34168 136394 34238
rect 136404 34232 136512 34244
rect 136408 34194 136454 34232
rect 136466 34194 136512 34232
rect 137136 34194 137170 34244
rect 137794 34194 137828 34244
rect 136408 34168 136523 34194
rect 136380 34164 136523 34168
rect 137136 34164 137181 34194
rect 137794 34164 137839 34194
rect 137908 34164 137942 34244
rect 143630 34164 143664 34608
rect 133412 34130 143664 34164
rect 124420 32894 132804 32928
rect 108802 29174 108878 29426
rect 108882 29234 108938 29486
rect 108966 29308 108992 29516
rect 108988 29303 108992 29308
rect 106212 29084 106295 29161
rect 108802 29090 108880 29174
rect 108882 29090 108940 29234
rect 97708 28958 97790 28982
rect 97708 28936 97750 28958
rect 97708 28926 97746 28936
rect 97686 28907 97688 28908
rect 97756 28907 97790 28958
rect 119458 29056 119848 29090
rect 97603 28874 98504 28907
rect 97548 28840 98504 28874
rect 97603 28804 98504 28840
rect 98702 28804 99694 28907
rect 97603 28769 97826 28804
rect 97603 28757 97844 28769
rect 99806 28757 99812 28806
rect 99834 28757 99868 28862
rect 100012 28757 101004 28907
rect 101180 28757 102172 28907
rect 97603 28723 102172 28757
rect 97603 28711 97844 28723
rect 97603 28644 97826 28711
rect 97892 28644 98144 28723
rect 98910 28717 99460 28723
rect 98938 28689 99432 28704
rect 95616 28592 95658 28638
rect 95513 28366 95578 28378
rect 95478 28294 95510 28328
rect 95528 28278 95536 28366
rect 95544 28340 95578 28366
rect 95620 28226 95654 28592
rect 85116 28192 95654 28226
rect 97603 28372 98176 28644
rect 99806 28562 99812 28723
rect 99834 28590 99868 28723
rect 85116 28094 91554 28192
rect 85116 28072 92388 28094
rect 85116 28050 91554 28072
rect 84854 27988 84926 28026
rect 84976 28016 91554 28050
rect 84892 27884 84926 27988
rect 84963 27922 84964 27923
rect 84964 27921 84965 27922
rect 85116 27884 91554 28016
rect 83942 27850 83978 27884
rect 83980 27850 84636 27884
rect 84790 27882 91554 27884
rect 93104 27882 93138 28192
rect 95442 27882 95476 28192
rect 97603 28111 97826 28372
rect 100012 28212 101004 28723
rect 101180 28220 102172 28723
rect 97603 28099 97844 28111
rect 102340 28099 105964 28907
rect 97603 28065 105964 28099
rect 97603 28060 97844 28065
rect 95517 28053 97844 28060
rect 95517 28049 97826 28053
rect 95528 28037 97826 28049
rect 95517 28026 97826 28037
rect 95544 27882 95578 28026
rect 97603 27957 97826 28026
rect 101496 28002 101862 28016
rect 101468 27974 101890 27988
rect 95617 27946 96984 27957
rect 97506 27946 97826 27957
rect 95628 27912 97826 27946
rect 84790 27850 97062 27882
rect 83980 27812 84016 27850
rect 84790 27782 84824 27850
rect 84892 27782 84926 27850
rect 85116 27848 97062 27850
rect 85116 27834 91560 27848
rect 85116 27782 91554 27834
rect 82672 27768 91554 27782
rect 92964 27768 93067 27780
rect 93104 27768 93138 27848
rect 95442 27768 95476 27848
rect 95513 27779 95616 27780
rect 95513 27772 96374 27779
rect 95506 27768 96374 27772
rect 96876 27768 96887 27779
rect 82672 27765 93067 27768
rect 82672 27748 93052 27765
rect 82516 27712 82586 27748
rect 82516 27246 82550 27712
rect 82574 27246 82584 27712
rect 82472 27186 82612 27246
rect 82276 27100 82612 27186
rect 82276 26798 82552 27100
rect 82574 26874 82584 27100
rect 82366 25495 82400 26798
rect 82368 25483 82400 25495
rect 78702 25436 80534 25483
rect 82338 25479 82400 25483
rect 82338 25436 82385 25479
rect 82402 25457 82436 26798
rect 82402 25445 82434 25457
rect 73238 25402 76269 25436
rect 76286 25402 76294 25436
rect 76296 25402 82385 25436
rect 73238 25386 73274 25402
rect 76224 25396 76260 25402
rect 76226 25334 76260 25396
rect 76286 25334 76362 25402
rect 76368 25396 76630 25402
rect 76368 25368 76630 25390
rect 76480 25340 76630 25368
rect 78456 25347 78490 25402
rect 78409 25334 78490 25347
rect 78558 25334 78592 25402
rect 78820 25334 79612 25402
rect 82480 25334 82514 26798
rect 73174 25300 73182 25334
rect 73216 25300 82448 25334
rect 82482 25300 82514 25334
rect 76226 24680 76260 25300
rect 76286 24680 76362 25300
rect 78456 24693 78490 25300
rect 78409 24680 78490 24693
rect 78558 24680 78592 25300
rect 78820 24680 79612 25300
rect 73216 24646 82448 24680
rect 73228 24625 73262 24646
rect 76226 24625 76260 24646
rect 73228 24578 74546 24625
rect 75286 24584 76260 24625
rect 76286 24612 76362 24646
rect 75286 24578 76270 24584
rect 73228 24510 73268 24578
rect 73278 24544 76270 24578
rect 73278 24538 73296 24544
rect 76224 24538 76270 24544
rect 76280 24578 76362 24612
rect 78456 24578 78490 24646
rect 78558 24578 78592 24646
rect 78820 24625 79612 24646
rect 82402 24625 82436 24646
rect 78702 24578 80534 24625
rect 82374 24584 82436 24625
rect 82368 24578 82436 24584
rect 76280 24544 82436 24578
rect 73228 22241 73262 24510
rect 76226 23536 76260 24538
rect 76280 24510 76362 24544
rect 76286 23678 76362 24510
rect 78456 23678 78490 24544
rect 76286 23662 76354 23678
rect 76286 23536 76320 23662
rect 78397 23650 78408 23661
rect 76421 23616 78408 23650
rect 78558 23536 78592 24544
rect 76226 23502 78592 23536
rect 76286 22241 76320 23502
rect 78820 23442 79612 24544
rect 82368 24538 82386 24544
rect 82396 24510 82436 24544
rect 79344 22241 79378 23442
rect 82402 22241 82436 24510
rect 73228 22194 74546 22241
rect 76258 22228 76320 22241
rect 79316 22228 79378 22241
rect 76258 22200 76326 22228
rect 79316 22200 79384 22228
rect 76252 22194 76326 22200
rect 76336 22194 76354 22200
rect 79310 22194 79384 22200
rect 79394 22194 79412 22200
rect 79628 22194 80542 22241
rect 82374 22200 82436 22241
rect 82368 22194 82436 22200
rect 73228 22126 73268 22194
rect 73278 22160 76326 22194
rect 76332 22160 79384 22194
rect 79390 22160 82436 22194
rect 73278 22154 73296 22160
rect 76252 22154 76270 22160
rect 76280 22126 76326 22160
rect 76336 22154 76354 22160
rect 79310 22154 79328 22160
rect 79338 22126 79384 22160
rect 79394 22154 79412 22160
rect 82368 22154 82386 22160
rect 82396 22126 82436 22160
rect 73228 22092 73262 22126
rect 76286 22092 76320 22126
rect 79344 22092 79378 22126
rect 82402 22092 82436 22126
rect 73210 22058 82470 22092
rect 82516 20464 82550 26798
rect 84790 25366 84824 27748
rect 85116 27734 93052 27748
rect 93070 27734 93138 27768
rect 95408 27734 96887 27768
rect 84908 27436 84932 27454
rect 84886 27408 84932 27436
rect 85116 27392 91554 27734
rect 92964 27722 93052 27734
rect 93002 27420 93036 27722
rect 92952 27392 92963 27403
rect 85116 27358 92963 27392
rect 85116 27310 91554 27358
rect 92964 27330 93036 27368
rect 93002 27322 93036 27330
rect 92964 27310 93052 27322
rect 93104 27310 93138 27734
rect 95442 27310 95476 27734
rect 95528 27722 95616 27734
rect 95544 27322 95616 27722
rect 96888 27706 96960 27744
rect 96926 27338 96960 27706
rect 95528 27321 95616 27322
rect 95528 27314 96374 27321
rect 95506 27310 96374 27314
rect 96876 27310 96887 27321
rect 85116 27294 93052 27310
rect 93070 27294 93138 27310
rect 85116 27276 93138 27294
rect 95408 27276 96887 27310
rect 85116 27270 93102 27276
rect 85116 27266 91554 27270
rect 92964 27266 93067 27270
rect 85116 27264 93074 27266
rect 85116 27242 92996 27264
rect 93042 27242 93074 27264
rect 85116 27196 91554 27242
rect 93104 27196 93138 27276
rect 95442 27196 95476 27276
rect 95513 27264 95616 27276
rect 97028 27196 97062 27848
rect 85116 27162 97062 27196
rect 97603 27453 97826 27912
rect 97603 27395 97844 27453
rect 85116 26076 91554 27162
rect 85116 26042 92952 26076
rect 85116 25234 91554 26042
rect 93104 25366 93138 27162
rect 85532 25224 85634 25226
rect 85532 25196 85606 25198
rect 85276 25080 86422 25140
rect 85116 24722 85516 24758
rect 85566 24722 85600 24754
rect 85761 24722 85937 24756
rect 86098 24722 86132 24754
rect 85116 24688 91422 24722
rect 85116 24544 85516 24688
rect 85566 24614 85606 24688
rect 85614 24614 85634 24688
rect 85668 24620 85702 24646
rect 85996 24620 86030 24646
rect 85566 24608 85600 24614
rect 85637 24608 85749 24620
rect 85949 24608 86061 24620
rect 86098 24608 86132 24688
rect 86142 24620 86224 24646
rect 85566 24582 86262 24608
rect 85566 24574 86132 24582
rect 85566 24544 85600 24574
rect 85116 24522 85606 24544
rect 85116 24520 85548 24522
rect 85116 24516 85516 24520
rect 85566 24516 85600 24522
rect 85116 24494 85634 24516
rect 86098 24494 86132 24574
rect 90580 24568 90836 24570
rect 90608 24540 90808 24542
rect 85116 24492 86132 24494
rect 85116 24446 85516 24492
rect 85566 24460 86132 24492
rect 85116 23970 85516 24392
rect 85566 24340 86132 24374
rect 85566 24018 85600 24340
rect 85937 24260 85948 24271
rect 85621 24198 85702 24245
rect 85761 24226 85948 24260
rect 85949 24198 86030 24245
rect 85668 24160 85702 24198
rect 85996 24160 86030 24198
rect 85937 24132 85948 24143
rect 85610 24096 85682 24102
rect 85761 24098 85948 24132
rect 85626 24040 85682 24046
rect 86098 24018 86132 24340
rect 85566 23984 86132 24018
rect 85152 23595 85186 23970
rect 85254 23962 85296 23970
rect 85279 23924 85296 23962
rect 86164 23898 86798 23908
rect 91484 23595 91518 24626
rect 84763 23561 92937 23595
rect 85152 23481 85186 23561
rect 85118 23447 85186 23481
rect 85207 23481 85335 23493
rect 91335 23481 91447 23493
rect 91484 23481 91518 23561
rect 85207 23478 91447 23481
rect 85207 23447 91432 23478
rect 91450 23447 91518 23481
rect 85152 22823 85186 23447
rect 85238 23435 85335 23447
rect 91335 23435 91432 23447
rect 85192 23406 85248 23420
rect 85254 23320 85288 23435
rect 91382 23320 91416 23435
rect 91323 23292 91334 23303
rect 85207 23230 85288 23277
rect 85347 23258 91334 23292
rect 91335 23230 91416 23277
rect 85254 22836 85288 23230
rect 91382 22836 91416 23230
rect 91424 22916 91480 22922
rect 91424 22860 91478 22866
rect 85118 22789 85186 22823
rect 85207 22835 85288 22836
rect 91335 22835 91416 22836
rect 85207 22823 85335 22835
rect 91335 22823 91432 22835
rect 91484 22823 91518 23447
rect 85207 22789 91432 22823
rect 91450 22789 91518 22823
rect 85152 22520 85186 22789
rect 85238 22777 85335 22789
rect 91335 22777 91432 22789
rect 85254 22662 85288 22777
rect 91382 22662 91416 22777
rect 91424 22682 91480 22706
rect 91323 22634 91334 22645
rect 85347 22600 91334 22634
rect 91484 22520 91518 22789
rect 85152 22486 91518 22520
rect 85192 22202 86280 22206
rect 84862 22131 92838 22165
rect 86280 22066 86916 22072
rect 86224 22010 86972 22044
rect 95442 21778 95476 27162
rect 95544 25460 95578 27162
rect 97603 26795 97826 27395
rect 97603 26737 97844 26795
rect 97603 26137 97826 26737
rect 102340 26624 105964 28065
rect 105971 26660 105982 28837
rect 108881 28614 108886 28878
rect 108881 28518 108892 28614
rect 119458 28558 119492 29056
rect 119672 28988 119719 29035
rect 119634 28954 119719 28988
rect 119561 28895 119606 28906
rect 119689 28895 119734 28906
rect 119572 28719 119606 28895
rect 119700 28719 119734 28895
rect 119672 28660 119719 28707
rect 119634 28626 119719 28660
rect 119814 28558 119848 29056
rect 119458 28524 119848 28558
rect 119934 29056 120324 29090
rect 119934 29028 119968 29056
rect 119934 28620 120002 29028
rect 120148 28988 120195 29035
rect 120110 28954 120195 28988
rect 120037 28895 120082 28906
rect 120165 28895 120210 28906
rect 120048 28719 120082 28895
rect 120176 28719 120210 28895
rect 120148 28660 120195 28707
rect 120110 28626 120195 28660
rect 119934 28558 119968 28620
rect 120290 28558 120324 29056
rect 119934 28524 120324 28558
rect 108922 27886 109032 28454
rect 110006 28234 110304 28250
rect 110022 27994 110304 28234
rect 119440 27861 119862 28474
rect 119347 27827 119915 27861
rect 119916 27854 120338 28474
rect 121824 28154 121840 29668
rect 122576 27904 122609 31554
rect 122610 27870 122643 31520
rect 127760 31411 127794 32894
rect 129283 32858 132804 32894
rect 124389 31375 127830 31411
rect 129319 31375 129353 32858
rect 133080 32022 133130 32028
rect 133136 32022 133158 32056
rect 133080 31828 133130 31836
rect 133136 31800 133158 31836
rect 129433 31375 129467 31409
rect 130091 31375 130125 31409
rect 130749 31375 130783 31409
rect 131407 31375 131441 31409
rect 132065 31375 132099 31409
rect 132723 31375 132729 31409
rect 124389 31341 132769 31375
rect 124389 27964 127830 31341
rect 129319 31261 129353 31341
rect 129433 31261 129467 31341
rect 130091 31261 130125 31341
rect 130749 31261 130783 31341
rect 131407 31261 131441 31341
rect 132065 31261 132099 31341
rect 132757 31313 132769 31341
rect 132723 31279 132769 31313
rect 132596 31261 132607 31272
rect 129319 31227 132607 31261
rect 129319 30603 129353 31227
rect 129433 30603 129467 31227
rect 129479 31215 129480 31216
rect 130078 31215 130079 31216
rect 129478 31214 129479 31215
rect 130079 31214 130080 31215
rect 129478 30615 129479 30616
rect 130079 30615 130080 30616
rect 129479 30614 129480 30615
rect 130078 30614 130079 30615
rect 130091 30603 130125 31227
rect 130137 31215 130138 31216
rect 130736 31215 130737 31216
rect 130136 31214 130137 31215
rect 130737 31214 130738 31215
rect 130136 30615 130137 30616
rect 130737 30615 130738 30616
rect 130137 30614 130138 30615
rect 130736 30614 130737 30615
rect 130749 30603 130783 31227
rect 130795 31215 130796 31216
rect 131394 31215 131395 31216
rect 130794 31214 130795 31215
rect 131395 31214 131396 31215
rect 130794 30615 130795 30616
rect 131395 30615 131396 30616
rect 130795 30614 130796 30615
rect 131394 30614 131395 30615
rect 131407 30603 131441 31227
rect 131453 31215 131454 31216
rect 132052 31215 132053 31216
rect 131452 31214 131453 31215
rect 132053 31214 132054 31215
rect 131452 30615 131453 30616
rect 132053 30615 132054 30616
rect 131453 30614 131454 30615
rect 132052 30614 132053 30615
rect 132065 30603 132099 31227
rect 132111 31215 132112 31216
rect 132110 31214 132111 31215
rect 132608 31211 132689 31246
rect 132717 31237 132723 31239
rect 132608 31199 132695 31211
rect 132621 31144 132640 31199
rect 132649 31144 132695 31199
rect 132717 31172 132727 31237
rect 132655 30696 132702 31144
rect 132110 30615 132111 30616
rect 132111 30614 132112 30615
rect 132596 30603 132607 30614
rect 129319 30569 132607 30603
rect 132621 30591 132640 30696
rect 132649 30631 132695 30696
rect 132649 30619 132668 30631
rect 132689 30619 132695 30631
rect 132717 30668 132730 31172
rect 132717 30593 132727 30668
rect 132717 30591 132723 30593
rect 129319 29945 129353 30569
rect 129433 29945 129467 30569
rect 129479 30557 129480 30558
rect 130078 30557 130079 30558
rect 129478 30556 129479 30557
rect 130079 30556 130080 30557
rect 129478 29957 129479 29958
rect 130079 29957 130080 29958
rect 129479 29956 129480 29957
rect 130078 29956 130079 29957
rect 130091 29945 130125 30569
rect 130137 30557 130138 30558
rect 130736 30557 130737 30558
rect 130136 30556 130137 30557
rect 130737 30556 130738 30557
rect 130136 29957 130137 29958
rect 130737 29957 130738 29958
rect 130137 29956 130138 29957
rect 130736 29956 130737 29957
rect 130749 29945 130783 30569
rect 130795 30557 130796 30558
rect 131394 30557 131395 30558
rect 130794 30556 130795 30557
rect 131395 30556 131396 30557
rect 130794 29957 130795 29958
rect 131395 29957 131396 29958
rect 130795 29956 130796 29957
rect 131394 29956 131395 29957
rect 131407 29945 131441 30569
rect 131453 30557 131454 30558
rect 132052 30557 132053 30558
rect 131452 30556 131453 30557
rect 132053 30556 132054 30557
rect 131452 29957 131453 29958
rect 132053 29957 132054 29958
rect 131453 29956 131454 29957
rect 132052 29956 132053 29957
rect 132065 29945 132099 30569
rect 132111 30557 132112 30558
rect 132110 30556 132111 30557
rect 132608 30553 132689 30588
rect 132717 30579 132723 30581
rect 132608 30541 132695 30553
rect 132621 30492 132640 30541
rect 132649 30492 132695 30541
rect 132717 30520 132727 30579
rect 132655 30044 132702 30492
rect 132110 29957 132111 29958
rect 132111 29956 132112 29957
rect 132596 29945 132607 29956
rect 129319 29911 132607 29945
rect 132621 29933 132640 30044
rect 132649 29973 132695 30044
rect 132649 29961 132668 29973
rect 132689 29961 132695 29973
rect 132717 30016 132730 30520
rect 132717 29935 132727 30016
rect 132717 29933 132723 29935
rect 129319 29287 129353 29911
rect 129433 29287 129467 29911
rect 129479 29899 129480 29900
rect 130078 29899 130079 29900
rect 129478 29898 129479 29899
rect 130079 29898 130080 29899
rect 129478 29299 129479 29300
rect 130079 29299 130080 29300
rect 129479 29298 129480 29299
rect 130078 29298 130079 29299
rect 130091 29287 130125 29911
rect 130137 29899 130138 29900
rect 130736 29899 130737 29900
rect 130136 29898 130137 29899
rect 130737 29898 130738 29899
rect 130136 29299 130137 29300
rect 130737 29299 130738 29300
rect 130137 29298 130138 29299
rect 130736 29298 130737 29299
rect 130749 29287 130783 29911
rect 130795 29899 130796 29900
rect 131394 29899 131395 29900
rect 130794 29898 130795 29899
rect 131395 29898 131396 29899
rect 130794 29299 130795 29300
rect 131395 29299 131396 29300
rect 130795 29298 130796 29299
rect 131394 29298 131395 29299
rect 131407 29287 131441 29911
rect 131453 29899 131454 29900
rect 132052 29899 132053 29900
rect 131452 29898 131453 29899
rect 132053 29898 132054 29899
rect 131452 29299 131453 29300
rect 132053 29299 132054 29300
rect 131453 29298 131454 29299
rect 132052 29298 132053 29299
rect 132065 29287 132099 29911
rect 132111 29899 132112 29900
rect 132110 29898 132111 29899
rect 132608 29895 132689 29930
rect 132717 29921 132723 29923
rect 132608 29883 132695 29895
rect 132621 29822 132640 29883
rect 132649 29822 132695 29883
rect 132717 29850 132727 29921
rect 132655 29374 132702 29822
rect 132110 29299 132111 29300
rect 132111 29298 132112 29299
rect 132596 29287 132607 29298
rect 129319 29253 132607 29287
rect 132621 29275 132640 29374
rect 132649 29315 132695 29374
rect 132649 29303 132668 29315
rect 132689 29303 132695 29315
rect 132717 29346 132730 29850
rect 132717 29277 132727 29346
rect 132717 29275 132723 29277
rect 128214 29056 128604 29090
rect 127838 28589 128094 28592
rect 127866 28561 128066 28564
rect 128214 28558 128248 29056
rect 128428 28988 128475 29035
rect 128390 28954 128475 28988
rect 128317 28895 128362 28906
rect 128445 28895 128490 28906
rect 128328 28719 128362 28895
rect 128456 28719 128490 28895
rect 128428 28663 128475 28707
rect 128390 28641 128475 28663
rect 128374 28629 128475 28641
rect 128374 28610 128444 28629
rect 128570 28592 128604 29056
rect 128314 28589 128604 28592
rect 128348 28572 128468 28589
rect 128342 28561 128542 28564
rect 128342 28558 128496 28561
rect 128570 28558 128604 28589
rect 128214 28524 128604 28558
rect 128690 29056 129080 29090
rect 128690 28558 128724 29056
rect 128904 28988 128951 29035
rect 128866 28954 128951 28988
rect 128793 28895 128838 28906
rect 128921 28895 128966 28906
rect 128804 28719 128838 28895
rect 128932 28719 128966 28895
rect 128904 28663 128951 28707
rect 128866 28641 128951 28663
rect 128850 28629 128951 28641
rect 128850 28610 128920 28629
rect 128824 28572 128944 28574
rect 129046 28558 129080 29056
rect 128690 28524 129080 28558
rect 129319 28629 129353 29253
rect 129433 28629 129467 29253
rect 129479 29241 129480 29242
rect 130078 29241 130079 29242
rect 129478 29240 129479 29241
rect 130079 29240 130080 29241
rect 129478 28641 129479 28642
rect 130079 28641 130080 28642
rect 129479 28640 129480 28641
rect 130078 28640 130079 28641
rect 130091 28629 130125 29253
rect 130137 29241 130138 29242
rect 130736 29241 130737 29242
rect 130136 29240 130137 29241
rect 130737 29240 130738 29241
rect 130136 28641 130137 28642
rect 130737 28641 130738 28642
rect 130137 28640 130138 28641
rect 130736 28640 130737 28641
rect 130749 28629 130783 29253
rect 130795 29241 130796 29242
rect 131394 29241 131395 29242
rect 130794 29240 130795 29241
rect 131395 29240 131396 29241
rect 130794 28641 130795 28642
rect 131395 28641 131396 28642
rect 130795 28640 130796 28641
rect 131394 28640 131395 28641
rect 131407 28629 131441 29253
rect 131453 29241 131454 29242
rect 132052 29241 132053 29242
rect 131452 29240 131453 29241
rect 132053 29240 132054 29241
rect 131452 28641 131453 28642
rect 132053 28641 132054 28642
rect 131453 28640 131454 28641
rect 132052 28640 132053 28641
rect 132065 28629 132099 29253
rect 132111 29241 132112 29242
rect 132110 29240 132111 29241
rect 132608 29237 132689 29272
rect 132717 29263 132723 29265
rect 132608 29225 132695 29237
rect 132621 29160 132640 29225
rect 132649 29160 132695 29225
rect 132717 29160 132727 29263
rect 132655 28712 132689 29160
rect 132723 28712 132727 29160
rect 132110 28641 132111 28642
rect 132111 28640 132112 28641
rect 132596 28629 132607 28640
rect 129319 28595 132607 28629
rect 132621 28617 132640 28712
rect 132649 28657 132695 28712
rect 132649 28645 132668 28657
rect 132689 28645 132695 28657
rect 132717 28619 132727 28712
rect 132717 28617 132723 28619
rect 128196 28368 128618 28474
rect 128672 28368 129094 28474
rect 128196 28156 129094 28368
rect 128196 27964 128618 28156
rect 128672 27964 129094 28156
rect 129319 27971 129353 28595
rect 129433 27971 129467 28595
rect 129479 28583 129480 28584
rect 130078 28583 130079 28584
rect 129478 28582 129479 28583
rect 130079 28582 130080 28583
rect 129478 27983 129479 27984
rect 130079 27983 130080 27984
rect 129479 27982 129480 27983
rect 130078 27982 130079 27983
rect 130091 27971 130125 28595
rect 130137 28583 130138 28584
rect 130736 28583 130737 28584
rect 130136 28582 130137 28583
rect 130737 28582 130738 28583
rect 130136 27983 130137 27984
rect 130737 27983 130738 27984
rect 130137 27982 130138 27983
rect 130736 27982 130737 27983
rect 130749 27971 130783 28595
rect 130795 28583 130796 28584
rect 131394 28583 131395 28584
rect 130794 28582 130795 28583
rect 131395 28582 131396 28583
rect 130794 27983 130795 27984
rect 131395 27983 131396 27984
rect 130795 27982 130796 27983
rect 131394 27982 131395 27983
rect 131407 27971 131441 28595
rect 131453 28583 131454 28584
rect 132052 28583 132053 28584
rect 131452 28582 131453 28583
rect 132053 28582 132054 28583
rect 131452 27983 131453 27984
rect 132053 27983 132054 27984
rect 131453 27982 131454 27983
rect 132052 27982 132053 27983
rect 132065 27971 132099 28595
rect 132111 28583 132112 28584
rect 132110 28582 132111 28583
rect 132608 28579 132689 28614
rect 132717 28605 132723 28607
rect 132608 28567 132695 28579
rect 132621 28502 132640 28567
rect 132649 28502 132695 28567
rect 132717 28530 132727 28605
rect 132655 28054 132702 28502
rect 132110 27983 132111 27984
rect 132111 27982 132112 27983
rect 132596 27971 132607 27982
rect 124389 27937 129096 27964
rect 129319 27937 132607 27971
rect 132621 27959 132640 28054
rect 132649 27999 132695 28054
rect 132649 27987 132668 27999
rect 132689 27987 132695 27999
rect 132717 28026 132730 28530
rect 132717 27961 132727 28026
rect 132717 27959 132723 27961
rect 121855 27852 121901 27867
rect 121876 27821 121901 27852
rect 124389 27857 127830 27937
rect 128196 27930 128618 27937
rect 128672 27930 129094 27937
rect 127848 27903 129094 27930
rect 128196 27860 128618 27903
rect 128672 27860 129094 27903
rect 127924 27857 129094 27860
rect 129319 27857 129353 27937
rect 129433 27920 129467 27937
rect 130091 27920 130125 27937
rect 130749 27920 130783 27937
rect 131407 27920 131441 27937
rect 132065 27920 132099 27937
rect 132757 27911 132769 31279
rect 129421 27908 129479 27911
rect 130079 27908 130137 27911
rect 130737 27908 130795 27911
rect 131395 27908 131453 27911
rect 132053 27908 132111 27911
rect 132711 27908 132769 27911
rect 129495 27861 130063 27891
rect 130153 27861 130721 27891
rect 130811 27861 131379 27891
rect 131469 27861 132037 27891
rect 132127 27861 132695 27891
rect 124389 27846 130090 27857
rect 130126 27846 130748 27857
rect 130784 27846 131406 27857
rect 131442 27846 132064 27857
rect 132100 27846 132722 27857
rect 124389 27834 130079 27846
rect 130137 27834 130737 27846
rect 130795 27834 131395 27846
rect 131453 27834 132053 27846
rect 132111 27834 132711 27846
rect 124389 27827 130090 27834
rect 130126 27827 130748 27834
rect 130784 27827 131406 27834
rect 131442 27827 132064 27834
rect 132100 27827 132722 27834
rect 124389 27823 132722 27827
rect 132837 27823 132845 31429
rect 134390 29782 134424 34130
rect 135820 33666 135854 34130
rect 135508 33224 135854 33666
rect 135820 29782 135854 33224
rect 136318 32554 136352 34130
rect 136380 34048 136394 34130
rect 136408 34076 136523 34130
rect 136386 33972 136394 34048
rect 136414 34012 136523 34076
rect 136414 34000 136460 34012
rect 136466 33997 136523 34012
rect 137136 33997 137181 34130
rect 136466 33996 136524 33997
rect 137124 33996 137125 33997
rect 137136 33996 137182 33997
rect 137782 33996 137783 33997
rect 137794 33996 137839 34130
rect 136472 33984 136512 33996
rect 136524 33995 136525 33996
rect 137123 33995 137124 33996
rect 136524 33984 137124 33995
rect 137136 33984 137170 33996
rect 137182 33995 137183 33996
rect 137781 33995 137782 33996
rect 137182 33984 137782 33995
rect 137794 33984 137828 33996
rect 137908 33984 137942 34130
rect 136472 33972 137942 33984
rect 136478 33962 137942 33972
rect 136386 33960 136394 33962
rect 136472 33960 137942 33962
rect 136382 33950 137942 33960
rect 136382 33938 136512 33950
rect 136524 33938 136525 33939
rect 137123 33938 137124 33939
rect 137136 33938 137170 33950
rect 137182 33938 137183 33939
rect 137781 33938 137782 33939
rect 137794 33938 137828 33950
rect 136382 33937 136524 33938
rect 137124 33937 137125 33938
rect 137136 33937 137182 33938
rect 137782 33937 137783 33938
rect 136382 33922 136523 33937
rect 136386 33314 136394 33922
rect 136414 33866 136523 33922
rect 136414 33418 136546 33866
rect 136414 33354 136523 33418
rect 136414 33342 136460 33354
rect 136466 33339 136523 33354
rect 137136 33339 137181 33937
rect 136466 33338 136524 33339
rect 137124 33338 137125 33339
rect 137136 33338 137182 33339
rect 137782 33338 137783 33339
rect 137794 33338 137839 33938
rect 136472 33326 136512 33338
rect 136524 33337 136525 33338
rect 137123 33337 137124 33338
rect 136524 33326 137124 33337
rect 137136 33326 137170 33338
rect 137182 33337 137183 33338
rect 137781 33337 137782 33338
rect 137182 33326 137782 33337
rect 137794 33326 137828 33338
rect 137908 33326 137942 33950
rect 136472 33314 137942 33326
rect 136478 33304 137942 33314
rect 136386 33302 136394 33304
rect 136472 33302 137942 33304
rect 136382 33292 137942 33302
rect 136382 33280 136512 33292
rect 136524 33280 136525 33281
rect 137123 33280 137124 33281
rect 137136 33280 137170 33292
rect 137182 33280 137183 33281
rect 137781 33280 137782 33281
rect 137794 33280 137828 33292
rect 136382 33279 136524 33280
rect 137124 33279 137125 33280
rect 137136 33279 137182 33280
rect 137782 33279 137783 33280
rect 136382 33264 136523 33279
rect 136386 33242 136394 33264
rect 136380 32738 136394 33242
rect 136414 33214 136523 33264
rect 136408 33172 136523 33214
rect 137136 33172 137181 33279
rect 137794 33172 137839 33280
rect 136408 32766 136454 33172
rect 136386 32656 136394 32738
rect 136414 32684 136460 32766
rect 136444 32680 136454 32684
rect 136466 32680 136512 33172
rect 136523 32680 136524 32681
rect 137124 32680 137125 32681
rect 136472 32668 136512 32680
rect 136524 32679 136525 32680
rect 137123 32679 137124 32680
rect 137136 32668 137170 33172
rect 137181 32680 137182 32681
rect 137782 32680 137783 32681
rect 137182 32679 137183 32680
rect 137781 32679 137782 32680
rect 137794 32668 137828 33172
rect 137908 32668 137942 33292
rect 136472 32656 137942 32668
rect 136478 32634 137942 32656
rect 136478 32554 136512 32634
rect 137136 32554 137170 32634
rect 137794 32554 137828 32634
rect 137908 32554 137942 32634
rect 144632 32616 144666 35244
rect 147742 34944 153662 35528
rect 147742 34928 153702 34944
rect 147742 34680 153662 34928
rect 153702 34864 153718 34928
rect 153950 34864 153954 34944
rect 147742 34577 153663 34680
rect 153701 34616 153702 34617
rect 153702 34615 153703 34616
rect 153716 34577 153743 34620
rect 147742 34576 153662 34577
rect 147742 34256 153886 34576
rect 154117 34493 154165 35995
rect 154245 36005 154279 36057
rect 154903 36036 154937 36057
rect 155561 36036 155595 36057
rect 156219 36036 156253 36057
rect 156877 36036 156911 36057
rect 154861 36005 154937 36036
rect 155519 36005 155595 36036
rect 156177 36005 156253 36036
rect 156835 36005 156911 36036
rect 154245 35908 154291 36005
rect 154861 35989 154949 36005
rect 155519 35989 155607 36005
rect 156177 35989 156265 36005
rect 156835 35989 156923 36005
rect 156934 35995 156948 36057
rect 157017 36036 157051 36057
rect 157131 36054 157176 36057
rect 157535 36054 157580 36057
rect 157131 36036 157165 36054
rect 157535 36036 157569 36054
rect 157017 35989 157064 36036
rect 157131 36005 157178 36036
rect 157119 35989 157178 36005
rect 157493 35989 157569 36036
rect 154293 35955 154949 35989
rect 154951 35955 155607 35989
rect 155609 35955 156265 35989
rect 156267 35955 156923 35989
rect 156925 35955 157569 35989
rect 154869 35949 154873 35955
rect 154897 35921 154901 35955
rect 154903 35908 154949 35955
rect 155561 35908 155607 35955
rect 156185 35949 156189 35955
rect 156213 35921 156217 35955
rect 156219 35908 156265 35955
rect 156877 35908 156923 35955
rect 154245 35896 154279 35908
rect 154878 35896 154891 35907
rect 154903 35896 154937 35908
rect 155536 35896 155549 35907
rect 155561 35896 155595 35908
rect 156194 35896 156207 35907
rect 156219 35896 156253 35908
rect 156852 35896 156865 35907
rect 156877 35896 156911 35908
rect 154231 34592 154279 35896
rect 154889 34592 154937 35896
rect 155547 34592 155595 35896
rect 154231 34520 154265 34592
rect 154889 34580 154923 34592
rect 155547 34580 155581 34592
rect 154267 34520 154271 34567
rect 154295 34533 154299 34539
rect 154875 34533 154923 34580
rect 155533 34533 155581 34580
rect 147742 34255 153662 34256
rect 147742 34148 153663 34255
rect 153702 34216 153703 34217
rect 153701 34215 153702 34216
rect 153716 34208 153743 34255
rect 147742 32944 153662 34148
rect 136318 32520 141848 32554
rect 137374 31604 137586 32052
rect 137908 31037 137942 32520
rect 136259 31001 137978 31037
rect 141501 31001 141535 31499
rect 136259 30967 144661 31001
rect 134504 27934 134538 27938
rect 134466 27896 134576 27900
rect 135128 27884 135140 28040
rect 135162 27918 135174 28074
rect 134294 27850 135134 27884
rect 124389 27820 127830 27823
rect 124206 27818 124242 27820
rect 124276 27818 127830 27820
rect 124389 27787 127830 27818
rect 127924 27787 128894 27823
rect 129319 27821 129353 27823
rect 124240 27784 124242 27786
rect 124276 27784 124496 27786
rect 127796 27504 127808 27786
rect 127830 27538 127842 27760
rect 136259 27712 137978 30967
rect 138362 29056 138752 29090
rect 138362 28913 138396 29056
rect 138576 28988 138623 29035
rect 138538 28954 138623 28988
rect 138522 28913 138592 28925
rect 138718 28913 138752 29056
rect 138362 28879 138752 28913
rect 138362 28558 138396 28879
rect 138476 28719 138510 28879
rect 138522 28867 138523 28868
rect 138591 28867 138592 28868
rect 138521 28866 138522 28867
rect 138592 28866 138593 28867
rect 138604 28719 138638 28879
rect 138458 28558 138468 28698
rect 138486 28568 138524 28670
rect 138576 28660 138623 28707
rect 138538 28626 138623 28660
rect 138718 28558 138752 28879
rect 138362 28524 138752 28558
rect 138838 29056 139228 29090
rect 138838 28913 138872 29056
rect 139052 29026 139099 29035
rect 138960 29000 139099 29026
rect 139052 28998 139099 29000
rect 138988 28972 139099 28998
rect 139014 28954 139099 28972
rect 138988 28946 139060 28947
rect 138998 28919 139068 28925
rect 138960 28918 139088 28919
rect 138998 28913 139068 28918
rect 139194 28913 139228 29056
rect 138838 28879 139228 28913
rect 138838 28558 138872 28879
rect 138952 28719 138986 28879
rect 138998 28867 138999 28868
rect 139067 28867 139068 28868
rect 138997 28866 138998 28867
rect 139068 28866 139069 28867
rect 139080 28719 139114 28879
rect 139052 28660 139099 28707
rect 139014 28626 139099 28660
rect 139194 28558 139228 28879
rect 138838 28524 139228 28558
rect 138344 27854 138766 28474
rect 138820 27854 139242 28474
rect 141501 28077 141535 30967
rect 141590 30916 141597 30921
rect 141643 30916 142796 30921
rect 144148 30916 144506 30921
rect 141556 30893 141684 30899
rect 144466 30893 144477 30898
rect 141556 30888 142796 30893
rect 144148 30888 144478 30893
rect 141556 30887 141684 30888
rect 144466 30887 144477 30888
rect 141556 30857 144477 30887
rect 144478 30857 144559 30872
rect 141556 30853 144559 30857
rect 141587 30847 142796 30853
rect 144148 30847 144559 30853
rect 141587 30841 141684 30847
rect 144478 30835 144559 30847
rect 144478 30829 144575 30835
rect 141684 30823 142796 30829
rect 144148 30823 144575 30829
rect 144627 30823 144661 30967
rect 141680 30819 144575 30823
rect 141556 30761 141637 30808
rect 141696 30798 144575 30819
rect 144593 30798 144695 30823
rect 141684 30789 144695 30798
rect 141684 30783 144606 30789
rect 144478 30777 144575 30783
rect 141574 30258 141597 30263
rect 141603 30242 141637 30761
rect 141656 30755 144519 30770
rect 141952 30263 143466 30291
rect 141643 30258 144506 30263
rect 144525 30257 144559 30777
rect 144565 30755 144578 30770
rect 141556 30241 141637 30242
rect 141556 30235 141684 30241
rect 144466 30235 144477 30240
rect 141546 30230 144478 30235
rect 141556 30229 141684 30230
rect 144466 30229 144477 30230
rect 141556 30199 144477 30229
rect 144478 30199 144559 30214
rect 141556 30195 144559 30199
rect 141587 30189 142008 30195
rect 143410 30189 144559 30195
rect 141587 30183 141684 30189
rect 144478 30177 144559 30189
rect 144478 30171 144575 30177
rect 141684 30165 142008 30171
rect 143410 30165 144575 30171
rect 144627 30165 144661 30789
rect 141680 30161 149672 30165
rect 141556 30103 141637 30150
rect 141696 30146 149672 30161
rect 141684 30131 149672 30146
rect 141684 30125 142008 30131
rect 143410 30125 144606 30131
rect 144478 30119 144575 30125
rect 141590 29596 141597 29605
rect 141603 29584 141637 30103
rect 141656 30097 142008 30118
rect 143410 30097 144519 30118
rect 141643 29596 142826 29605
rect 144178 29596 144506 29605
rect 144525 29599 144559 30119
rect 144565 30097 144578 30118
rect 141556 29583 141637 29584
rect 141556 29577 141684 29583
rect 144466 29577 144477 29582
rect 141556 29571 142826 29577
rect 144178 29571 144478 29577
rect 141556 29568 144478 29571
rect 141556 29541 144477 29568
rect 144478 29541 144559 29556
rect 141556 29537 144559 29541
rect 141587 29531 142826 29537
rect 144178 29531 144559 29537
rect 141587 29525 141684 29531
rect 144478 29519 144559 29531
rect 144478 29513 144575 29519
rect 141684 29507 142826 29513
rect 144178 29507 144575 29513
rect 144627 29507 144661 30131
rect 154117 29782 154151 34493
rect 154231 34431 154271 34520
rect 154291 34520 154299 34533
rect 154307 34520 154923 34533
rect 154291 34499 154923 34520
rect 154949 34499 154957 34533
rect 154965 34499 155581 34533
rect 154295 34493 154348 34499
rect 154290 34465 154348 34492
rect 154877 34483 154923 34499
rect 155535 34483 155581 34499
rect 154290 34431 154299 34465
rect 154889 34431 154923 34483
rect 155547 34431 155581 34483
rect 155583 34465 155587 34567
rect 156128 34539 156130 35636
rect 156156 34539 156158 35608
rect 156205 34592 156253 35896
rect 156863 34592 156911 35896
rect 156934 34882 156948 35949
rect 157017 34727 157051 35955
rect 157119 35908 157177 35955
rect 157131 34888 157165 35908
rect 157535 35907 157569 35955
rect 157510 35896 157569 35907
rect 157521 34876 157569 35896
rect 157509 34829 157581 34876
rect 157193 34795 157581 34829
rect 157450 34727 157452 34782
rect 157478 34727 157480 34782
rect 157509 34779 157581 34795
rect 157521 34764 157581 34779
rect 157521 34727 157569 34764
rect 157635 34727 157683 36057
rect 158426 35632 158500 36258
rect 158412 35478 158566 35632
rect 159071 34848 159090 37372
rect 159099 34876 159118 37372
rect 159166 36132 160605 40784
rect 161948 39626 161982 40784
rect 161210 38932 161672 39570
rect 161882 39544 161982 39626
rect 161268 38848 161618 38882
rect 161268 38820 161302 38848
rect 161268 38430 161336 38820
rect 161460 38780 161498 38818
rect 161426 38746 161498 38780
rect 161371 38696 161416 38707
rect 161459 38696 161504 38707
rect 161382 38520 161416 38696
rect 161470 38520 161504 38696
rect 161460 38470 161498 38508
rect 161426 38436 161498 38470
rect 161268 38368 161302 38430
rect 161584 38368 161618 38848
rect 161268 38334 161618 38368
rect 161910 38216 161946 38302
rect 159152 36096 160605 36132
rect 160632 36096 160666 36130
rect 161290 36096 161324 36130
rect 161948 36096 161982 39544
rect 162018 39150 162020 39228
rect 162018 36096 162020 36262
rect 162088 36096 162122 40784
rect 162202 39910 162247 40784
rect 162202 36096 162236 39910
rect 162606 39884 162651 40784
rect 162606 36096 162640 39884
rect 162720 36096 162754 40784
rect 162860 36127 162894 42136
rect 163170 41524 163632 42162
rect 163646 41524 164108 42162
rect 163224 41440 163574 41474
rect 163224 40960 163258 41440
rect 163416 41372 163454 41410
rect 163382 41338 163454 41372
rect 163327 41288 163372 41299
rect 163415 41288 163460 41299
rect 163338 41112 163372 41288
rect 163426 41112 163460 41288
rect 163416 41062 163454 41100
rect 163382 41028 163454 41062
rect 163540 40960 163574 41440
rect 163224 40926 163574 40960
rect 163700 41440 164050 41474
rect 163700 40960 163734 41440
rect 163892 41372 163930 41410
rect 163858 41338 163930 41372
rect 163803 41288 163848 41299
rect 163891 41288 163936 41299
rect 163814 41112 163848 41288
rect 163902 41112 163936 41288
rect 163892 41062 163930 41100
rect 163858 41028 163930 41062
rect 164016 40960 164050 41440
rect 163700 40926 164050 40960
rect 162896 40808 162932 40894
rect 165492 36127 165526 42878
rect 159152 36062 162754 36096
rect 159152 36032 160605 36062
rect 159152 35960 160628 36032
rect 160632 36010 160666 36062
rect 161248 36028 161286 36032
rect 159152 34829 160605 35960
rect 160632 35922 160678 36010
rect 161248 35994 161288 36028
rect 160680 35960 161288 35994
rect 161244 35954 161260 35960
rect 161284 35954 161288 35960
rect 161272 35926 161288 35954
rect 161290 36010 161324 36062
rect 161290 35922 161336 36010
rect 161906 35994 161944 36032
rect 161338 35960 161944 35994
rect 161948 36010 161982 36062
rect 161948 35922 161994 36010
rect 162004 36000 162020 36062
rect 162074 36026 162076 36062
rect 162060 36000 162076 36026
rect 162088 36032 162122 36062
rect 162202 36032 162236 36062
rect 162088 35994 162126 36032
rect 162202 36010 162240 36032
rect 162190 35994 162248 36010
rect 162564 35994 162602 36032
rect 161996 35960 162602 35994
rect 160607 35910 160620 35921
rect 160632 35910 160666 35922
rect 161265 35910 161278 35921
rect 161290 35910 161324 35922
rect 161923 35910 161936 35921
rect 161948 35910 161982 35922
rect 159151 34795 160605 34829
rect 159152 34727 160605 34795
rect 157017 34693 160605 34727
rect 156205 34580 156239 34592
rect 156863 34580 156897 34592
rect 155611 34533 155615 34539
rect 156191 34533 156239 34580
rect 156849 34533 156897 34580
rect 155607 34499 155615 34533
rect 155623 34499 156239 34533
rect 156265 34499 156273 34533
rect 156281 34499 156897 34533
rect 155611 34493 155615 34499
rect 156128 34486 156130 34493
rect 156156 34458 156158 34493
rect 156193 34483 156239 34499
rect 156851 34483 156897 34499
rect 156205 34431 156239 34483
rect 156863 34431 156897 34483
rect 156899 34465 156903 34567
rect 157450 34539 157452 34693
rect 157478 34539 157480 34693
rect 157521 34592 157569 34693
rect 157521 34580 157555 34592
rect 156927 34533 156931 34539
rect 157507 34533 157555 34580
rect 156923 34499 156931 34533
rect 156939 34499 157555 34533
rect 156927 34493 156931 34499
rect 157450 34486 157452 34493
rect 157478 34458 157480 34493
rect 157509 34483 157555 34499
rect 157521 34431 157555 34483
rect 157635 34493 157683 34693
rect 159152 34657 160605 34693
rect 159188 34516 159236 34657
rect 159302 34606 159350 34657
rect 154219 34397 157567 34431
rect 154262 34264 154271 34397
rect 154290 34292 154299 34397
rect 156864 34052 156903 34397
rect 156920 34052 156931 34348
rect 157635 29782 157669 34493
rect 159188 29782 159222 34516
rect 159302 34454 159336 34606
rect 159338 34488 159342 34590
rect 159888 34562 159896 34657
rect 159916 34562 159924 34657
rect 159960 34606 160008 34657
rect 160618 34606 160666 35910
rect 161276 34606 161324 35910
rect 161352 34804 161372 35328
rect 161934 34606 161982 35910
rect 162004 34860 162020 35954
rect 162060 34818 162076 35954
rect 162088 34750 162122 35960
rect 162190 35922 162248 35960
rect 162202 34902 162236 35922
rect 162606 35921 162640 36062
rect 162581 35910 162640 35921
rect 162592 34890 162640 35910
rect 162580 34852 162652 34890
rect 162264 34818 162652 34852
rect 162516 34750 162522 34806
rect 162544 34750 162550 34806
rect 162580 34802 162652 34818
rect 162592 34787 162652 34802
rect 162592 34750 162640 34787
rect 162706 34750 162754 36062
rect 162837 36091 165676 36127
rect 165773 36091 165807 42963
rect 165887 36091 165921 42864
rect 162837 36058 166425 36091
rect 162837 36057 166450 36058
rect 162762 35350 162782 35980
rect 162837 35952 165676 36057
rect 165681 35955 165687 35989
rect 162790 35936 165676 35952
rect 162790 35674 165687 35936
rect 162790 35458 165676 35674
rect 162790 35378 165687 35458
rect 162837 35258 165687 35378
rect 162837 35236 165676 35258
rect 162762 34934 162782 35190
rect 162826 35162 165676 35236
rect 165692 35202 165746 35228
rect 162790 35058 165676 35162
rect 162790 34962 165687 35058
rect 162778 34858 162782 34934
rect 162837 34932 165687 34962
rect 162806 34858 165687 34932
rect 162837 34812 165676 34858
rect 162778 34806 162782 34812
rect 162806 34762 165676 34812
rect 162790 34750 165676 34762
rect 162088 34716 165676 34750
rect 159960 34594 159994 34606
rect 160618 34594 160652 34606
rect 161276 34594 161310 34606
rect 161934 34594 161968 34606
rect 162516 34594 162522 34716
rect 162544 34594 162550 34716
rect 162592 34606 162640 34716
rect 162592 34594 162626 34606
rect 159366 34556 159370 34562
rect 159946 34556 159994 34594
rect 160604 34556 160652 34594
rect 159362 34522 159370 34556
rect 159378 34522 159994 34556
rect 160020 34522 160028 34556
rect 160036 34522 160652 34556
rect 159366 34516 159370 34522
rect 159888 34510 159896 34516
rect 159916 34482 159924 34516
rect 159948 34506 159994 34522
rect 160606 34506 160652 34522
rect 159960 34454 159994 34506
rect 160618 34454 160652 34506
rect 160654 34488 160658 34590
rect 160682 34556 160686 34562
rect 161262 34556 161310 34594
rect 161920 34556 161968 34594
rect 160678 34522 160686 34556
rect 160694 34522 161310 34556
rect 161336 34522 161344 34556
rect 161352 34522 161968 34556
rect 160682 34516 160686 34522
rect 161264 34506 161310 34522
rect 161922 34506 161968 34522
rect 161276 34454 161310 34506
rect 161934 34454 161968 34506
rect 161970 34488 161976 34590
rect 161998 34556 162004 34562
rect 162086 34556 162626 34594
rect 161994 34522 162004 34556
rect 162010 34522 162626 34556
rect 161998 34516 162004 34522
rect 162516 34504 162522 34516
rect 162544 34482 162550 34516
rect 162580 34506 162626 34522
rect 162592 34454 162626 34506
rect 162706 34516 162754 34716
rect 162837 34680 165676 34716
rect 165773 34727 165807 36057
rect 165887 36020 165934 36036
rect 165875 35989 165934 36020
rect 166060 36024 166450 36057
rect 166060 35996 166094 36024
rect 166249 36003 166296 36024
rect 166026 35989 166128 35996
rect 166249 35989 166321 36003
rect 165875 35955 166321 35989
rect 165875 35908 165933 35955
rect 165887 34898 165921 35908
rect 166060 35526 166094 35955
rect 166236 35922 166321 35955
rect 166277 35907 166311 35912
rect 166266 35896 166311 35907
rect 166277 35879 166311 35896
rect 166277 35874 166322 35879
rect 166163 35863 166208 35874
rect 166174 35687 166208 35863
rect 166277 35687 166336 35874
rect 166277 35675 166322 35687
rect 166274 35671 166322 35675
rect 166274 35628 166321 35671
rect 166236 35594 166321 35628
rect 166277 35526 166311 35594
rect 166391 35526 166450 36024
rect 166060 35492 166450 35526
rect 166536 36024 166926 36058
rect 166536 35996 166570 36024
rect 166536 35588 166604 35996
rect 166750 35956 166797 36003
rect 166712 35922 166797 35956
rect 166639 35863 166684 35874
rect 166767 35863 166812 35874
rect 166650 35687 166684 35863
rect 166778 35687 166812 35863
rect 166750 35628 166797 35675
rect 166712 35594 166797 35628
rect 166536 35526 166570 35588
rect 166892 35526 166926 36024
rect 166536 35492 166926 35526
rect 166277 35442 166311 35492
rect 166391 35442 166425 35492
rect 165887 34888 165932 34898
rect 166042 34876 166464 35442
rect 165902 34829 166464 34876
rect 165949 34822 166464 34829
rect 166518 34822 166940 35442
rect 167827 34848 167830 37372
rect 167855 34876 167858 37372
rect 167908 36096 169361 36132
rect 170844 36096 170878 42968
rect 220506 39050 221858 39052
rect 214604 38548 214660 38564
rect 214170 37779 222146 37813
rect 167908 36062 171496 36096
rect 167908 34829 169361 36062
rect 170000 35954 170016 35982
rect 170028 35928 170044 35954
rect 170712 35926 170732 36028
rect 170740 35954 170760 36000
rect 165949 34795 166425 34822
rect 167907 34795 169361 34829
rect 166265 34779 166323 34795
rect 166277 34764 166323 34779
rect 166277 34727 166311 34764
rect 166391 34727 166425 34795
rect 167908 34727 169361 34795
rect 165773 34693 169361 34727
rect 170844 34750 170878 36062
rect 170958 36025 170996 36032
rect 170946 36010 170996 36025
rect 170946 35994 171004 36010
rect 171320 35994 171358 36032
rect 170946 35960 171358 35994
rect 170946 35922 171004 35960
rect 170958 34902 170992 35922
rect 171337 35910 171382 35921
rect 171348 34890 171382 35910
rect 171336 34852 171394 34890
rect 171020 34818 171394 34852
rect 171336 34802 171394 34818
rect 171379 34787 171394 34802
rect 171348 34750 171382 34784
rect 171462 34750 171496 36062
rect 174950 35540 175070 35560
rect 175256 35542 175496 36094
rect 175256 35540 175546 35542
rect 174944 35512 175098 35532
rect 175256 35514 175496 35540
rect 175256 35512 175574 35514
rect 175256 35456 175496 35512
rect 175885 35456 175972 36348
rect 214633 36112 218293 36145
rect 219704 36112 222312 36146
rect 185098 35540 185218 35560
rect 185404 35542 185644 36094
rect 214651 36066 218275 36112
rect 219758 36084 222312 36096
rect 219758 36078 222380 36084
rect 214651 36054 218442 36066
rect 219792 36062 222226 36078
rect 222278 36062 222380 36078
rect 214651 36032 218275 36054
rect 219758 36037 222172 36044
rect 219758 36034 219792 36037
rect 219724 36032 219826 36034
rect 210508 36000 210534 36032
rect 210938 36000 210956 36032
rect 214648 36020 218476 36032
rect 219724 36028 222176 36032
rect 185404 35540 185694 35542
rect 185092 35512 185246 35532
rect 185404 35514 185644 35540
rect 185404 35512 185722 35514
rect 185404 35456 185644 35512
rect 170844 34716 174300 34750
rect 159290 34420 162638 34454
rect 159960 29782 159994 34420
rect 162706 29782 162740 34516
rect 162949 34444 162950 34530
rect 162806 34384 162981 34404
rect 162768 33654 162816 33662
rect 162768 33620 162782 33628
rect 162987 29782 163021 34680
rect 163156 34526 163578 34680
rect 163632 34526 164054 34680
rect 165636 34624 165659 34680
rect 166277 34586 166311 34693
rect 165620 34176 165659 34404
rect 165613 34120 165659 34176
rect 165620 33858 165659 34120
rect 165613 33104 165659 33858
rect 165676 33160 165687 34348
rect 166391 29782 166425 34693
rect 167908 34657 169361 34693
rect 171462 29782 171496 34716
rect 174398 34472 174410 34754
rect 174432 34506 174444 34728
rect 183516 33104 183716 33126
rect 209762 31966 209764 32022
rect 209762 31710 209764 31766
rect 209762 31566 209764 31622
rect 209762 31310 209764 31366
rect 141680 29503 144575 29507
rect 141556 29445 141637 29492
rect 141696 29476 144575 29503
rect 144593 29476 144695 29507
rect 141684 29473 144695 29476
rect 141684 29467 144606 29473
rect 144478 29461 144575 29467
rect 141590 28926 141597 28947
rect 141603 28926 141637 29445
rect 141656 29439 144519 29448
rect 142770 29411 144234 29439
rect 141930 28947 143444 28975
rect 141643 28926 144506 28947
rect 144525 28941 144559 29461
rect 144565 29439 144578 29448
rect 141556 28925 141637 28926
rect 141556 28919 141684 28925
rect 144466 28919 144477 28924
rect 141556 28898 144478 28919
rect 141556 28883 144477 28898
rect 144478 28883 144559 28898
rect 141556 28879 144559 28883
rect 141587 28873 141986 28879
rect 143388 28873 144559 28879
rect 141587 28867 141684 28873
rect 144478 28861 144559 28873
rect 144478 28855 144575 28861
rect 141684 28849 141986 28855
rect 143388 28849 144575 28855
rect 144627 28849 144661 29473
rect 172106 29090 172140 29782
rect 172186 29090 172194 29280
rect 172214 29124 172222 29308
rect 172214 29090 172244 29124
rect 163160 29056 163550 29090
rect 141680 28845 144575 28849
rect 141556 28787 141637 28834
rect 141696 28815 144575 28845
rect 144593 28815 144695 28849
rect 143388 28814 144228 28815
rect 144478 28814 144575 28815
rect 141684 28809 141986 28814
rect 143388 28809 144575 28814
rect 144478 28803 144575 28809
rect 141590 28274 141597 28289
rect 141603 28268 141637 28787
rect 141656 28781 141986 28786
rect 143388 28781 144519 28786
rect 141643 28274 142820 28289
rect 144172 28274 144506 28289
rect 144525 28283 144559 28803
rect 141556 28267 141637 28268
rect 141556 28261 141684 28267
rect 144466 28261 144477 28266
rect 141556 28255 142820 28261
rect 144172 28255 144478 28261
rect 141556 28246 144478 28255
rect 141556 28225 144477 28246
rect 144478 28225 144559 28240
rect 141556 28221 144559 28225
rect 141587 28215 142820 28221
rect 144172 28215 144559 28221
rect 141587 28209 141684 28215
rect 144478 28203 144559 28215
rect 144478 28197 144575 28203
rect 141684 28191 142820 28197
rect 144172 28191 144575 28197
rect 144627 28191 144661 28815
rect 163160 28558 163194 29056
rect 163374 28988 163421 29035
rect 163336 28954 163421 28988
rect 163263 28895 163308 28906
rect 163391 28895 163436 28906
rect 163274 28719 163308 28895
rect 163402 28719 163436 28895
rect 163374 28660 163421 28707
rect 163336 28626 163421 28660
rect 163516 28558 163550 29056
rect 163160 28524 163550 28558
rect 163636 29056 164026 29090
rect 172012 29056 172306 29090
rect 163636 29028 163670 29056
rect 163636 28620 163704 29028
rect 163850 28988 163897 29035
rect 163812 28954 163897 28988
rect 163739 28895 163784 28906
rect 163867 28895 163912 28906
rect 163750 28719 163784 28895
rect 163878 28719 163912 28895
rect 163850 28660 163897 28707
rect 163812 28626 163897 28660
rect 163636 28558 163670 28620
rect 163992 28558 164026 29056
rect 172106 29022 172140 29056
rect 172106 28954 172164 29022
rect 172106 28694 172140 28954
rect 172158 28703 172174 28911
rect 172186 28907 172194 29056
rect 172214 28961 172222 29056
rect 172238 28961 172254 29056
rect 172186 28902 172198 28907
rect 172186 28895 172192 28902
rect 172182 28719 172192 28895
rect 172186 28703 172192 28719
rect 172208 28732 172258 28961
rect 172208 28707 172266 28732
rect 172106 28626 172164 28694
rect 172106 28592 172140 28626
rect 172166 28592 172170 28668
rect 172050 28572 172170 28592
rect 172106 28564 172140 28572
rect 172194 28564 172198 28696
rect 172044 28558 172198 28564
rect 172210 28558 172266 28707
rect 172272 28558 172306 29056
rect 163636 28524 164026 28558
rect 172012 28524 172306 28558
rect 172392 29056 172782 29090
rect 172392 28558 172426 29056
rect 172606 28988 172653 29035
rect 172568 28954 172653 28988
rect 172495 28895 172540 28906
rect 172623 28895 172668 28906
rect 172506 28719 172540 28895
rect 172634 28719 172668 28895
rect 172444 28558 172464 28706
rect 172606 28660 172653 28707
rect 172568 28626 172653 28660
rect 172748 28558 172782 29056
rect 172392 28524 172782 28558
rect 204826 29056 205216 29090
rect 204826 28558 204860 29056
rect 205040 28988 205087 29035
rect 205002 28954 205087 28988
rect 204929 28895 204974 28906
rect 205057 28895 205102 28906
rect 204940 28719 204974 28895
rect 205068 28719 205102 28895
rect 205040 28660 205087 28707
rect 205002 28626 205087 28660
rect 205182 28558 205216 29056
rect 204826 28524 205216 28558
rect 205302 29056 205692 29090
rect 205302 29028 205336 29056
rect 205302 28620 205370 29028
rect 205516 28988 205563 29035
rect 205478 28954 205563 28988
rect 205405 28895 205450 28906
rect 205533 28895 205578 28906
rect 205416 28719 205450 28895
rect 205544 28719 205578 28895
rect 205516 28660 205563 28707
rect 205478 28626 205563 28660
rect 205302 28558 205336 28620
rect 205658 28558 205692 29056
rect 205302 28524 205692 28558
rect 172106 28474 172140 28524
rect 172210 28522 172266 28524
rect 172146 28474 172266 28522
rect 141680 28187 144575 28191
rect 141696 28160 144575 28187
rect 141696 28157 144590 28160
rect 144593 28157 144695 28191
rect 144478 28156 144590 28157
rect 141684 28151 144606 28156
rect 144478 28145 144590 28151
rect 141656 28123 144519 28128
rect 144565 28123 144578 28128
rect 142764 28095 144228 28123
rect 144627 28077 144661 28157
rect 141501 28043 149771 28077
rect 136414 27625 136431 27684
rect 136452 27597 136469 27646
rect 136534 27597 137154 27712
rect 137204 27676 137238 27712
rect 137582 27700 137615 27704
rect 137736 27700 137770 27712
rect 137582 27681 137790 27700
rect 137388 27680 137790 27681
rect 137388 27676 137586 27680
rect 137204 27638 137244 27676
rect 137388 27672 137587 27676
rect 137736 27672 137770 27680
rect 137388 27670 137790 27672
rect 137259 27648 137387 27655
rect 137252 27638 137387 27648
rect 137194 27624 137202 27630
rect 137204 27618 137238 27638
rect 137244 27624 137387 27638
rect 137399 27652 137790 27670
rect 137399 27636 137586 27652
rect 137259 27618 137387 27624
rect 137587 27618 137715 27652
rect 137736 27618 137770 27652
rect 137204 27597 137860 27618
rect 136452 27564 137154 27597
rect 137170 27564 141848 27597
rect 136452 27563 141848 27564
rect 136534 27413 137154 27563
rect 137204 27551 137860 27563
rect 137206 27544 137860 27551
rect 144627 27545 144661 28043
rect 163142 27861 163564 28474
rect 163049 27827 163617 27861
rect 163618 27854 164040 28474
rect 172070 28110 172320 28474
rect 172374 28110 172796 28474
rect 172136 28060 172170 28070
rect 172524 28060 172558 28070
rect 172612 28060 172646 28070
rect 172152 28026 172204 28036
rect 172490 28026 172680 28036
rect 172118 27992 172142 28026
rect 172152 27958 172176 28026
rect 172250 27924 172284 27936
rect 172028 27890 172284 27924
rect 172410 27924 172444 27936
rect 172726 27924 172760 27936
rect 172410 27890 172760 27924
rect 204808 27861 205230 28474
rect 204715 27827 205283 27861
rect 205284 27854 205706 28474
rect 210508 27950 210534 35954
rect 210938 27950 210956 35954
rect 212350 35910 212396 35922
rect 212356 35898 212396 35910
rect 211658 34224 211670 35328
rect 212386 32614 212396 35898
rect 214651 35122 218275 36020
rect 219724 35998 219792 36028
rect 219884 35998 222176 36028
rect 222312 36010 222323 36021
rect 222335 36010 222346 36021
rect 219758 35374 219792 35998
rect 219918 35964 220540 35998
rect 220576 35964 221198 35998
rect 221234 35964 221856 35998
rect 221892 35994 222172 35998
rect 222312 35994 222346 36010
rect 221892 35964 222346 35994
rect 219934 35960 220540 35964
rect 220592 35960 221198 35964
rect 221250 35960 221856 35964
rect 221908 35960 222346 35964
rect 222171 35922 222172 35923
rect 222172 35921 222173 35922
rect 219861 35910 219906 35921
rect 220519 35910 220564 35921
rect 221177 35910 221222 35921
rect 221835 35910 221880 35921
rect 219872 35374 219906 35910
rect 219917 35386 219918 35387
rect 220518 35386 220519 35387
rect 219918 35385 219919 35386
rect 220517 35385 220518 35386
rect 220530 35374 220564 35910
rect 220575 35386 220576 35387
rect 221176 35386 221177 35387
rect 220576 35385 220577 35386
rect 221175 35385 221176 35386
rect 221188 35374 221222 35910
rect 221233 35386 221234 35387
rect 221834 35386 221835 35387
rect 221234 35385 221235 35386
rect 221833 35385 221834 35386
rect 221846 35374 221880 35910
rect 222210 35402 222244 35960
rect 221891 35386 221892 35387
rect 221892 35385 221893 35386
rect 222160 35374 222171 35385
rect 219724 35340 222171 35374
rect 214651 34910 218316 35122
rect 214651 32628 218275 34910
rect 219758 34716 219792 35340
rect 219872 34716 219906 35340
rect 219918 35328 219919 35329
rect 220517 35328 220518 35329
rect 219917 35327 219918 35328
rect 220518 35327 220519 35328
rect 219917 34728 219918 34729
rect 220518 34728 220519 34729
rect 219918 34727 219919 34728
rect 220517 34727 220518 34728
rect 220530 34716 220564 35340
rect 220576 35328 220577 35329
rect 221175 35328 221176 35329
rect 220575 35327 220576 35328
rect 221176 35327 221177 35328
rect 220575 34728 220576 34729
rect 221176 34728 221177 34729
rect 220576 34727 220577 34728
rect 221175 34727 221176 34728
rect 221188 34716 221222 35340
rect 221778 35334 221840 35340
rect 221234 35328 221235 35329
rect 221833 35328 221834 35329
rect 221233 35327 221234 35328
rect 221806 35306 221840 35328
rect 221233 34728 221234 34729
rect 221834 34728 221835 34729
rect 221234 34727 221235 34728
rect 221833 34727 221834 34728
rect 221846 34716 221880 35340
rect 221886 35334 221970 35340
rect 221892 35328 221893 35329
rect 221886 35306 221942 35328
rect 222172 35312 222244 35350
rect 222210 34744 222244 35312
rect 221891 34728 221892 34729
rect 221892 34727 221893 34728
rect 222160 34716 222171 34727
rect 219724 34682 222171 34716
rect 219758 34058 219792 34682
rect 219872 34058 219906 34682
rect 219918 34670 219919 34671
rect 220517 34670 220518 34671
rect 219917 34669 219918 34670
rect 220518 34669 220519 34670
rect 219917 34070 219918 34071
rect 219918 34069 219919 34070
rect 220446 34064 220452 34126
rect 220474 34064 220480 34098
rect 220518 34070 220519 34071
rect 220517 34069 220518 34070
rect 220530 34058 220564 34682
rect 220576 34670 220577 34671
rect 221175 34670 221176 34671
rect 220575 34669 220576 34670
rect 221176 34669 221177 34670
rect 220575 34070 220576 34071
rect 221176 34070 221177 34071
rect 220576 34069 220577 34070
rect 221175 34069 221176 34070
rect 221188 34058 221222 34682
rect 221234 34670 221235 34671
rect 221833 34670 221834 34671
rect 221233 34669 221234 34670
rect 221834 34669 221835 34670
rect 221233 34070 221234 34071
rect 221834 34070 221835 34071
rect 221234 34069 221235 34070
rect 221833 34069 221834 34070
rect 221846 34058 221880 34682
rect 221892 34670 221893 34671
rect 221891 34669 221892 34670
rect 222172 34654 222244 34692
rect 222210 34086 222244 34654
rect 221891 34070 221892 34071
rect 221892 34069 221893 34070
rect 222160 34058 222171 34069
rect 219724 34024 222171 34058
rect 219758 33400 219792 34024
rect 219872 33400 219906 34024
rect 219918 34012 219919 34013
rect 219917 34011 219918 34012
rect 220446 33934 220452 34018
rect 220474 33962 220480 34018
rect 220517 34012 220518 34013
rect 220518 34011 220519 34012
rect 219917 33412 219918 33413
rect 220518 33412 220519 33413
rect 219918 33411 219919 33412
rect 220517 33411 220518 33412
rect 220530 33400 220564 34024
rect 220576 34012 220577 34013
rect 221175 34012 221176 34013
rect 220575 34011 220576 34012
rect 221176 34011 221177 34012
rect 220575 33412 220576 33413
rect 221176 33412 221177 33413
rect 220576 33411 220577 33412
rect 221175 33411 221176 33412
rect 221188 33400 221222 34024
rect 221234 34012 221235 34013
rect 221833 34012 221834 34013
rect 221233 34011 221234 34012
rect 221834 34011 221835 34012
rect 221233 33412 221234 33413
rect 221834 33412 221835 33413
rect 221234 33411 221235 33412
rect 221833 33411 221834 33412
rect 221846 33400 221880 34024
rect 221892 34012 221893 34013
rect 221891 34011 221892 34012
rect 222172 33996 222244 34034
rect 222210 33428 222244 33996
rect 221891 33412 221892 33413
rect 221892 33411 221893 33412
rect 222160 33400 222171 33411
rect 219724 33366 222171 33400
rect 219758 32742 219792 33366
rect 219872 32742 219906 33366
rect 219918 33354 219919 33355
rect 220517 33354 220518 33355
rect 219917 33353 219918 33354
rect 220518 33353 220519 33354
rect 219917 32754 219918 32755
rect 219918 32753 219919 32754
rect 220448 32748 220452 32818
rect 220476 32748 220480 32790
rect 220518 32754 220519 32755
rect 220517 32753 220518 32754
rect 220530 32742 220564 33366
rect 220576 33354 220577 33355
rect 221175 33354 221176 33355
rect 220575 33353 220576 33354
rect 221176 33353 221177 33354
rect 220575 32754 220576 32755
rect 221176 32754 221177 32755
rect 220576 32753 220577 32754
rect 221175 32753 221176 32754
rect 221188 32742 221222 33366
rect 221234 33354 221235 33355
rect 221833 33354 221834 33355
rect 221233 33353 221234 33354
rect 221834 33353 221835 33354
rect 221233 32754 221234 32755
rect 221834 32754 221835 32755
rect 221234 32753 221235 32754
rect 221833 32753 221834 32754
rect 221846 32742 221880 33366
rect 221892 33354 221893 33355
rect 221891 33353 221892 33354
rect 222172 33338 222244 33376
rect 222210 32770 222244 33338
rect 221891 32754 221892 32755
rect 221892 32753 221893 32754
rect 222160 32742 222171 32753
rect 219724 32708 222171 32742
rect 219758 32628 219792 32708
rect 219872 32628 219906 32708
rect 220448 32628 220452 32702
rect 220476 32654 220480 32702
rect 220530 32628 220564 32708
rect 221188 32628 221222 32708
rect 221846 32628 221880 32708
rect 222312 32628 222346 35960
rect 214651 32594 222346 32628
rect 214651 32558 218275 32594
rect 218880 32558 219342 32594
rect 214687 32223 214721 32558
rect 215421 32420 215432 32506
rect 215459 32382 215470 32544
rect 218205 32223 218239 32558
rect 218916 32223 218950 32470
rect 219272 32223 219306 32470
rect 219758 32259 219792 32594
rect 219722 32223 222395 32259
rect 214089 32189 222395 32223
rect 214104 32109 214724 32189
rect 214801 32174 214835 32189
rect 214774 32140 215340 32174
rect 214774 32112 214835 32140
rect 215306 32128 215340 32140
rect 215459 32128 215493 32189
rect 214740 32109 214835 32112
rect 214904 32109 215558 32128
rect 216117 32109 216151 32189
rect 216775 32109 216809 32189
rect 217433 32109 217467 32189
rect 218091 32109 218125 32189
rect 218205 32109 218239 32189
rect 214104 32078 218239 32109
rect 214104 32047 214724 32078
rect 214740 32075 218239 32078
rect 214095 32008 214724 32047
rect 214022 31922 214724 32008
rect 214095 31770 214724 31922
rect 214774 32045 214835 32075
rect 214847 32063 214848 32064
rect 214846 32062 214847 32063
rect 214904 32054 215558 32075
rect 216104 32063 216105 32064
rect 216105 32062 216106 32063
rect 214953 32045 215232 32054
rect 214774 31998 214910 32045
rect 214953 32041 215238 32045
rect 214969 32026 215238 32041
rect 214774 31818 214835 31998
rect 214876 31960 214910 31998
rect 215020 31960 215238 32026
rect 215020 31932 215232 31960
rect 214969 31898 215232 31932
rect 215020 31818 215232 31898
rect 215306 31818 215340 32054
rect 215421 31944 215432 32030
rect 214774 31784 215340 31818
rect 214095 31716 214129 31770
rect 214687 31716 214721 31770
rect 214095 31479 214724 31716
rect 214801 31698 214835 31784
rect 215020 31698 215232 31784
rect 214104 31294 214724 31479
rect 214774 31664 215340 31698
rect 214774 31569 214835 31664
rect 215020 31650 215232 31664
rect 215145 31584 215156 31595
rect 214774 31522 214910 31569
rect 214969 31550 215156 31584
rect 215157 31522 215238 31569
rect 214774 31451 214835 31522
rect 214876 31468 214910 31522
rect 215204 31468 215238 31522
rect 214846 31463 214847 31464
rect 214847 31462 214848 31463
rect 215145 31462 215156 31467
rect 215306 31462 215340 31664
rect 215459 31464 215504 32054
rect 215447 31463 215448 31464
rect 215459 31463 215505 31464
rect 216105 31463 216106 31464
rect 215446 31462 215447 31463
rect 214953 31456 214969 31462
rect 215145 31456 215161 31462
rect 214953 31451 215161 31456
rect 215306 31451 215447 31462
rect 215459 31451 215493 31463
rect 215505 31462 215506 31463
rect 216104 31462 216105 31463
rect 215505 31451 215530 31462
rect 216117 31451 216151 32075
rect 216163 32063 216164 32064
rect 216762 32063 216763 32064
rect 216162 32062 216163 32063
rect 216763 32062 216764 32063
rect 216162 31463 216163 31464
rect 216763 31463 216764 31464
rect 216163 31462 216164 31463
rect 216762 31462 216763 31463
rect 216775 31451 216809 32075
rect 216821 32063 216822 32064
rect 217420 32063 217421 32064
rect 216820 32062 216821 32063
rect 217421 32062 217422 32063
rect 216820 31463 216821 31464
rect 217421 31463 217422 31464
rect 216821 31462 216822 31463
rect 217420 31462 217421 31463
rect 217433 31451 217467 32075
rect 217479 32063 217480 32064
rect 218078 32063 218079 32064
rect 217478 32062 217479 32063
rect 218079 32062 218080 32063
rect 218091 31890 218125 32075
rect 218205 31890 218239 32075
rect 218916 32034 218950 32189
rect 219092 32136 219130 32143
rect 219061 32109 219177 32121
rect 219061 32106 219161 32109
rect 219076 32086 219146 32106
rect 219272 32034 219306 32189
rect 218916 32000 219306 32034
rect 218340 31918 218458 31998
rect 218314 31890 218458 31918
rect 217918 31866 218458 31890
rect 217918 31678 218366 31866
rect 217478 31463 217479 31464
rect 218079 31463 218080 31464
rect 217479 31462 217480 31463
rect 218078 31462 218079 31463
rect 218091 31451 218125 31678
rect 218205 31451 218239 31678
rect 214740 31417 218239 31451
rect 218902 31440 219324 31950
rect 218900 31417 219706 31440
rect 214774 31342 214835 31417
rect 214847 31405 214848 31406
rect 214846 31404 214847 31405
rect 215306 31342 215340 31417
rect 215446 31405 215447 31406
rect 215459 31405 215493 31417
rect 215505 31405 215506 31406
rect 216104 31405 216105 31406
rect 215447 31404 215448 31405
rect 215459 31404 215505 31405
rect 216105 31404 216106 31405
rect 214774 31308 215340 31342
rect 215459 31310 215504 31404
rect 214687 30793 214721 31294
rect 214801 30793 214835 31308
rect 214846 30805 214847 30806
rect 215447 30805 215448 30806
rect 214847 30804 214848 30805
rect 215446 30804 215447 30805
rect 215459 30793 215493 31310
rect 215504 30805 215505 30806
rect 216105 30805 216106 30806
rect 215505 30804 215506 30805
rect 216104 30804 216105 30805
rect 216117 30793 216151 31417
rect 216163 31405 216164 31406
rect 216762 31405 216763 31406
rect 216162 31404 216163 31405
rect 216763 31404 216764 31405
rect 216162 30805 216163 30806
rect 216763 30805 216764 30806
rect 216163 30804 216164 30805
rect 216762 30804 216763 30805
rect 216775 30793 216809 31417
rect 216821 31405 216822 31406
rect 217420 31405 217421 31406
rect 216820 31404 216821 31405
rect 217421 31404 217422 31405
rect 216820 30805 216821 30806
rect 217421 30805 217422 30806
rect 216821 30804 216822 30805
rect 217420 30804 217421 30805
rect 217433 30793 217467 31417
rect 217479 31405 217480 31406
rect 218078 31405 218079 31406
rect 217478 31404 217479 31405
rect 218079 31404 218080 31405
rect 217478 30805 217479 30806
rect 218079 30805 218080 30806
rect 217479 30804 217480 30805
rect 218078 30804 218079 30805
rect 218091 30793 218125 31417
rect 218205 30793 218239 31417
rect 218902 31406 219324 31417
rect 218902 31383 219672 31406
rect 218902 31330 219324 31383
rect 214653 30759 218239 30793
rect 214687 30700 214721 30759
rect 214602 30690 214795 30700
rect 214687 30672 214721 30690
rect 214574 30662 214795 30672
rect 214687 30135 214721 30662
rect 214801 30135 214835 30759
rect 214847 30747 214848 30748
rect 215446 30747 215447 30748
rect 214846 30746 214847 30747
rect 215447 30746 215448 30747
rect 214846 30147 214847 30148
rect 215447 30147 215448 30148
rect 214847 30146 214848 30147
rect 215446 30146 215447 30147
rect 215459 30135 215493 30759
rect 215505 30747 215506 30748
rect 216104 30747 216105 30748
rect 215504 30746 215505 30747
rect 216105 30746 216106 30747
rect 215504 30147 215505 30148
rect 216105 30147 216106 30148
rect 215505 30146 215506 30147
rect 216104 30146 216105 30147
rect 216117 30135 216151 30759
rect 216163 30747 216164 30748
rect 216762 30747 216763 30748
rect 216162 30746 216163 30747
rect 216763 30746 216764 30747
rect 216162 30147 216163 30148
rect 216763 30147 216764 30148
rect 216163 30146 216164 30147
rect 216762 30146 216763 30147
rect 216775 30135 216809 30759
rect 216821 30747 216822 30748
rect 217420 30747 217421 30748
rect 216820 30746 216821 30747
rect 217421 30746 217422 30747
rect 216820 30147 216821 30148
rect 217421 30147 217422 30148
rect 216821 30146 216822 30147
rect 217420 30146 217421 30147
rect 217433 30135 217467 30759
rect 217479 30747 217480 30748
rect 218078 30747 218079 30748
rect 217478 30746 217479 30747
rect 218079 30746 218080 30747
rect 217478 30147 217479 30148
rect 218079 30147 218080 30148
rect 217479 30146 217480 30147
rect 218078 30146 218079 30147
rect 218091 30135 218125 30759
rect 218205 30135 218239 30759
rect 214653 30101 218239 30135
rect 212404 28188 212428 29590
rect 214687 29477 214721 30101
rect 214801 29477 214835 30101
rect 214847 30089 214848 30090
rect 215446 30089 215447 30090
rect 214846 30088 214847 30089
rect 215447 30088 215448 30089
rect 214846 29489 214847 29490
rect 215447 29489 215448 29490
rect 214847 29488 214848 29489
rect 215446 29488 215447 29489
rect 215459 29477 215493 30101
rect 215505 30089 215506 30090
rect 216104 30089 216105 30090
rect 215504 30088 215505 30089
rect 216105 30088 216106 30089
rect 215504 29489 215505 29490
rect 216105 29489 216106 29490
rect 215505 29488 215506 29489
rect 216104 29488 216105 29489
rect 216117 29477 216151 30101
rect 216163 30089 216164 30090
rect 216762 30089 216763 30090
rect 216162 30088 216163 30089
rect 216763 30088 216764 30089
rect 216162 29489 216163 29490
rect 216763 29489 216764 29490
rect 216163 29488 216164 29489
rect 216762 29488 216763 29489
rect 216775 29477 216809 30101
rect 216821 30089 216822 30090
rect 217420 30089 217421 30090
rect 216820 30088 216821 30089
rect 217421 30088 217422 30089
rect 216820 29489 216821 29490
rect 217421 29489 217422 29490
rect 216821 29488 216822 29489
rect 217420 29488 217421 29489
rect 217433 29477 217467 30101
rect 217479 30089 217480 30090
rect 218078 30089 218079 30090
rect 217478 30088 217479 30089
rect 218079 30088 218080 30089
rect 217478 29489 217479 29490
rect 218079 29489 218080 29490
rect 217479 29488 217480 29489
rect 218078 29488 218079 29489
rect 218091 29477 218125 30101
rect 218205 29477 218239 30101
rect 214653 29443 218239 29477
rect 213646 28902 213648 29308
rect 213674 28902 213704 29280
rect 213993 29090 214027 29144
rect 213993 29058 214026 29090
rect 213959 28637 213972 29058
rect 213993 28705 214027 29058
rect 214058 29056 214448 29090
rect 214058 28705 214092 29056
rect 214095 28831 214126 29056
rect 214272 28988 214319 29035
rect 214234 28954 214319 28988
rect 214414 28924 214448 29056
rect 214160 28906 214176 28907
rect 214160 28819 214206 28906
rect 214289 28895 214334 28906
rect 214340 28902 214634 28924
rect 214414 28896 214448 28902
rect 214217 28831 214218 28832
rect 214288 28831 214289 28832
rect 214218 28830 214219 28831
rect 214287 28830 214288 28831
rect 214300 28819 214334 28895
rect 214340 28874 214606 28896
rect 214414 28819 214448 28874
rect 214687 28819 214721 29443
rect 214801 28819 214835 29443
rect 214847 29431 214848 29432
rect 215446 29431 215447 29432
rect 214846 29430 214847 29431
rect 215447 29430 215448 29431
rect 214846 28831 214847 28832
rect 215447 28831 215448 28832
rect 214847 28830 214848 28831
rect 215446 28830 215447 28831
rect 215459 28819 215493 29443
rect 215505 29431 215506 29432
rect 216104 29431 216105 29432
rect 215504 29430 215505 29431
rect 216105 29430 216106 29431
rect 215504 28831 215505 28832
rect 216105 28831 216106 28832
rect 215505 28830 215506 28831
rect 216104 28830 216105 28831
rect 216117 28819 216151 29443
rect 216163 29431 216164 29432
rect 216762 29431 216763 29432
rect 216162 29430 216163 29431
rect 216763 29430 216764 29431
rect 216162 28831 216163 28832
rect 216763 28831 216764 28832
rect 216163 28830 216164 28831
rect 216762 28830 216763 28831
rect 216775 28819 216809 29443
rect 216821 29431 216822 29432
rect 217420 29431 217421 29432
rect 216820 29430 216821 29431
rect 217421 29430 217422 29431
rect 216820 28831 216821 28832
rect 217421 28831 217422 28832
rect 216821 28830 216822 28831
rect 217420 28830 217421 28831
rect 217433 28819 217467 29443
rect 217479 29431 217480 29432
rect 218078 29431 218079 29432
rect 217478 29430 217479 29431
rect 218079 29430 218080 29431
rect 217478 28831 217479 28832
rect 218079 28831 218080 28832
rect 217479 28830 217480 28831
rect 218078 28830 218079 28831
rect 218091 28819 218125 29443
rect 218205 28819 218239 29443
rect 214160 28816 214448 28819
rect 214172 28785 214448 28816
rect 214653 28785 218239 28819
rect 214172 28759 214206 28785
rect 214300 28759 214334 28785
rect 214160 28707 214218 28759
rect 214288 28707 214346 28759
rect 214414 28705 214448 28785
rect 214687 28705 214721 28785
rect 214801 28705 214835 28785
rect 215459 28705 215493 28785
rect 216117 28705 216151 28785
rect 216775 28705 216809 28785
rect 217433 28705 217467 28785
rect 218091 28705 218125 28785
rect 218205 28705 218239 28785
rect 219722 28705 222395 32189
rect 223708 29044 224080 29748
rect 213993 28671 214026 28705
rect 214058 28671 222395 28705
rect 214058 28635 214092 28671
rect 214218 28637 214288 28660
rect 213716 28572 213836 28592
rect 214022 28574 214262 28635
rect 214414 28620 214448 28671
rect 214687 28635 214721 28671
rect 214022 28572 214312 28574
rect 213710 28544 213864 28564
rect 214022 28546 214262 28572
rect 214022 28544 214340 28546
rect 214022 28488 214262 28544
rect 214651 28488 214738 28635
rect 212356 27934 212396 27946
rect 212350 27922 212396 27934
rect 172228 27712 172232 27802
rect 172256 27728 172260 27774
rect 137399 27537 137575 27542
rect 137224 27522 137244 27530
rect 137252 27528 137272 27530
rect 137204 27490 137238 27517
rect 137387 27496 137587 27537
rect 137736 27490 137770 27517
rect 213164 27504 213176 27786
rect 213198 27538 213210 27760
rect 213690 27712 213704 28066
rect 214687 27821 214721 28488
rect 218205 28008 218239 28671
rect 219722 28635 222395 28671
rect 221170 28624 221244 28635
rect 224170 28488 224410 29126
rect 217598 27759 218239 28008
rect 217598 27689 218218 27759
rect 218234 27725 218239 27759
rect 218268 27725 218293 27994
rect 218268 27700 218273 27725
rect 137387 27482 137587 27483
rect 137238 27449 137736 27482
rect 213732 27428 213808 27430
rect 213732 27426 213804 27428
rect 213704 27400 213836 27402
rect 213704 27398 213832 27400
rect 128178 26968 128640 27215
rect 145903 27156 145920 27212
rect 213696 27183 213730 27188
rect 213824 27183 213858 27188
rect 213662 27149 213764 27154
rect 213790 27149 213892 27154
rect 213962 27152 213972 27206
rect 213980 26968 214008 27188
rect 214016 27004 214026 27152
rect 214202 27004 222178 27038
rect 117588 26874 118376 26892
rect 117622 26840 118342 26858
rect 127866 26844 128066 26845
rect 127838 26816 128094 26817
rect 97603 26079 97844 26137
rect 95617 25574 96374 25585
rect 97603 25574 97826 26079
rect 95628 25540 97826 25574
rect 97603 25479 97826 25540
rect 97603 25460 97844 25479
rect 95497 25426 97844 25460
rect 97603 25421 97844 25426
rect 97603 25283 97826 25421
rect 96374 24854 96412 24884
rect 96374 24820 96378 24850
rect 95482 21950 95502 23622
rect 95538 21846 95558 23678
rect 51001 20428 59439 20464
rect 44868 20394 59439 20428
rect 73078 20394 82586 20464
rect 44868 19766 44902 20394
rect 46400 20366 46434 20378
rect 45712 20326 45750 20364
rect 46366 20332 46386 20338
rect 46394 20332 46434 20366
rect 46400 20326 46434 20332
rect 45044 20292 45750 20326
rect 45802 20292 46486 20326
rect 46361 20254 46362 20255
rect 46362 20253 46363 20254
rect 44971 20242 45016 20253
rect 45729 20242 45774 20253
rect 44982 19766 45016 20242
rect 45027 19778 45028 19779
rect 45728 19778 45729 19779
rect 45028 19777 45029 19778
rect 45727 19777 45728 19778
rect 45740 19766 45774 20242
rect 46400 19850 46434 20292
rect 46464 19850 46472 20282
rect 45785 19778 45786 19779
rect 45786 19777 45787 19778
rect 46350 19766 46361 19777
rect 44834 19732 46361 19766
rect 46366 19754 46386 19850
rect 46394 19794 46434 19850
rect 46492 19822 46500 20254
rect 46394 19782 46414 19794
rect 46366 19742 46386 19744
rect 44868 19108 44902 19732
rect 44982 19108 45016 19732
rect 45028 19720 45029 19721
rect 45727 19720 45728 19721
rect 45027 19719 45028 19720
rect 45728 19719 45729 19720
rect 45027 19120 45028 19121
rect 45728 19120 45729 19121
rect 45028 19119 45029 19120
rect 45727 19119 45728 19120
rect 45740 19108 45774 19732
rect 45786 19720 45787 19721
rect 45785 19719 45786 19720
rect 46362 19704 46434 19742
rect 46366 19634 46386 19704
rect 46394 19634 46434 19704
rect 46400 19186 46434 19634
rect 45785 19120 45786 19121
rect 45786 19119 45787 19120
rect 46350 19108 46361 19119
rect 44834 19074 46361 19108
rect 46366 19096 46386 19186
rect 46394 19136 46434 19186
rect 46394 19124 46414 19136
rect 46366 19084 46386 19086
rect 44868 18450 44902 19074
rect 44982 18450 45016 19074
rect 45028 19062 45029 19063
rect 45727 19062 45728 19063
rect 45027 19061 45028 19062
rect 45728 19061 45729 19062
rect 45027 18462 45028 18463
rect 45728 18462 45729 18463
rect 45028 18461 45029 18462
rect 45727 18461 45728 18462
rect 45740 18450 45774 19074
rect 45786 19062 45787 19063
rect 45785 19061 45786 19062
rect 46362 19046 46434 19084
rect 46366 18982 46386 19046
rect 46394 18982 46434 19046
rect 46400 18534 46434 18982
rect 46464 18534 46466 18982
rect 45785 18462 45786 18463
rect 45786 18461 45787 18462
rect 46350 18450 46361 18461
rect 44834 18416 46361 18450
rect 46366 18438 46386 18534
rect 46394 18478 46434 18534
rect 46492 18506 46494 19010
rect 46394 18466 46414 18478
rect 44868 18336 44902 18416
rect 44982 18336 45016 18416
rect 45740 18336 45774 18416
rect 46502 18336 46536 20394
rect 46544 20292 46583 20326
rect 41048 18302 46536 18336
rect 51001 18315 59439 20394
rect 60250 20390 60450 20392
rect 73018 20332 73028 20338
rect 73074 20332 82586 20394
rect 73078 20286 82586 20332
rect 43978 18146 43992 18296
rect 44006 18174 44020 18302
rect 38984 17696 39004 17754
rect 39012 17696 39032 17748
rect 43978 17746 43992 18002
rect 44006 17774 44020 17974
rect 38928 17456 39566 17696
rect 38984 17124 38986 17300
rect 39012 17152 39014 17272
rect 44868 16663 44902 18302
rect 38792 16398 38992 16424
rect 38764 16370 39020 16396
rect 23390 16026 23410 16084
rect 23418 16026 23438 16078
rect 23334 15786 23972 16026
rect 21062 15630 22184 15678
rect 21006 15574 22240 15622
rect 23390 15454 23392 15630
rect 23418 15482 23420 15602
rect 44832 15542 46467 16663
rect 48884 15650 48900 16654
rect 48912 15650 48956 16710
rect 57110 15862 57144 18315
rect 60194 17134 60222 17190
rect 55352 15828 58904 15862
rect 54836 15694 54876 15706
rect 54830 15682 54876 15694
rect 55352 15542 55386 15828
rect 55460 15766 55476 15822
rect 57110 15798 57144 15828
rect 55594 15776 55632 15798
rect 55582 15760 55640 15776
rect 56096 15760 56134 15798
rect 56352 15776 56390 15798
rect 56340 15760 56398 15776
rect 56754 15760 56792 15798
rect 57110 15776 57148 15798
rect 57098 15760 57156 15776
rect 57412 15760 57450 15798
rect 57868 15776 57906 15798
rect 57856 15760 57914 15776
rect 58070 15760 58108 15798
rect 58626 15776 58664 15798
rect 58614 15760 58672 15776
rect 58728 15760 58766 15798
rect 58768 15766 58796 15822
rect 55528 15726 56134 15760
rect 56186 15726 56792 15760
rect 56844 15726 57450 15760
rect 57502 15726 58108 15760
rect 58160 15726 58766 15760
rect 55582 15688 55640 15726
rect 56340 15688 56398 15726
rect 57098 15688 57156 15726
rect 57856 15688 57914 15726
rect 58614 15688 58672 15726
rect 58750 15687 58752 15688
rect 55455 15682 55500 15687
rect 56113 15682 56158 15687
rect 56771 15682 56816 15687
rect 57429 15682 57474 15687
rect 58087 15682 58132 15687
rect 58745 15682 58790 15687
rect 55454 15644 55512 15682
rect 55566 15644 55604 15682
rect 56112 15644 56170 15682
rect 56324 15644 56362 15682
rect 56770 15644 56828 15682
rect 57082 15644 57120 15682
rect 57428 15644 57486 15682
rect 57840 15644 57878 15682
rect 58086 15644 58144 15682
rect 58598 15644 58636 15682
rect 58744 15680 58802 15682
rect 58726 15650 58802 15680
rect 58744 15644 58802 15650
rect 55454 15610 55604 15644
rect 55656 15610 56362 15644
rect 56414 15610 57120 15644
rect 57172 15610 57878 15644
rect 57930 15610 58636 15644
rect 58688 15610 58802 15644
rect 55454 15594 55512 15610
rect 56112 15594 56170 15610
rect 56770 15594 56828 15610
rect 57428 15594 57486 15610
rect 58086 15594 58144 15610
rect 58744 15594 58802 15610
rect 55454 15579 55469 15594
rect 58787 15579 58802 15594
rect 55466 15542 55500 15576
rect 56124 15542 56158 15576
rect 56782 15542 56816 15576
rect 57440 15542 57474 15576
rect 58098 15542 58132 15576
rect 58756 15542 58790 15576
rect 58870 15542 58904 15828
rect 59378 15682 59424 15706
rect 60136 15682 60182 15706
rect 60311 15542 63935 20157
rect 65418 20092 68970 20126
rect 72396 20112 72416 20242
rect 72434 20170 72610 20222
rect 72430 20146 72912 20170
rect 72506 20108 72912 20146
rect 73018 20108 73028 20286
rect 73074 20108 82586 20286
rect 64540 15994 65002 16632
rect 64598 15910 64948 15944
rect 64598 15542 64632 15910
rect 64690 15804 64724 15910
rect 64730 15896 64774 15910
rect 64730 15880 64820 15894
rect 64730 15868 64828 15880
rect 64790 15842 64828 15868
rect 64740 15808 64828 15842
rect 64802 15804 64820 15808
rect 64690 15772 64730 15804
rect 64736 15800 64758 15804
rect 64802 15800 64812 15804
rect 64830 15776 64848 15910
rect 64830 15772 64840 15776
rect 64690 15758 64724 15772
rect 64736 15758 64746 15769
rect 64789 15758 64834 15769
rect 64690 15694 64746 15758
rect 64712 15682 64746 15694
rect 64800 15682 64834 15758
rect 64712 15644 64758 15682
rect 64788 15644 64846 15682
rect 64712 15610 64846 15644
rect 64712 15596 64758 15610
rect 64700 15594 64758 15596
rect 64788 15594 64846 15610
rect 64700 15582 64746 15594
rect 64700 15576 64740 15582
rect 64806 15576 64846 15594
rect 64700 15570 64746 15576
rect 64712 15566 64746 15570
rect 64800 15570 64846 15576
rect 64800 15566 64834 15570
rect 64722 15542 64824 15566
rect 64914 15542 64948 15910
rect 65418 15706 65452 20092
rect 66162 20058 66200 20062
rect 66162 20024 66202 20058
rect 65594 19990 66202 20024
rect 66172 19984 66174 19990
rect 65562 19951 65572 19952
rect 65521 19940 65572 19951
rect 65418 15682 65488 15706
rect 65532 15682 65572 19940
rect 65418 15610 65436 15682
rect 65520 15644 65578 15682
rect 65590 15650 65600 19980
rect 66200 19956 66202 19990
rect 66206 20040 66240 20092
rect 66842 20062 66844 20066
rect 66206 20024 66252 20040
rect 66820 20024 66858 20062
rect 66964 20040 67002 20062
rect 66952 20024 67010 20040
rect 67478 20024 67516 20062
rect 67582 20030 67610 20092
rect 67638 20030 67666 20050
rect 67722 20040 67760 20062
rect 67710 20024 67768 20040
rect 68136 20024 68174 20062
rect 68480 20040 68518 20062
rect 68468 20024 68526 20040
rect 68794 20024 68832 20062
rect 66206 19990 66858 20024
rect 66910 19990 67516 20024
rect 67568 19990 68174 20024
rect 68226 19990 68832 20024
rect 66206 19952 66252 19990
rect 66952 19952 67010 19990
rect 66179 19940 66194 19951
rect 66206 19940 66240 19952
rect 66868 19951 66888 19952
rect 66837 19940 66888 19951
rect 66190 15706 66240 19940
rect 66848 18680 66888 19940
rect 66190 15682 66246 15706
rect 66848 15682 66882 18680
rect 66964 15706 66998 19952
rect 67495 19940 67540 19951
rect 66958 15694 66998 15706
rect 66958 15682 67004 15694
rect 67506 15682 67540 19940
rect 66178 15644 66230 15682
rect 66256 15644 66286 15650
rect 66836 15644 66894 15682
rect 66936 15650 67004 15682
rect 66902 15644 67004 15650
rect 67494 15644 67552 15682
rect 67582 15650 67610 19984
rect 67638 15650 67666 19984
rect 67710 19952 67768 19990
rect 68468 19952 68526 19990
rect 67722 15694 67756 19952
rect 68153 19940 68198 19951
rect 68164 15682 68198 19940
rect 68480 15694 68514 19952
rect 68811 19940 68856 19951
rect 68822 17388 68856 19940
rect 68936 17388 68970 20092
rect 71336 19970 71696 20108
rect 72232 19970 82586 20108
rect 84631 20428 93069 20464
rect 97126 20428 97160 20554
rect 97240 20428 97274 20462
rect 97898 20428 97932 20462
rect 98012 20428 98046 20554
rect 98316 20428 98350 20554
rect 98430 20428 98464 20462
rect 84631 20394 99060 20428
rect 84631 20007 93069 20394
rect 97126 20326 97160 20394
rect 97228 20326 97406 20364
rect 97420 20326 97944 20364
rect 95942 20292 96610 20326
rect 96700 20292 97406 20326
rect 97458 20292 97944 20326
rect 71336 19936 82586 19970
rect 70964 18180 71286 18232
rect 70884 17810 71286 18180
rect 70964 17724 71286 17810
rect 71336 17670 71696 19936
rect 72232 18278 82586 19936
rect 83798 19462 84160 19828
rect 89024 19524 89050 19600
rect 89052 19524 89078 19628
rect 83706 19314 84160 19462
rect 89024 19402 89050 19426
rect 89052 19402 89078 19426
rect 89212 19402 92178 19992
rect 83798 18772 84160 19314
rect 87508 19150 87528 19350
rect 87536 19122 87556 19378
rect 88308 19310 88856 19344
rect 88308 19028 88342 19310
rect 88670 19230 88681 19241
rect 88366 19108 88370 19230
rect 88372 19186 88444 19224
rect 88494 19196 88681 19230
rect 88682 19186 88754 19224
rect 88394 19136 88398 19186
rect 88410 19152 88444 19186
rect 88670 19142 88681 19153
rect 88720 19152 88754 19186
rect 88494 19108 88681 19142
rect 88822 19028 88856 19310
rect 88308 18994 88856 19028
rect 88906 19054 92178 19402
rect 88906 18940 89544 19054
rect 88262 18666 88276 18752
rect 88300 18628 88314 18790
rect 89096 18564 89098 18940
rect 89124 18592 89126 18940
rect 83782 18448 83786 18560
rect 92724 18558 94374 19996
rect 95832 19994 95842 20148
rect 94810 18556 96460 19994
rect 83816 18448 83820 18526
rect 84690 18490 93038 18524
rect 72232 17670 73728 18278
rect 74968 17786 75002 18278
rect 75082 17938 75127 18278
rect 75414 17926 75459 18278
rect 76172 17926 76217 18278
rect 76930 17926 76975 18278
rect 77688 17926 77733 18278
rect 78446 17926 78491 18278
rect 79204 17926 79249 18278
rect 79962 17926 80007 18278
rect 80140 17938 80185 18278
rect 75106 17888 80150 17926
rect 75144 17854 80150 17888
rect 75402 17838 75460 17854
rect 76160 17838 76218 17854
rect 76918 17838 76976 17854
rect 77676 17838 77734 17854
rect 78434 17838 78492 17854
rect 79192 17838 79250 17854
rect 79950 17838 80008 17854
rect 80254 17786 80288 18278
rect 74968 17752 80288 17786
rect 71626 17442 71660 17670
rect 71690 17580 71700 17588
rect 71718 17524 71756 17588
rect 72268 17442 72302 17670
rect 71348 17408 81696 17442
rect 68764 17348 71264 17388
rect 68822 17332 68856 17348
rect 68936 17332 68970 17348
rect 68708 17292 71320 17332
rect 68822 15682 68856 17292
rect 67694 15644 67732 15682
rect 68152 15644 68210 15682
rect 68452 15644 68490 15682
rect 68810 15644 68868 15682
rect 65520 15622 66230 15644
rect 66252 15622 67004 15644
rect 65520 15610 66224 15622
rect 66252 15610 66258 15622
rect 66268 15610 66974 15622
rect 67026 15610 67732 15644
rect 67784 15610 68490 15644
rect 68542 15610 68868 15644
rect 65418 15542 65452 15610
rect 65520 15594 65578 15610
rect 66178 15594 66224 15610
rect 66836 15594 66894 15610
rect 67494 15594 67552 15610
rect 68152 15594 68210 15610
rect 68810 15594 68868 15610
rect 65520 15579 65535 15594
rect 65532 15542 65566 15576
rect 66190 15542 66224 15594
rect 66848 15542 66882 15576
rect 67506 15542 67540 15594
rect 68853 15579 68868 15594
rect 68164 15542 68198 15576
rect 68822 15542 68856 15576
rect 68936 15542 68970 17292
rect 71348 16756 71382 17408
rect 71512 17328 71546 17408
rect 71626 17328 71660 17408
rect 72268 17328 72302 17408
rect 72382 17328 72416 17408
rect 72428 17328 73128 17339
rect 73140 17328 73174 17408
rect 73186 17328 73886 17339
rect 73898 17328 73932 17408
rect 73944 17328 74546 17339
rect 74656 17328 74690 17408
rect 75414 17328 75448 17408
rect 76172 17328 76206 17408
rect 76930 17328 76964 17408
rect 77688 17328 77722 17408
rect 78446 17328 78480 17408
rect 79204 17328 79238 17408
rect 79628 17328 79950 17339
rect 79962 17328 79996 17408
rect 80008 17328 80542 17339
rect 80720 17328 80754 17408
rect 81478 17328 81512 17408
rect 71512 17306 71660 17328
rect 71412 17278 71484 17304
rect 71506 17294 71660 17306
rect 72234 17294 81512 17328
rect 71506 17282 71546 17294
rect 71412 17266 71490 17278
rect 71450 17198 71490 17266
rect 71450 16954 71484 17198
rect 71450 16898 71490 16954
rect 71478 16886 71490 16898
rect 71478 16882 71484 16886
rect 71500 16882 71546 17282
rect 71506 16870 71546 16882
rect 71626 16870 71660 17294
rect 72268 16870 72302 17294
rect 72316 17288 72376 17294
rect 72382 17282 72416 17294
rect 72422 17288 72496 17294
rect 72428 17282 72429 17283
rect 73127 17282 73128 17283
rect 73140 17282 73174 17294
rect 73186 17282 73187 17283
rect 73885 17282 73886 17283
rect 73898 17282 73932 17294
rect 73944 17282 73945 17283
rect 74643 17282 74644 17283
rect 72382 17281 72428 17282
rect 73128 17281 73129 17282
rect 73140 17281 73186 17282
rect 73886 17281 73887 17282
rect 73898 17281 73944 17282
rect 74644 17281 74645 17282
rect 72382 17278 72427 17281
rect 72344 17260 72376 17278
rect 72382 17260 72468 17278
rect 72382 16883 72427 17260
rect 73140 16883 73185 17281
rect 73898 16883 73943 17281
rect 72382 16882 72428 16883
rect 73128 16882 73129 16883
rect 73140 16882 73186 16883
rect 73886 16882 73887 16883
rect 73898 16882 73944 16883
rect 74644 16882 74645 16883
rect 72382 16870 72416 16882
rect 72428 16881 72429 16882
rect 73127 16881 73128 16882
rect 72428 16870 73128 16881
rect 73140 16870 73174 16882
rect 73186 16881 73187 16882
rect 73885 16881 73886 16882
rect 73186 16870 73886 16881
rect 73898 16870 73932 16882
rect 73944 16881 73945 16882
rect 74643 16881 74644 16882
rect 73944 16870 74546 16881
rect 74656 16870 74690 17294
rect 74702 17282 74703 17283
rect 75401 17282 75402 17283
rect 74701 17281 74702 17282
rect 75402 17281 75403 17282
rect 74701 16882 74702 16883
rect 75402 16882 75403 16883
rect 74702 16881 74703 16882
rect 75401 16881 75402 16882
rect 75414 16870 75448 17294
rect 75460 17282 75461 17283
rect 76159 17282 76160 17283
rect 75459 17281 75460 17282
rect 76160 17281 76161 17282
rect 75459 16882 75460 16883
rect 76160 16882 76161 16883
rect 75460 16881 75461 16882
rect 76159 16881 76160 16882
rect 76172 16870 76206 17294
rect 76858 17288 76924 17294
rect 76218 17282 76219 17283
rect 76917 17282 76918 17283
rect 76217 17281 76218 17282
rect 76918 17281 76919 17282
rect 76886 17260 76924 17270
rect 76217 16882 76218 16883
rect 76918 16882 76919 16883
rect 76218 16881 76219 16882
rect 76917 16881 76918 16882
rect 76930 16870 76964 17294
rect 76970 17288 77038 17294
rect 76976 17282 76977 17283
rect 77675 17282 77676 17283
rect 76975 17281 76976 17282
rect 77676 17281 77677 17282
rect 76970 17260 77010 17270
rect 76975 16882 76976 16883
rect 77676 16882 77677 16883
rect 76976 16881 76977 16882
rect 77675 16881 77676 16882
rect 77688 16870 77722 17294
rect 78374 17288 78440 17294
rect 77734 17282 77735 17283
rect 78433 17282 78434 17283
rect 77733 17281 77734 17282
rect 78434 17281 78435 17282
rect 78402 17260 78440 17278
rect 77733 16882 77734 16883
rect 78434 16882 78435 16883
rect 77734 16881 77735 16882
rect 78433 16881 78434 16882
rect 78446 16870 78480 17294
rect 78486 17288 78554 17294
rect 78492 17282 78493 17283
rect 79191 17282 79192 17283
rect 78491 17281 78492 17282
rect 79192 17281 79193 17282
rect 78486 17260 78526 17278
rect 78491 16882 78492 16883
rect 79192 16882 79193 16883
rect 78492 16881 78493 16882
rect 79191 16881 79192 16882
rect 79204 16870 79238 17294
rect 79896 17288 79956 17294
rect 79250 17282 79251 17283
rect 79949 17282 79950 17283
rect 79962 17282 79996 17294
rect 80002 17288 80076 17294
rect 80008 17282 80009 17283
rect 80707 17282 80708 17283
rect 79249 17281 79250 17282
rect 79950 17281 79951 17282
rect 79962 17281 80008 17282
rect 80708 17281 80709 17282
rect 79962 17280 80007 17281
rect 79924 17260 79956 17280
rect 79962 17260 80048 17280
rect 79962 16883 80007 17260
rect 79249 16882 79250 16883
rect 79950 16882 79951 16883
rect 79962 16882 80008 16883
rect 80708 16882 80709 16883
rect 79250 16881 79251 16882
rect 79949 16881 79950 16882
rect 79628 16870 79950 16881
rect 79962 16870 79996 16882
rect 80008 16881 80009 16882
rect 80707 16881 80708 16882
rect 80008 16870 80542 16881
rect 80720 16870 80754 17294
rect 80766 17282 80767 17283
rect 81465 17282 81466 17283
rect 80765 17281 80766 17282
rect 81466 17281 81467 17282
rect 80765 16882 80766 16883
rect 81466 16882 81467 16883
rect 80766 16881 80767 16882
rect 81465 16881 81466 16882
rect 81478 16870 81512 17294
rect 81524 17282 81594 17304
rect 81522 17278 81594 17282
rect 81522 17266 81600 17278
rect 81522 16882 81524 17266
rect 81560 17198 81600 17266
rect 81618 17226 81628 17306
rect 81560 16954 81616 17198
rect 81560 16898 81600 16954
rect 81590 16886 81600 16898
rect 81618 16926 81644 17226
rect 71506 16858 71660 16870
rect 71512 16836 71660 16858
rect 72234 16836 81512 16870
rect 81618 16858 81628 16926
rect 71512 16756 71546 16836
rect 71626 16756 71660 16836
rect 72268 16756 72302 16836
rect 72382 16756 72416 16836
rect 73140 16756 73174 16836
rect 73898 16756 73932 16836
rect 74656 16756 74690 16836
rect 75414 16756 75448 16836
rect 76172 16756 76206 16836
rect 76930 16756 76964 16836
rect 77688 16756 77722 16836
rect 78446 16756 78480 16836
rect 79204 16756 79238 16836
rect 79962 16756 79996 16836
rect 80720 16756 80754 16836
rect 81478 16756 81512 16836
rect 81662 16756 81696 17408
rect 71348 16722 81696 16756
rect 69232 15682 69278 15706
rect 69990 15682 70036 15706
rect 70748 15682 70794 15706
rect 71506 15694 71546 15706
rect 71506 15682 71552 15694
rect 71626 15604 71660 16722
rect 44832 15508 71564 15542
rect 44832 15472 46467 15508
rect 23857 14958 24272 14989
rect 20304 14953 24272 14958
rect 28928 14958 29349 14989
rect 28928 14953 34288 14958
rect 15233 14919 19069 14953
rect 20304 14924 34288 14953
rect 23857 14919 29349 14924
rect 15613 14867 15624 14878
rect 15636 14867 15647 14878
rect 15137 13153 15171 14857
rect 15613 14851 15647 14867
rect 18655 14851 18689 14889
rect 20684 14872 20695 14883
rect 20707 14872 20718 14883
rect 15313 14817 18989 14851
rect 15251 13153 15285 13187
rect 15613 13153 15647 14817
rect 15716 14758 15772 14769
rect 15898 14758 15954 14769
rect 16374 14758 16430 14769
rect 16556 14758 16612 14769
rect 17032 14758 17088 14769
rect 17214 14758 17270 14769
rect 17690 14758 17735 14769
rect 17872 14758 17917 14769
rect 18348 14758 18393 14769
rect 18530 14758 18575 14769
rect 15727 13153 15772 14758
rect 15788 13153 15816 14434
rect 15909 13153 15954 14758
rect 16385 13153 16430 14758
rect 16446 13153 16474 14434
rect 16502 13153 16530 14434
rect 16567 13153 16612 14758
rect 17043 13153 17088 14758
rect 17108 13153 17136 14434
rect 17164 13153 17192 14434
rect 17225 13153 17270 14758
rect 13841 13119 17297 13153
rect 15137 13051 15171 13119
rect 15251 13082 15298 13098
rect 15239 13070 15298 13082
rect 15239 13057 15319 13070
rect 15239 13051 15298 13057
rect 15613 13051 15647 13119
rect 15727 13116 15772 13119
rect 15727 13098 15761 13116
rect 15788 13098 15816 13119
rect 15909 13116 15954 13119
rect 16385 13116 16430 13119
rect 15909 13098 15943 13116
rect 16385 13098 16419 13116
rect 16446 13098 16474 13119
rect 16502 13113 16530 13119
rect 16567 13116 16612 13119
rect 17043 13116 17088 13119
rect 16502 13098 16531 13113
rect 15727 13051 15774 13098
rect 15788 13051 15852 13098
rect 15909 13067 15956 13098
rect 15897 13051 15956 13067
rect 16385 13051 16432 13098
rect 16446 13057 16531 13098
rect 16567 13098 16601 13116
rect 17043 13098 17077 13116
rect 17108 13098 17136 13119
rect 17164 13098 17192 13119
rect 16567 13067 16614 13098
rect 16446 13051 16510 13057
rect 16555 13051 16614 13067
rect 17043 13051 17090 13098
rect 17108 13051 17192 13098
rect 15137 13017 15163 13051
rect 15167 13017 15171 13024
rect 13859 12850 13893 12958
rect 13825 12622 13848 12822
rect 13853 12594 13893 12850
rect 13859 12450 13893 12594
rect 13825 12222 13848 12422
rect 13853 12194 13893 12450
rect 13859 12050 13893 12194
rect 13825 11822 13848 12022
rect 13853 11794 13893 12050
rect 15137 11944 15171 13017
rect 15239 13017 15852 13051
rect 15895 13017 16510 13051
rect 16553 13017 17192 13051
rect 15239 13011 15297 13017
rect 15175 11944 15205 12974
rect 15239 12970 15319 13011
rect 15251 12726 15291 12970
rect 15245 12424 15291 12726
rect 15296 12424 15319 12970
rect 15245 11944 15319 12424
rect 15613 11944 15647 13017
rect 15727 12424 15761 13017
rect 15771 13011 15817 13017
rect 15771 12670 15816 13011
rect 15844 12983 15845 13017
rect 15897 12970 15955 13017
rect 15827 12969 15844 12970
rect 15822 12958 15867 12969
rect 15827 12670 15867 12958
rect 15833 12424 15867 12670
rect 15909 12424 15943 12970
rect 16385 12424 16419 13017
rect 16429 13011 16475 13017
rect 16502 13011 16503 13017
rect 16429 12424 16474 13011
rect 16502 12970 16531 13011
rect 16555 12970 16613 13017
rect 16485 12969 16531 12970
rect 16480 12958 16531 12969
rect 15727 11944 15772 12424
rect 15833 12126 15878 12424
rect 15812 11944 15882 12126
rect 15909 11944 15954 12424
rect 16385 11944 16474 12424
rect 16485 12424 16530 12958
rect 16567 12424 16601 12970
rect 17043 12424 17077 13017
rect 17087 12640 17136 13017
rect 17164 12970 17192 13017
rect 17143 12969 17192 12970
rect 17138 12958 17192 12969
rect 17143 12640 17192 12958
rect 17225 13116 17297 13119
rect 17149 12424 17183 12640
rect 17225 12424 17259 13116
rect 17263 12424 17297 13116
rect 16485 11944 16536 12424
rect 16567 11944 16612 12424
rect 17043 11944 17088 12424
rect 17149 12104 17194 12424
rect 17134 11944 17204 12104
rect 17225 11944 17297 12424
rect 17701 12424 17735 14758
rect 17701 11944 17746 12424
rect 17778 11944 17806 14434
rect 17834 11944 17862 14434
rect 17883 12424 17917 14758
rect 18359 12424 18393 14758
rect 17883 11944 17928 12424
rect 13859 11650 13893 11794
rect 13825 11422 13848 11622
rect 13853 11394 13893 11650
rect 13859 11250 13893 11394
rect 13825 11022 13848 11222
rect 13853 10994 13893 11250
rect 15096 11910 17990 11944
rect 15096 11112 15130 11910
rect 15137 11112 15171 11910
rect 15175 11799 15205 11910
rect 15245 11892 15319 11910
rect 15245 11876 15291 11892
rect 15238 11848 15291 11876
rect 15296 11848 15319 11892
rect 15613 11889 15647 11910
rect 15727 11892 15772 11910
rect 15727 11889 15761 11892
rect 15238 11842 15285 11848
rect 15613 11842 15660 11889
rect 15727 11842 15774 11889
rect 15812 11842 15882 11910
rect 15909 11892 15954 11910
rect 16385 11892 16474 11910
rect 15909 11876 15943 11892
rect 15896 11842 15943 11876
rect 16385 11889 16419 11892
rect 16429 11889 16474 11892
rect 16385 11848 16474 11889
rect 16485 11892 16536 11910
rect 16567 11892 16612 11910
rect 17043 11892 17088 11910
rect 16485 11889 16530 11892
rect 16485 11848 16538 11889
rect 16567 11876 16601 11892
rect 16385 11842 16432 11848
rect 16491 11842 16538 11848
rect 16554 11842 16601 11876
rect 17043 11889 17077 11892
rect 17043 11842 17090 11889
rect 17134 11842 17204 11910
rect 17225 11892 17297 11910
rect 17225 11876 17259 11892
rect 17212 11842 17259 11876
rect 17263 11889 17297 11892
rect 17701 11892 17746 11910
rect 17701 11889 17735 11892
rect 17263 11842 17310 11889
rect 17701 11842 17748 11889
rect 17778 11848 17806 11910
rect 17834 11904 17862 11910
rect 17834 11889 17882 11904
rect 17814 11848 17882 11889
rect 17883 11892 17928 11910
rect 17778 11842 17861 11848
rect 15251 11808 15882 11842
rect 15251 11802 15285 11808
rect 15175 11223 15209 11799
rect 15210 11761 15244 11765
rect 15245 11761 15291 11802
rect 15210 11262 15291 11761
rect 15210 11257 15244 11262
rect 15251 11248 15291 11262
rect 15175 11112 15205 11223
rect 15238 11220 15291 11248
rect 15296 11220 15319 11802
rect 15613 11261 15647 11808
rect 15727 11261 15761 11808
rect 15812 11765 15882 11808
rect 15909 11808 16538 11842
rect 16567 11808 17204 11842
rect 15812 11754 15902 11765
rect 15909 11754 15943 11808
rect 15812 11670 15943 11754
rect 15833 11578 15943 11670
rect 15833 11318 15867 11578
rect 15771 11261 15816 11318
rect 15238 11214 15285 11220
rect 15613 11214 15660 11261
rect 15727 11220 15816 11261
rect 15827 11261 15867 11318
rect 15868 11261 15902 11578
rect 15827 11257 15902 11261
rect 15827 11220 15880 11257
rect 15909 11248 15943 11578
rect 16046 11442 16342 11504
rect 15727 11214 15774 11220
rect 15833 11214 15880 11220
rect 15896 11214 15943 11248
rect 16385 11261 16419 11808
rect 16491 11802 16525 11808
rect 16429 11261 16474 11802
rect 16385 11220 16474 11261
rect 16485 11765 16530 11802
rect 16485 11257 16560 11765
rect 16485 11220 16538 11257
rect 16567 11248 16601 11808
rect 16385 11214 16432 11220
rect 16491 11214 16538 11220
rect 16554 11214 16601 11248
rect 17043 11261 17077 11808
rect 17134 11765 17204 11808
rect 17225 11808 17861 11842
rect 17134 11736 17218 11765
rect 17225 11736 17259 11808
rect 17134 11648 17259 11736
rect 17149 11594 17259 11648
rect 17149 11288 17183 11594
rect 17184 11288 17218 11594
rect 17087 11261 17136 11288
rect 17043 11220 17136 11261
rect 17143 11257 17218 11288
rect 17225 11470 17259 11594
rect 17263 11470 17297 11808
rect 17390 11470 17686 11504
rect 17701 11470 17735 11808
rect 17778 11802 17826 11808
rect 17834 11802 17854 11808
rect 17778 11470 17806 11802
rect 17834 11760 17882 11802
rect 17831 11749 17882 11760
rect 17834 11470 17876 11749
rect 17883 11470 17917 11892
rect 17956 11470 17990 11910
rect 18359 11892 18404 12424
rect 17225 11430 18082 11470
rect 17225 11414 17259 11430
rect 17263 11414 17297 11430
rect 17701 11414 17735 11430
rect 17772 11414 17806 11430
rect 17834 11414 17876 11430
rect 17883 11414 17917 11430
rect 17956 11414 17990 11430
rect 17225 11402 18026 11414
rect 17225 11374 17446 11402
rect 17630 11374 18026 11402
rect 17143 11220 17196 11257
rect 17225 11248 17259 11374
rect 17043 11214 17090 11220
rect 17149 11214 17196 11220
rect 17212 11214 17259 11248
rect 17263 11261 17297 11374
rect 17701 11261 17735 11374
rect 17794 11268 17806 11374
rect 17822 11273 17876 11374
rect 17822 11272 17882 11273
rect 17828 11268 17882 11272
rect 17263 11214 17310 11261
rect 17701 11214 17748 11261
rect 17772 11220 17806 11268
rect 17834 11261 17882 11268
rect 17814 11220 17882 11261
rect 17772 11214 17861 11220
rect 15251 11180 15880 11214
rect 15909 11180 16538 11214
rect 16567 11180 17196 11214
rect 17225 11180 17861 11214
rect 15251 11174 15285 11180
rect 15251 11112 15291 11174
rect 15296 11112 15319 11174
rect 15613 11112 15647 11180
rect 15727 11112 15761 11180
rect 15833 11174 15867 11180
rect 15771 11112 15816 11174
rect 15827 11112 15867 11174
rect 15909 11112 15943 11180
rect 16385 11112 16419 11180
rect 16491 11174 16525 11180
rect 16429 11112 16474 11174
rect 16485 11112 16530 11174
rect 16567 11112 16601 11180
rect 17043 11112 17077 11180
rect 17149 11174 17183 11180
rect 17087 11112 17136 11174
rect 17143 11112 17192 11174
rect 17225 11112 17259 11180
rect 17263 11112 17297 11180
rect 17701 11112 17735 11180
rect 17778 11174 17826 11180
rect 17834 11174 17854 11180
rect 17778 11112 17806 11174
rect 17834 11118 17882 11174
rect 17834 11112 17862 11118
rect 17883 11112 17917 11374
rect 17956 11112 17990 11374
rect 15096 11078 17990 11112
rect 13859 10850 13893 10994
rect 13825 10622 13848 10822
rect 13853 10594 13893 10850
rect 13859 10450 13893 10594
rect 13825 10222 13848 10422
rect 13853 10194 13893 10450
rect 15137 10236 15171 11078
rect 15175 10236 15205 11078
rect 15251 10236 15291 11078
rect 15296 10236 15319 11078
rect 15613 10236 15647 11078
rect 15727 10236 15761 11078
rect 15771 10236 15816 11078
rect 15827 10236 15867 11078
rect 15909 10236 15943 11078
rect 15946 10952 16158 10960
rect 15946 10512 16358 10952
rect 16146 10504 16358 10512
rect 13859 9758 13893 10194
rect 13825 9530 13848 9730
rect 13853 9622 13893 9758
rect 14074 10202 16310 10236
rect 13853 9502 13876 9622
rect 14074 9160 14108 10202
rect 15137 10181 15171 10202
rect 15175 10181 15205 10202
rect 15251 10181 15291 10202
rect 15296 10181 15319 10202
rect 15613 10181 15647 10202
rect 15727 10181 15761 10202
rect 15771 10181 15816 10202
rect 14517 10150 14564 10181
rect 14505 10134 14564 10150
rect 14818 10134 14865 10181
rect 15137 10134 15222 10181
rect 15251 10140 15319 10181
rect 15251 10134 15298 10140
rect 15476 10134 15523 10181
rect 15613 10134 15660 10181
rect 15727 10140 15816 10181
rect 15827 10181 15867 10202
rect 15909 10181 15943 10202
rect 15827 10140 15880 10181
rect 15727 10134 15774 10140
rect 15833 10134 15880 10140
rect 15909 10134 15956 10181
rect 16134 10134 16181 10181
rect 14250 10100 14865 10134
rect 14908 10100 15523 10134
rect 15566 10100 16181 10134
rect 14505 10053 14563 10100
rect 15137 10053 15221 10100
rect 14177 10041 14222 10052
rect 14188 9296 14222 10041
rect 14168 9160 14244 9296
rect 14074 9006 14290 9160
rect 14517 9053 14551 10053
rect 14835 10041 14880 10052
rect 14846 9065 14880 10041
rect 15137 9053 15171 10053
rect 15175 9053 15209 10053
rect 15251 9053 15285 10100
rect 15493 10041 15538 10052
rect 15504 9328 15538 10041
rect 15482 9160 15562 9328
rect 14505 9006 14564 9053
rect 14818 9006 14865 9053
rect 15137 9006 15222 9053
rect 15251 9006 15298 9053
rect 15400 9006 15612 9160
rect 15613 9053 15647 10100
rect 15727 9053 15761 10100
rect 15833 9053 15867 10100
rect 15909 9053 15943 10100
rect 16151 10041 16196 10052
rect 16162 9065 16196 10041
rect 15613 9006 15660 9053
rect 15727 9006 15774 9053
rect 15833 9006 15880 9053
rect 15909 9006 15956 9053
rect 16134 9006 16181 9053
rect 14074 8972 14865 9006
rect 14908 8972 16181 9006
rect 14074 8904 14290 8972
rect 14505 8956 14563 8972
rect 15137 8956 15221 8972
rect 15251 8966 15285 8972
rect 15137 8904 15171 8956
rect 15175 8904 15205 8956
rect 15251 8904 15291 8966
rect 15296 8904 15319 8966
rect 15400 8904 15612 8972
rect 15613 8904 15647 8972
rect 15727 8904 15761 8972
rect 15833 8966 15867 8972
rect 15771 8904 15816 8966
rect 15827 8904 15867 8966
rect 15909 8904 15943 8972
rect 16276 8904 16310 10202
rect 14074 8870 16310 8904
rect 14078 8712 14290 8870
rect 14062 7266 15054 8686
rect 15137 8564 15171 8870
rect 15175 8564 15205 8870
rect 15251 8686 15291 8870
rect 15296 8686 15319 8870
rect 15400 8712 15612 8870
rect 15613 8686 15647 8870
rect 15727 8686 15761 8870
rect 15771 8686 15816 8870
rect 15827 8686 15867 8870
rect 15909 8686 15943 8870
rect 15251 8610 16244 8686
rect 15137 8468 15215 8564
rect 15245 8508 16244 8610
rect 15132 8228 15215 8468
rect 15100 8122 15110 8228
rect 15137 8098 15215 8228
rect 15132 8060 15215 8098
rect 15137 7342 15215 8060
rect 14517 6432 14551 7266
rect 15137 6621 15171 7342
rect 15175 7078 15215 7342
rect 15218 7106 15243 8508
rect 15251 7266 16244 8508
rect 15251 7106 15296 7266
rect 15175 6621 15205 7078
rect 15251 6782 15319 7106
rect 15268 6770 15291 6782
rect 15296 6770 15319 6782
rect 15613 6770 15647 7266
rect 15727 7166 15816 7266
rect 15827 7166 15878 7266
rect 15727 6828 15772 7166
rect 15833 6828 15878 7166
rect 15727 6782 15816 6828
rect 15771 6770 15816 6782
rect 15827 6770 15878 6828
rect 15909 6782 15954 7266
rect 16385 6782 16419 11078
rect 15266 6723 16254 6770
rect 16429 6729 16474 11078
rect 16485 6770 16530 11078
rect 16567 8694 16601 11078
rect 16792 10952 17004 10960
rect 16622 10512 17004 10952
rect 16622 10504 16834 10512
rect 17043 10242 17077 11078
rect 17087 10242 17136 11078
rect 17143 10242 17192 11078
rect 17225 10242 17259 11078
rect 17263 10242 17297 11078
rect 17476 10952 17480 10960
rect 17488 10512 17492 10952
rect 17701 10242 17735 11078
rect 17778 10242 17806 11078
rect 17834 10242 17862 11078
rect 17883 10242 17917 11078
rect 17964 10504 18346 10952
rect 18359 10242 18393 11892
rect 18430 10622 18458 11908
rect 18486 10242 18514 14434
rect 18541 12424 18575 14758
rect 18541 11892 18586 12424
rect 18655 11948 18689 14817
rect 18780 13158 19201 13194
rect 20208 13158 20242 14862
rect 20684 14856 20718 14872
rect 22848 14862 22876 14882
rect 22904 14862 22932 14882
rect 23556 14862 23584 14882
rect 23726 14856 23760 14903
rect 20684 14822 23760 14856
rect 20322 13158 20356 13192
rect 20684 13158 20718 14822
rect 20787 14772 20832 14783
rect 20969 14772 21025 14783
rect 21445 14772 21501 14783
rect 21627 14772 21683 14783
rect 22103 14772 22159 14783
rect 22285 14772 22341 14783
rect 22761 14772 22817 14783
rect 20798 13158 20832 14772
rect 20874 14032 20902 14434
rect 20980 14336 21025 14772
rect 21456 14424 21501 14772
rect 21526 14424 21554 14434
rect 21582 14424 21610 14434
rect 21638 14424 21683 14772
rect 22114 14424 22159 14772
rect 22184 14424 22212 14434
rect 22240 14424 22268 14434
rect 22296 14424 22341 14772
rect 22772 14424 22817 14772
rect 22848 14424 22876 14816
rect 22904 14424 22932 14816
rect 22943 14772 22999 14783
rect 23419 14772 23475 14783
rect 22954 14424 22999 14772
rect 23430 14424 23475 14772
rect 23556 14424 23584 14816
rect 23601 14772 23657 14783
rect 23612 14424 23657 14772
rect 23726 14424 23760 14822
rect 23857 14424 24272 14919
rect 20942 13848 20948 13854
rect 20874 13158 20902 13832
rect 20980 13158 21014 14336
rect 21128 13486 24272 14424
rect 25761 14867 25772 14878
rect 25784 14867 25795 14878
rect 25761 14851 25795 14867
rect 27411 14851 27445 14889
rect 28928 14851 29349 14919
rect 25761 14817 27445 14851
rect 28450 14817 28479 14851
rect 25761 14392 25795 14817
rect 25864 14758 25920 14769
rect 25970 14758 26026 14769
rect 26522 14758 26578 14769
rect 26628 14758 26684 14769
rect 27180 14758 27236 14769
rect 27286 14758 27342 14769
rect 25875 14392 25920 14758
rect 25932 14392 25943 14470
rect 25981 14392 26026 14758
rect 24676 14358 26254 14392
rect 21456 13158 21490 13486
rect 21526 13158 21554 13486
rect 21582 13158 21610 13486
rect 21638 13158 21672 13486
rect 22114 13158 22148 13486
rect 22184 13158 22212 13486
rect 22240 13158 22268 13486
rect 22296 13158 22330 13486
rect 18780 13124 22368 13158
rect 18780 11984 19201 13124
rect 20208 13056 20242 13124
rect 20344 13094 20362 13122
rect 20322 13087 20362 13094
rect 20310 13072 20362 13087
rect 20310 13056 20368 13072
rect 20372 13062 20390 13094
rect 20684 13056 20718 13124
rect 20798 13094 20832 13124
rect 20874 13094 20902 13124
rect 20980 13094 21014 13124
rect 21456 13094 21490 13124
rect 21526 13094 21554 13124
rect 20798 13056 20836 13094
rect 20874 13056 20914 13094
rect 20980 13072 21018 13094
rect 20968 13056 21026 13072
rect 21456 13056 21494 13094
rect 21526 13056 21572 13094
rect 20208 13022 20234 13056
rect 20238 13022 20242 13038
rect 20174 12716 20180 12768
rect 20208 12716 20242 13022
rect 20310 13022 20914 13056
rect 20966 13022 21572 13056
rect 20246 12716 20276 12988
rect 20310 12984 20368 13022
rect 20316 12716 20362 12984
rect 20372 12716 20390 13016
rect 20684 12716 20718 13022
rect 20798 12716 20832 13022
rect 20874 12984 20902 13022
rect 20968 12984 21026 13022
rect 20893 12972 20938 12983
rect 20904 12716 20938 12972
rect 20980 12716 21014 12984
rect 21456 12716 21490 13022
rect 21500 12983 21554 13022
rect 21582 12984 21610 13124
rect 21638 13094 21672 13124
rect 22114 13094 22148 13124
rect 22184 13094 22212 13124
rect 21638 13072 21676 13094
rect 21626 13056 21684 13072
rect 22114 13056 22152 13094
rect 22184 13056 22230 13094
rect 21624 13022 22230 13056
rect 21626 12984 21684 13022
rect 21556 12983 21610 12984
rect 21500 12972 21610 12983
rect 21500 12716 21554 12972
rect 21556 12716 21610 12972
rect 21638 12716 21672 12984
rect 22114 12716 22148 13022
rect 22158 12983 22212 13022
rect 22240 12984 22268 13124
rect 22214 12983 22268 12984
rect 22158 12972 22268 12983
rect 22158 12716 22212 12972
rect 22214 12716 22268 12972
rect 22296 12716 22330 13124
rect 22334 12716 22368 13124
rect 22772 12722 22806 13486
rect 22848 12722 22876 13486
rect 22904 12722 22932 13486
rect 22954 12722 22988 13486
rect 23430 12722 23464 13486
rect 23500 13032 23528 13486
rect 23556 12722 23584 13486
rect 23612 12722 23646 13486
rect 23726 12722 23760 13486
rect 23857 12722 24272 13486
rect 24622 13112 24628 14248
rect 24676 13060 24710 14358
rect 25444 14337 25488 14352
rect 25323 14306 25370 14337
rect 24726 13452 24750 14296
rect 25311 14290 25370 14306
rect 25420 14296 25488 14337
rect 25761 14337 25795 14358
rect 25875 14337 25920 14358
rect 25388 14290 25467 14296
rect 25761 14290 25808 14337
rect 25875 14290 25922 14337
rect 25932 14296 25943 14358
rect 25981 14337 26026 14358
rect 25981 14290 26028 14337
rect 26078 14290 26125 14337
rect 24852 14256 25467 14290
rect 25510 14256 26125 14290
rect 25311 14250 25432 14256
rect 25311 14209 25386 14250
rect 25444 14222 25460 14256
rect 24779 14197 24824 14208
rect 24790 14044 24824 14197
rect 25323 14044 25357 14209
rect 25364 14204 25386 14209
rect 25437 14204 25482 14208
rect 25420 14197 25482 14204
rect 24790 13221 24835 14044
rect 24726 13122 24750 13212
rect 25323 13209 25368 14044
rect 25420 13936 25442 14197
rect 25448 14044 25482 14197
rect 25448 13221 25493 14044
rect 25761 13209 25795 14256
rect 25875 14044 25909 14256
rect 25981 14044 26015 14256
rect 26095 14197 26140 14208
rect 26106 14044 26140 14197
rect 25875 13254 25920 14044
rect 25981 13254 26026 14044
rect 25832 13209 26026 13254
rect 26106 13221 26151 14044
rect 24805 13162 26125 13209
rect 24852 13128 25467 13162
rect 25510 13128 26125 13162
rect 25311 13112 25369 13128
rect 25388 13122 25432 13128
rect 25444 13122 25460 13128
rect 25323 13104 25357 13112
rect 25444 13104 25488 13122
rect 25761 13104 25795 13128
rect 25875 13104 25920 13128
rect 25932 13118 25943 13122
rect 25981 13104 26026 13128
rect 26220 13104 26254 14358
rect 26533 14350 26578 14758
rect 26639 14520 26684 14758
rect 26605 14350 26618 14464
rect 26533 14336 26618 14350
rect 26533 14044 26567 14336
rect 26577 14044 26618 14336
rect 26533 13112 26618 14044
rect 26633 14336 26684 14520
rect 27191 14390 27236 14758
rect 27254 14390 27259 14440
rect 27297 14390 27342 14758
rect 27411 14390 27445 14817
rect 28488 14779 28517 14846
rect 28569 14817 29349 14851
rect 26762 14356 28340 14390
rect 26633 14044 26674 14336
rect 26533 13104 26578 13112
rect 26633 13104 26684 14044
rect 26762 13104 26796 14356
rect 27191 14336 27236 14356
rect 27191 14335 27225 14336
rect 27226 14335 27231 14336
rect 27191 14288 27238 14335
rect 27254 14294 27259 14356
rect 27297 14336 27342 14356
rect 27297 14335 27331 14336
rect 27411 14335 27445 14356
rect 27297 14288 27344 14335
rect 27411 14288 27458 14335
rect 27506 14288 27553 14335
rect 27849 14304 27896 14335
rect 27837 14288 27896 14304
rect 28164 14288 28211 14335
rect 26938 14254 27553 14288
rect 27596 14254 28211 14288
rect 26865 14195 26910 14206
rect 26876 14044 26910 14195
rect 27191 14044 27225 14254
rect 27297 14044 27331 14254
rect 26876 13219 26921 14044
rect 27191 13856 27236 14044
rect 27297 13904 27342 14044
rect 27282 13856 27352 13904
rect 27100 13702 27352 13856
rect 27191 13207 27236 13702
rect 27282 13448 27352 13702
rect 27297 13207 27342 13448
rect 27411 13207 27445 14254
rect 27837 14207 27895 14254
rect 27523 14195 27568 14206
rect 27534 14044 27568 14195
rect 27849 14044 27883 14207
rect 28181 14195 28226 14206
rect 28192 14044 28226 14195
rect 27534 13219 27579 14044
rect 27849 13926 27894 14044
rect 27828 13852 27898 13926
rect 27748 13706 27998 13852
rect 27828 13470 27898 13706
rect 27849 13207 27894 13470
rect 28192 13219 28237 14044
rect 26891 13160 28211 13207
rect 26938 13126 27553 13160
rect 27596 13126 28211 13160
rect 24770 13070 27090 13104
rect 24770 13060 24804 13070
rect 25444 13066 25488 13070
rect 25761 13060 25795 13070
rect 25875 13060 25920 13070
rect 25981 13060 26026 13070
rect 26220 13060 26254 13070
rect 24676 13026 26254 13060
rect 26533 13049 26578 13070
rect 26633 13056 26684 13070
rect 26639 13049 26684 13056
rect 26762 13058 26796 13070
rect 27056 13058 27090 13070
rect 27191 13058 27236 13126
rect 27254 13088 27259 13120
rect 27297 13058 27342 13126
rect 27411 13058 27445 13126
rect 27837 13110 27895 13126
rect 28306 13058 28340 14356
rect 20106 11984 22414 12716
rect 18780 11948 22414 11984
rect 18608 11914 22414 11948
rect 18541 11452 18575 11892
rect 18608 11452 18642 11914
rect 18655 11452 18689 11914
rect 18722 11764 18723 11769
rect 18711 11753 18756 11764
rect 18722 11452 18756 11753
rect 18780 11452 22414 11914
rect 18541 11430 22414 11452
rect 18541 11424 18575 11430
rect 18608 11424 18642 11430
rect 18655 11424 18689 11430
rect 18722 11424 18756 11430
rect 18780 11424 22414 11430
rect 18541 11374 22414 11424
rect 18541 10242 18575 11374
rect 18608 10952 18642 11374
rect 18655 10990 18689 11374
rect 18722 10990 18756 11374
rect 18780 11278 22414 11374
rect 22684 12686 24272 12722
rect 24770 12686 24804 13026
rect 25323 13018 25370 13026
rect 25311 13002 25370 13018
rect 25761 13002 25795 13026
rect 25875 13002 25922 13026
rect 25981 13018 26028 13026
rect 25969 13002 26028 13018
rect 26533 13002 26580 13049
rect 26639 13018 26686 13049
rect 26762 13024 28340 13058
rect 26627 13002 26686 13018
rect 26914 13002 26961 13024
rect 24930 12992 26961 13002
rect 24946 12968 26961 12992
rect 25311 12921 25369 12968
rect 24873 12909 24918 12920
rect 24884 12766 24918 12909
rect 24884 12686 24929 12766
rect 22684 12652 24956 12686
rect 22684 12584 24272 12652
rect 24770 12631 24804 12652
rect 24665 12600 24712 12631
rect 24653 12584 24712 12600
rect 24770 12584 24817 12631
rect 22684 12550 24817 12584
rect 22684 12088 24272 12550
rect 24653 12503 24711 12550
rect 24770 12544 24804 12550
rect 24665 12424 24699 12503
rect 22684 12034 24612 12088
rect 22684 12032 24272 12034
rect 22684 12006 24612 12032
rect 22684 11948 24272 12006
rect 24665 11948 24710 12424
rect 24726 11948 24750 12544
rect 24770 12502 24806 12544
rect 24808 12502 24838 12507
rect 24770 12491 24842 12502
rect 24770 11948 24806 12491
rect 24808 12424 24842 12491
rect 24808 11948 24853 12424
rect 24884 11948 24956 12652
rect 25323 12424 25357 12921
rect 25323 11948 25368 12424
rect 25761 11948 25795 12968
rect 25875 12424 25909 12968
rect 25969 12921 26027 12968
rect 25981 12424 26015 12921
rect 25875 11948 25920 12424
rect 25981 11948 26026 12424
rect 22684 11914 26350 11948
rect 22684 11503 24272 11914
rect 24665 11893 24710 11914
rect 24665 11862 24712 11893
rect 24653 11846 24712 11862
rect 24726 11852 24750 11914
rect 24770 11893 24806 11914
rect 24808 11893 24853 11914
rect 24884 11893 24956 11914
rect 25323 11893 25368 11914
rect 25761 11893 25795 11914
rect 25875 11893 25920 11914
rect 25981 11893 26026 11914
rect 24770 11846 24855 11893
rect 24858 11846 25284 11893
rect 25323 11846 25370 11893
rect 25516 11846 25563 11893
rect 25761 11846 25808 11893
rect 25875 11846 25922 11893
rect 25981 11846 26028 11893
rect 26174 11846 26221 11893
rect 24290 11812 25563 11846
rect 25606 11812 26221 11846
rect 24653 11765 24711 11812
rect 24665 11503 24699 11765
rect 24770 11503 24804 11812
rect 24808 11515 24842 11812
rect 24808 11503 24838 11515
rect 22684 11456 24283 11503
rect 24665 11456 24712 11503
rect 24770 11499 24838 11503
rect 24770 11456 24817 11499
rect 22684 11422 24817 11456
rect 22684 11354 24272 11422
rect 24665 11354 24699 11422
rect 24770 11354 24804 11422
rect 24884 11354 24956 11812
rect 22684 11320 24956 11354
rect 22684 11284 24272 11320
rect 18780 11094 20276 11278
rect 20316 11240 20362 11278
rect 20372 11240 20390 11278
rect 20322 11094 20356 11240
rect 20658 11094 22330 11278
rect 18780 11060 22330 11094
rect 18655 10952 18772 10990
rect 18780 10952 20280 11060
rect 20322 11044 20356 11060
rect 20362 11044 20372 11054
rect 20316 11026 20362 11044
rect 20308 10998 20362 11026
rect 20372 10998 20390 11044
rect 20308 10992 20356 10998
rect 20362 10992 20372 10998
rect 20658 10992 22330 11060
rect 20322 10958 22330 10992
rect 20322 10952 20356 10958
rect 18608 10908 20280 10952
rect 20288 10908 20314 10924
rect 18608 10826 20314 10908
rect 18608 10582 20242 10826
rect 18610 10546 20242 10582
rect 18610 10504 19201 10546
rect 18655 10242 18689 10504
rect 18780 10242 19201 10504
rect 16652 10208 19201 10242
rect 19388 10262 19422 10546
rect 19502 10414 19536 10546
rect 19588 10414 19624 10546
rect 19634 10414 19635 10546
rect 19588 10402 19622 10414
rect 19502 10286 19510 10400
rect 19576 10380 19578 10402
rect 19580 10380 19622 10402
rect 19530 10314 19538 10372
rect 19576 10364 19622 10380
rect 19546 10330 19622 10364
rect 19576 10314 19622 10330
rect 19588 10262 19622 10314
rect 19704 10262 19738 10546
rect 19388 10228 19738 10262
rect 19864 10262 19898 10546
rect 19978 10414 20012 10546
rect 20066 10414 20100 10546
rect 20056 10364 20094 10402
rect 20022 10330 20094 10364
rect 20166 10262 20242 10546
rect 19864 10228 20242 10262
rect 16652 8910 16686 10208
rect 17043 10187 17077 10208
rect 17087 10187 17136 10208
rect 17043 10146 17136 10187
rect 17143 10187 17192 10208
rect 17225 10187 17259 10208
rect 17263 10187 17297 10208
rect 17701 10187 17735 10208
rect 17143 10146 17196 10187
rect 17043 10140 17090 10146
rect 17149 10140 17196 10146
rect 17225 10140 17310 10187
rect 17396 10140 17443 10187
rect 17701 10140 17748 10187
rect 17778 10146 17806 10208
rect 17834 10146 17862 10208
rect 17883 10187 17917 10208
rect 18359 10187 18393 10208
rect 17883 10140 17930 10187
rect 18054 10140 18101 10187
rect 18359 10140 18406 10187
rect 18486 10146 18514 10208
rect 18541 10187 18575 10208
rect 18655 10187 18689 10208
rect 18541 10140 18588 10187
rect 18655 10140 18702 10187
rect 18712 10140 18759 10187
rect 16828 10106 17443 10140
rect 17486 10106 18101 10140
rect 18144 10106 18759 10140
rect 16755 10047 16800 10058
rect 16766 9340 16800 10047
rect 16740 9152 16822 9340
rect 16740 9076 16954 9152
rect 16742 9012 16954 9076
rect 17043 9059 17077 10106
rect 17149 9059 17183 10106
rect 17225 9059 17259 10106
rect 17263 9059 17297 10106
rect 17413 10047 17458 10058
rect 17424 9071 17458 10047
rect 17701 9059 17735 10106
rect 17883 9059 17917 10106
rect 18071 10047 18116 10058
rect 18082 9818 18116 10047
rect 18359 9818 18393 10106
rect 18541 9818 18575 10106
rect 18082 9628 18127 9818
rect 18359 9628 18404 9818
rect 17974 9596 18404 9628
rect 18541 9596 18586 9818
rect 18610 9638 18613 9720
rect 17974 9594 18393 9596
rect 17974 9096 18008 9594
rect 18082 9449 18116 9594
rect 18188 9526 18235 9573
rect 18134 9492 18235 9526
rect 18330 9566 18393 9594
rect 18082 9433 18127 9449
rect 18205 9433 18250 9444
rect 18082 9330 18122 9433
rect 18054 9198 18144 9330
rect 18216 9257 18250 9433
rect 18188 9198 18235 9245
rect 18054 9164 18235 9198
rect 18054 9124 18214 9164
rect 18330 9158 18398 9566
rect 18054 9096 18144 9124
rect 18330 9096 18393 9158
rect 17974 9062 18393 9096
rect 18359 9059 18393 9062
rect 18541 9059 18575 9596
rect 18655 9059 18689 10106
rect 18729 10047 18774 10058
rect 18740 9071 18774 10047
rect 17043 9012 17090 9059
rect 17149 9012 17196 9059
rect 17225 9012 17310 9059
rect 17396 9012 17443 9059
rect 17701 9012 17748 9059
rect 17883 9012 17930 9059
rect 18054 9012 18101 9059
rect 18359 9012 18406 9059
rect 18541 9012 18588 9059
rect 18655 9012 18702 9059
rect 18712 9012 18759 9059
rect 16742 8978 17443 9012
rect 17486 8978 18759 9012
rect 16742 8910 16954 8978
rect 17043 8910 17077 8978
rect 17149 8972 17183 8978
rect 17087 8910 17136 8972
rect 17143 8910 17192 8972
rect 17225 8910 17259 8978
rect 17263 8910 17297 8978
rect 17701 8910 17735 8978
rect 17883 8910 17917 8978
rect 17960 8910 18393 8978
rect 18486 8910 18514 8972
rect 18541 8910 18575 8978
rect 18655 8910 18689 8978
rect 18780 8910 19201 10208
rect 20166 9780 20200 10228
rect 20208 9780 20242 10228
rect 20246 10268 20314 10826
rect 20316 10598 20362 10952
rect 20372 10598 20390 10952
rect 20658 10932 22330 10958
rect 20322 10404 20356 10598
rect 20566 10544 22330 10932
rect 20566 10500 20778 10544
rect 20798 10500 20832 10544
rect 20316 10268 20362 10404
rect 20246 10050 20367 10268
rect 20246 9932 20314 10050
rect 20246 9780 20280 9932
rect 20288 9916 20314 9932
rect 20316 9916 20362 10050
rect 20308 9888 20362 9916
rect 20372 9888 20390 10404
rect 20422 10376 20850 10500
rect 20684 9920 20718 10376
rect 20798 9920 20832 10376
rect 20308 9882 20356 9888
rect 20684 9882 20722 9920
rect 20798 9882 20836 9920
rect 20904 9916 20972 10544
rect 20904 9882 20944 9916
rect 20322 9848 20944 9882
rect 20322 9842 20356 9848
rect 20316 9796 20362 9842
rect 20316 9780 20367 9796
rect 20372 9780 20390 9842
rect 20684 9780 20718 9848
rect 20798 9796 20832 9848
rect 20904 9796 20938 9848
rect 20980 9796 21014 10544
rect 21042 10484 21444 10544
rect 20798 9780 20843 9796
rect 20904 9780 20949 9796
rect 20980 9780 21025 9796
rect 21052 9780 21086 10484
rect 21098 10102 21136 10484
rect 21158 10162 21196 10484
rect 21232 10480 21444 10484
rect 20166 9746 21086 9780
rect 21356 9780 21390 10480
rect 21456 9916 21554 10544
rect 21456 9784 21490 9916
rect 21500 9888 21554 9916
rect 21556 10496 21610 10544
rect 21638 10496 21672 10544
rect 21708 10496 22092 10544
rect 21556 10484 22092 10496
rect 21556 10372 22024 10484
rect 21556 9888 21610 10372
rect 21638 9920 21672 10372
rect 22114 10254 22212 10544
rect 22214 10254 22276 10544
rect 22114 9944 22162 10254
rect 22220 9944 22276 10254
rect 22114 9920 22212 9944
rect 21562 9882 21600 9888
rect 21638 9882 21676 9920
rect 22100 9916 22212 9920
rect 22100 9882 22148 9916
rect 21516 9848 21524 9882
rect 21532 9848 22148 9882
rect 21562 9842 21596 9848
rect 21500 9784 21554 9842
rect 21456 9780 21554 9784
rect 21556 9780 21610 9842
rect 21638 9784 21672 9848
rect 22114 9784 22148 9848
rect 22158 9784 22212 9916
rect 21638 9780 21683 9784
rect 22114 9780 22212 9784
rect 22214 9780 22276 9944
rect 21356 9746 22276 9780
rect 16652 8876 19201 8910
rect 16742 8704 16954 8876
rect 17043 8694 17077 8876
rect 17087 8694 17136 8876
rect 17143 8694 17192 8876
rect 17225 8694 17259 8876
rect 17263 8694 17297 8876
rect 17701 8702 17735 8876
rect 17760 8702 17806 8876
rect 17816 8702 17862 8876
rect 17883 8702 17917 8876
rect 17960 8702 18393 8876
rect 18486 8798 18514 8876
rect 18541 8702 18575 8876
rect 18655 8702 18689 8876
rect 16562 6770 17554 8694
rect 16479 6723 16537 6770
rect 16548 6723 17554 6770
rect 17701 6766 18722 8702
rect 17730 6758 18722 6766
rect 17720 6732 18722 6758
rect 17730 6723 18722 6732
rect 18780 8670 19201 8876
rect 20208 8670 20242 9746
rect 20246 8670 20276 9746
rect 20316 8670 20367 9746
rect 20372 8670 20390 9746
rect 20684 8670 20718 9746
rect 20760 9278 20794 9550
rect 20798 8670 20843 9746
rect 20904 8670 20949 9746
rect 20980 8670 21025 9746
rect 21456 8670 21554 9746
rect 21556 8670 21610 9746
rect 21620 9308 21634 9546
rect 21638 8670 21683 9746
rect 22114 8670 22212 9746
rect 22214 8670 22268 9746
rect 22296 8670 22330 10544
rect 22334 10932 22368 11278
rect 22762 11146 24272 11284
rect 24665 11146 24699 11320
rect 24770 11146 24804 11320
rect 22762 11102 24804 11146
rect 22666 11068 24804 11102
rect 22334 10926 22568 10932
rect 22666 10926 22700 11068
rect 22334 10922 22760 10926
rect 22762 10922 24804 11068
rect 24884 11258 24931 11320
rect 24884 10952 24920 11258
rect 25323 11150 25357 11812
rect 25533 11753 25578 11764
rect 25544 11150 25578 11753
rect 25761 11150 25795 11812
rect 25875 11150 25909 11812
rect 25981 11150 26015 11812
rect 26191 11753 26236 11764
rect 26202 11150 26236 11753
rect 26316 11150 26350 11914
rect 26533 11150 26567 12968
rect 26627 12921 26685 12968
rect 26639 11150 26673 12921
rect 26931 12909 26976 12920
rect 26942 11150 26976 12909
rect 27056 11150 27090 13024
rect 27191 11150 27225 13024
rect 27297 11150 27331 13024
rect 27411 11150 27445 13024
rect 28507 11968 28541 14758
rect 28928 14428 29349 14817
rect 30832 14872 30843 14883
rect 30855 14872 30866 14883
rect 30832 14856 30866 14872
rect 32482 14856 32516 14903
rect 30832 14822 32516 14856
rect 30832 14428 30866 14822
rect 30935 14772 30991 14783
rect 31041 14772 31097 14783
rect 31593 14772 31649 14783
rect 31699 14772 31755 14783
rect 32251 14772 32307 14783
rect 32357 14772 32413 14783
rect 30946 14428 30991 14772
rect 31052 14428 31097 14772
rect 31604 14428 31649 14772
rect 31710 14428 31755 14772
rect 32262 14428 32307 14772
rect 32368 14428 32413 14772
rect 28928 14392 32454 14428
rect 28866 14358 32454 14392
rect 28866 11968 28900 14358
rect 28928 11968 32454 14358
rect 28330 11932 32454 11968
rect 32482 11932 32516 14822
rect 32920 11932 32954 11966
rect 33578 11932 33624 11966
rect 28330 11898 33686 11932
rect 28330 11830 32454 11898
rect 32482 11830 32516 11898
rect 32920 11846 32958 11868
rect 32908 11830 32966 11846
rect 33026 11830 33548 11868
rect 28330 11796 33548 11830
rect 28330 11428 32454 11796
rect 28122 11394 32454 11428
rect 28122 11150 28156 11394
rect 28330 11326 32454 11394
rect 28298 11292 32454 11326
rect 28225 11233 28270 11244
rect 28236 11150 28270 11233
rect 28330 11150 32454 11292
rect 24958 10952 32454 11150
rect 24884 10933 32454 10952
rect 22334 10772 24804 10922
rect 24886 10920 32454 10933
rect 32482 10920 32516 11796
rect 32908 11758 32966 11796
rect 32920 10958 32954 11758
rect 33527 11746 33566 11757
rect 33476 10972 33500 11118
rect 33504 11000 33528 11090
rect 33538 10970 33572 11746
rect 32908 10920 32966 10958
rect 33026 10920 33548 10958
rect 33578 10932 33610 11784
rect 24886 10886 33548 10920
rect 24886 10818 32454 10886
rect 32482 10818 32516 10886
rect 32908 10870 32966 10886
rect 32920 10818 32954 10852
rect 33578 10818 33624 10852
rect 33652 10818 33686 11898
rect 24886 10784 33686 10818
rect 24886 10772 32454 10784
rect 22334 10748 32454 10772
rect 22334 10738 28582 10748
rect 22334 10710 24790 10738
rect 22334 10484 22760 10710
rect 22334 8670 22368 10484
rect 22548 10478 22760 10484
rect 22762 10510 24790 10710
rect 24886 10510 28582 10738
rect 28758 10510 32454 10748
rect 22666 9188 22700 10478
rect 22762 10474 32454 10510
rect 32482 10474 32516 10784
rect 32920 10474 32954 10508
rect 33578 10474 33612 10508
rect 34236 10474 34270 10508
rect 34350 10474 34384 14862
rect 42356 13039 45830 13278
rect 45868 13039 46467 13282
rect 55352 13189 55386 15508
rect 57440 15112 57474 15508
rect 56998 14874 57712 15112
rect 56990 14554 57712 14874
rect 56990 14502 57694 14554
rect 57440 13189 57474 14502
rect 53910 13028 53944 13046
rect 42646 12398 42680 12892
rect 48992 12626 49010 12802
rect 44652 12532 44708 12550
rect 44652 12486 44708 12514
rect 44940 12486 45236 12548
rect 42760 12398 42794 12432
rect 42436 12364 42906 12398
rect 45382 12372 45434 12442
rect 42646 12156 42680 12364
rect 42748 12318 42777 12350
rect 42712 12305 42777 12318
rect 42712 12294 42751 12305
rect 42712 12266 42723 12290
rect 42806 12246 42842 12258
rect 42786 12238 42842 12246
rect 42772 12234 42842 12238
rect 42772 12194 42804 12234
rect 42806 12224 42842 12234
rect 42770 12168 42804 12194
rect 42872 12156 42906 12364
rect 45266 12316 45434 12372
rect 45266 12236 45402 12316
rect 42646 12122 42723 12156
rect 42736 12134 45444 12156
rect 42742 12122 45444 12134
rect 42872 12104 42906 12122
rect 47656 11836 47660 12160
rect 46210 11812 46336 11836
rect 46266 11809 46312 11812
rect 46924 11809 46970 11836
rect 47552 11812 47660 11836
rect 47582 11809 47628 11812
rect 46182 11784 46364 11808
rect 46238 11781 46340 11784
rect 46896 11781 46998 11808
rect 47524 11784 47688 11808
rect 47554 11781 47656 11784
rect 49754 11658 49776 12936
rect 49788 11658 49810 12936
rect 50488 12298 51480 13028
rect 51678 12298 52670 13028
rect 52988 12360 53944 13028
rect 54336 12712 54346 13070
rect 54336 12498 54364 12712
rect 54336 12492 54346 12498
rect 52988 12290 53936 12360
rect 51120 12114 51154 12148
rect 51778 12114 51812 12148
rect 52436 12114 52470 12148
rect 50500 12080 52736 12114
rect 53752 12108 53786 12142
rect 53866 12108 53900 12290
rect 54479 12282 55148 13189
rect 55244 12414 55250 12664
rect 54515 12108 54549 12282
rect 55316 12278 58103 13189
rect 58870 12410 58904 15508
rect 60311 15472 63935 15508
rect 64598 15492 64632 15508
rect 64914 15492 64948 15508
rect 60347 13402 60381 15472
rect 59320 13368 62776 13402
rect 59996 13194 60030 13223
rect 60032 13194 60036 13219
rect 60347 13194 60381 13368
rect 60461 13331 60508 13347
rect 60449 13300 60508 13331
rect 60626 13300 60673 13347
rect 61119 13316 61166 13347
rect 61107 13300 61166 13316
rect 61284 13300 61331 13347
rect 61777 13316 61824 13347
rect 61765 13300 61824 13316
rect 61942 13300 61989 13347
rect 62435 13316 62482 13347
rect 62423 13300 62482 13316
rect 62600 13300 62647 13347
rect 60449 13266 60673 13300
rect 60716 13266 61331 13300
rect 61374 13266 61989 13300
rect 62032 13266 62647 13300
rect 60449 13219 60507 13266
rect 60461 13194 60495 13219
rect 60654 13218 60688 13223
rect 61107 13219 61165 13266
rect 60643 13207 60688 13218
rect 60654 13194 60688 13207
rect 61119 13194 61153 13219
rect 61312 13218 61346 13223
rect 61765 13219 61823 13266
rect 61301 13207 61346 13218
rect 61312 13194 61346 13207
rect 61777 13194 61811 13219
rect 61970 13218 62004 13223
rect 62423 13219 62481 13266
rect 61959 13207 62004 13218
rect 61970 13194 62004 13207
rect 62435 13194 62469 13219
rect 62540 13194 62562 13260
rect 62568 13218 62618 13260
rect 62628 13218 62662 13223
rect 62568 13207 62662 13218
rect 62568 13194 62618 13207
rect 62628 13194 62662 13207
rect 62742 13194 62776 13368
rect 54629 12108 54663 12142
rect 50466 12018 50496 12052
rect 46122 11590 46472 11592
rect 22762 10440 34998 10474
rect 22762 10360 32454 10440
rect 32482 10360 32516 10440
rect 32920 10360 32954 10440
rect 33026 10360 33566 10371
rect 33578 10360 33612 10440
rect 33624 10360 33940 10371
rect 34236 10360 34270 10440
rect 34350 10360 34384 10440
rect 22762 10326 34384 10360
rect 22762 9990 32454 10326
rect 22762 9902 29349 9990
rect 29724 9914 29725 9915
rect 29723 9913 29724 9914
rect 29736 9902 29770 9990
rect 29781 9914 29782 9915
rect 30382 9914 30383 9915
rect 29782 9913 29783 9914
rect 30381 9913 30382 9914
rect 30394 9902 30428 9990
rect 30439 9914 30440 9915
rect 30440 9913 30441 9914
rect 30832 9902 30866 9990
rect 30946 9902 30980 9990
rect 31052 9902 31086 9990
rect 31604 9902 31638 9990
rect 31710 9902 31744 9990
rect 32262 9902 32296 9990
rect 32368 9902 32402 9990
rect 32482 9902 32516 10326
rect 32907 10314 32908 10315
rect 32908 10313 32909 10314
rect 32908 9914 32909 9915
rect 32907 9913 32908 9914
rect 32920 9902 32954 10326
rect 32966 10314 32967 10315
rect 33565 10314 33566 10315
rect 33578 10314 33612 10326
rect 33624 10314 33625 10315
rect 34223 10314 34224 10315
rect 32965 10313 32966 10314
rect 33566 10313 33567 10314
rect 33578 10313 33624 10314
rect 34224 10313 34225 10314
rect 33578 9915 33623 10313
rect 32965 9914 32966 9915
rect 33566 9914 33567 9915
rect 33578 9914 33624 9915
rect 34224 9914 34225 9915
rect 32966 9913 32967 9914
rect 33565 9913 33566 9914
rect 33026 9902 33566 9913
rect 33578 9902 33612 9914
rect 33624 9913 33625 9914
rect 34223 9913 34224 9914
rect 33624 9902 33940 9913
rect 34236 9902 34270 10326
rect 34350 9902 34384 10326
rect 22762 9868 34384 9902
rect 41588 9878 43896 11316
rect 44166 9884 46472 11322
rect 50348 11014 50382 11140
rect 50428 10866 50452 11122
rect 50456 10838 50480 11150
rect 50500 10782 50534 12080
rect 51120 12028 51167 12059
rect 51108 12012 51167 12028
rect 51244 12012 51291 12059
rect 51778 12028 51825 12059
rect 51766 12012 51825 12028
rect 51902 12012 51949 12059
rect 52436 12028 52483 12059
rect 52424 12012 52483 12028
rect 52560 12012 52607 12059
rect 50676 11978 51291 12012
rect 51334 11978 51949 12012
rect 51992 11978 52607 12012
rect 51108 11931 51166 11978
rect 51766 11972 51824 11978
rect 51766 11931 51864 11972
rect 50603 11919 50648 11930
rect 50614 11466 50648 11919
rect 50614 11408 51006 11466
rect 51120 11408 51154 11931
rect 51261 11919 51306 11930
rect 50614 11304 51180 11408
rect 50614 11302 51006 11304
rect 50614 10943 50648 11302
rect 51120 10931 51154 11304
rect 51272 10943 51306 11919
rect 51392 11408 51584 11450
rect 51778 11408 51864 11931
rect 51392 11336 51864 11408
rect 51502 11302 51864 11336
rect 51778 10931 51864 11302
rect 51108 10884 51167 10931
rect 51244 10884 51291 10931
rect 51766 10890 51864 10931
rect 51868 11930 51920 11972
rect 52424 11931 52482 11978
rect 51868 11919 51964 11930
rect 51868 10931 51920 11919
rect 51930 10943 51964 11919
rect 52036 11406 52228 11456
rect 52436 11406 52470 11931
rect 52036 11342 52470 11406
rect 52160 11300 52470 11342
rect 52436 10931 52470 11300
rect 51868 10890 51949 10931
rect 51766 10884 51825 10890
rect 51902 10884 51949 10890
rect 52424 10884 52483 10931
rect 52512 10890 52524 11972
rect 52540 11930 52580 11972
rect 52540 11919 52622 11930
rect 52540 10931 52580 11919
rect 52588 10943 52622 11919
rect 52540 10890 52607 10931
rect 52560 10884 52607 10890
rect 50676 10850 51291 10884
rect 51334 10850 51949 10884
rect 51992 10850 52607 10884
rect 51108 10834 51166 10850
rect 51766 10834 51824 10850
rect 52424 10834 52482 10850
rect 51120 10782 51154 10816
rect 51778 10782 51812 10816
rect 52436 10782 52470 10816
rect 52702 10782 52736 12080
rect 50500 10748 52736 10782
rect 53078 12074 55314 12108
rect 53078 12046 53112 12074
rect 53078 10838 53146 12046
rect 53752 12022 53798 12053
rect 53740 12006 53798 12022
rect 53254 11972 53798 12006
rect 53832 11972 53838 12006
rect 53740 11925 53798 11972
rect 53156 11622 53162 11918
rect 53181 11913 53226 11924
rect 53192 10937 53226 11913
rect 53332 11388 53524 11440
rect 53752 11388 53786 11925
rect 53308 11320 53786 11388
rect 53752 10925 53786 11320
rect 53788 11140 53820 11504
rect 53844 11140 53848 11925
rect 53788 10930 53848 11140
rect 53788 10925 53820 10930
rect 53844 10925 53848 10930
rect 53740 10878 53820 10925
rect 53254 10844 53798 10878
rect 53078 10776 53112 10838
rect 53740 10828 53820 10844
rect 53754 10813 53820 10828
rect 53754 10810 53786 10813
rect 53752 10776 53786 10810
rect 53788 10776 53820 10813
rect 53866 10776 53900 12074
rect 54481 11972 54496 12006
rect 54515 10776 54549 12074
rect 54629 12037 54676 12053
rect 54617 12006 54676 12037
rect 55138 12006 55185 12053
rect 54554 11972 54587 12006
rect 54617 11972 55185 12006
rect 55280 12046 55314 12074
rect 54617 11925 54675 11972
rect 54629 11504 54663 11925
rect 55155 11913 55200 11924
rect 55166 11504 55200 11913
rect 54629 10925 54674 11504
rect 55166 10937 55211 11504
rect 54570 10844 54587 10878
rect 54617 10844 55185 10925
rect 54617 10828 54675 10844
rect 55280 10838 55348 12046
rect 54617 10813 54632 10828
rect 54629 10776 54663 10810
rect 55280 10776 55314 10838
rect 53078 10742 55314 10776
rect 53754 10294 53786 10742
rect 53788 10328 53820 10742
rect 51778 9906 51812 9940
rect 52436 9906 52470 9940
rect 53094 9906 53128 9940
rect 53752 9906 53786 9940
rect 53866 9906 53900 10742
rect 54515 10196 54549 10742
rect 55287 10402 55321 10436
rect 55945 10402 55979 10436
rect 57261 10404 57295 10438
rect 57919 10404 57953 10438
rect 58033 10404 58067 12278
rect 59550 11891 63174 13194
rect 65418 13189 65452 15508
rect 67506 13189 67540 15508
rect 64799 12990 64802 13016
rect 64827 13011 64830 13044
rect 59550 11857 63185 11891
rect 59550 11719 63174 11857
rect 65382 11742 68251 13189
rect 68854 11952 68862 12180
rect 68882 11952 68890 12152
rect 68936 11874 68970 15508
rect 72268 13864 72302 16722
rect 84690 16684 84724 18490
rect 85132 18416 85158 18474
rect 85160 18416 85186 18446
rect 85268 18410 85302 18490
rect 86026 18410 86060 18490
rect 86784 18410 86818 18490
rect 87542 18410 87576 18490
rect 88300 18410 88334 18490
rect 89058 18410 89092 18490
rect 89816 18410 89850 18490
rect 90574 18410 90608 18490
rect 91332 18410 91366 18490
rect 92090 18410 92124 18490
rect 92848 18410 92882 18490
rect 84876 18388 92882 18410
rect 84876 18386 92888 18388
rect 84754 18348 84826 18386
rect 84876 18376 92936 18386
rect 84792 17780 84826 18348
rect 85132 18310 85158 18370
rect 85160 18338 85186 18370
rect 85255 18364 85256 18365
rect 85256 18363 85257 18364
rect 85256 17764 85257 17765
rect 85255 17763 85256 17764
rect 85268 17752 85302 18376
rect 85314 18364 85315 18365
rect 86013 18364 86014 18365
rect 85313 18363 85314 18364
rect 86014 18363 86015 18364
rect 85313 17764 85314 17765
rect 86014 17764 86015 17765
rect 85314 17763 85315 17764
rect 86013 17763 86014 17764
rect 86026 17752 86060 18376
rect 86072 18364 86073 18365
rect 86771 18364 86772 18365
rect 86071 18363 86072 18364
rect 86772 18363 86773 18364
rect 86071 17764 86072 17765
rect 86772 17764 86773 17765
rect 86072 17763 86073 17764
rect 86771 17763 86772 17764
rect 86784 17752 86818 18376
rect 86830 18364 86831 18365
rect 87529 18364 87530 18365
rect 86829 18363 86830 18364
rect 87530 18363 87531 18364
rect 86829 17764 86830 17765
rect 87530 17764 87531 17765
rect 86830 17763 86831 17764
rect 87529 17763 87530 17764
rect 87542 17752 87576 18376
rect 87588 18364 87589 18365
rect 88287 18364 88288 18365
rect 87587 18363 87588 18364
rect 88288 18363 88289 18364
rect 88300 18284 88334 18376
rect 88346 18364 88347 18365
rect 89045 18364 89046 18365
rect 88345 18363 88346 18364
rect 89046 18363 89047 18364
rect 89058 18284 89092 18376
rect 89104 18364 89105 18365
rect 89803 18364 89804 18365
rect 89103 18363 89104 18364
rect 89804 18363 89805 18364
rect 89816 18284 89850 18376
rect 89862 18364 89863 18365
rect 90561 18364 90562 18365
rect 89861 18363 89862 18364
rect 90562 18363 90563 18364
rect 87770 17884 88148 18112
rect 87587 17764 87588 17765
rect 87588 17763 87589 17764
rect 87770 17763 88092 17884
rect 88190 17763 90498 18284
rect 90562 17764 90563 17765
rect 90561 17763 90562 17764
rect 87770 17752 90498 17763
rect 90574 17752 90608 18376
rect 90620 18364 90621 18365
rect 91319 18364 91320 18365
rect 90619 18363 90620 18364
rect 91320 18363 91321 18364
rect 91332 18290 91366 18376
rect 91378 18364 91379 18365
rect 92077 18364 92078 18365
rect 91377 18363 91378 18364
rect 92078 18363 92079 18364
rect 92090 18290 92124 18376
rect 92136 18364 92137 18365
rect 92835 18364 92836 18365
rect 92135 18363 92136 18364
rect 92836 18363 92837 18364
rect 92848 18348 92936 18376
rect 92848 18290 92894 18348
rect 92896 18290 92936 18348
rect 92990 18290 93002 18306
rect 93004 18290 93038 18490
rect 90619 17764 90620 17765
rect 90620 17763 90621 17764
rect 90768 17752 93076 18290
rect 84754 17690 84826 17728
rect 84876 17718 93076 17752
rect 85255 17706 85256 17707
rect 85256 17705 85257 17706
rect 84792 17122 84826 17690
rect 85138 17100 85158 17164
rect 85166 17100 85186 17136
rect 85256 17106 85257 17107
rect 85255 17105 85256 17106
rect 85268 17094 85302 17718
rect 85314 17706 85315 17707
rect 86013 17706 86014 17707
rect 85313 17705 85314 17706
rect 86014 17705 86015 17706
rect 85313 17106 85314 17107
rect 86014 17106 86015 17107
rect 85314 17105 85315 17106
rect 86013 17105 86014 17106
rect 86026 17094 86060 17718
rect 86072 17706 86073 17707
rect 86771 17706 86772 17707
rect 86071 17705 86072 17706
rect 86772 17705 86773 17706
rect 86071 17106 86072 17107
rect 86772 17106 86773 17107
rect 86072 17105 86073 17106
rect 86771 17105 86772 17106
rect 86784 17094 86818 17718
rect 86830 17706 86831 17707
rect 87529 17706 87530 17707
rect 86829 17705 86830 17706
rect 87530 17705 87531 17706
rect 86829 17106 86830 17107
rect 87530 17106 87531 17107
rect 86830 17105 86831 17106
rect 87529 17105 87530 17106
rect 87542 17094 87576 17718
rect 87588 17706 87589 17707
rect 87587 17705 87588 17706
rect 87816 17556 87984 17718
rect 87587 17106 87588 17107
rect 87588 17105 87589 17106
rect 88190 17105 90498 17718
rect 90561 17706 90562 17707
rect 90562 17705 90563 17706
rect 87896 17094 90498 17105
rect 90524 17100 90532 17178
rect 90562 17106 90563 17107
rect 90561 17105 90562 17106
rect 90574 17094 90608 17718
rect 90620 17706 90621 17707
rect 90619 17705 90620 17706
rect 90619 17106 90620 17107
rect 90620 17105 90621 17106
rect 90768 17094 93076 17718
rect 84754 17032 84826 17070
rect 84876 17060 93076 17094
rect 84792 16688 84826 17032
rect 85138 17000 85158 17054
rect 85166 17028 85186 17054
rect 85255 17048 85256 17049
rect 85256 17047 85257 17048
rect 84754 16684 84826 16688
rect 85268 16684 85302 17060
rect 85314 17048 85315 17049
rect 86013 17048 86014 17049
rect 85313 17047 85314 17048
rect 86014 17047 86015 17048
rect 86026 16684 86060 17060
rect 86072 17048 86073 17049
rect 86771 17048 86772 17049
rect 86071 17047 86072 17048
rect 86772 17047 86773 17048
rect 86784 16684 86818 17060
rect 86830 17048 86831 17049
rect 87529 17048 87530 17049
rect 86829 17047 86830 17048
rect 87530 17047 87531 17048
rect 87542 16684 87576 17060
rect 87588 17048 87589 17049
rect 87587 17047 87588 17048
rect 88190 16846 90498 17060
rect 90524 16978 90532 17054
rect 90561 17048 90562 17049
rect 90562 17047 90563 17048
rect 88300 16684 88334 16846
rect 89058 16684 89092 16846
rect 89816 16684 89850 16846
rect 90574 16684 90608 17060
rect 90620 17048 90621 17049
rect 90619 17047 90620 17048
rect 90768 16852 93076 17060
rect 91332 16684 91366 16852
rect 92090 16684 92124 16852
rect 92848 16688 92894 16852
rect 92902 16688 92936 16852
rect 92848 16684 92936 16688
rect 92962 16684 92974 16852
rect 92990 16684 93002 16852
rect 93004 16684 93038 16852
rect 96638 16684 96672 20242
rect 97126 19996 97160 20292
rect 97228 20254 97286 20292
rect 97886 20254 97944 20292
rect 97240 19996 97285 20254
rect 97385 20242 97441 20253
rect 97396 19996 97441 20242
rect 97898 19996 97943 20254
rect 98012 19996 98046 20394
rect 98316 19996 98350 20394
rect 98418 20292 98922 20364
rect 99026 20332 99060 20394
rect 98418 20254 98476 20292
rect 98430 19996 98475 20254
rect 98901 20242 98957 20253
rect 98912 19996 98957 20242
rect 99026 20142 99078 20332
rect 99026 19996 99060 20142
rect 99088 19996 99094 20366
rect 104042 20157 104076 22644
rect 116196 21314 116222 21402
rect 106598 20162 106632 20191
rect 107256 20162 107290 20191
rect 107914 20162 107948 20191
rect 108572 20162 108606 20191
rect 109230 20162 109264 20191
rect 117278 20164 117312 20180
rect 100512 19996 100546 20014
rect 96914 19266 99272 19996
rect 99590 19328 100546 19996
rect 100938 19680 100948 20038
rect 100938 19466 100966 19680
rect 100938 19460 100948 19466
rect 96914 19082 99096 19266
rect 99590 19258 100538 19328
rect 96914 19048 99338 19082
rect 100354 19076 100388 19110
rect 100468 19076 100502 19258
rect 101081 19250 101750 20157
rect 101846 19382 101852 19632
rect 101117 19076 101151 19250
rect 101918 19246 104705 20157
rect 101231 19076 101265 19110
rect 96914 18980 99096 19048
rect 99162 18980 99209 19027
rect 96914 18946 99209 18980
rect 96852 18276 96860 18288
rect 96864 18238 96872 18276
rect 96914 18108 99096 18946
rect 96878 17982 99096 18108
rect 96914 17852 99096 17982
rect 99114 17858 99126 18940
rect 99142 18898 99182 18940
rect 99142 18887 99224 18898
rect 99142 17899 99182 18887
rect 99190 17911 99224 18887
rect 99142 17858 99209 17899
rect 99162 17852 99209 17858
rect 96914 17818 99209 17852
rect 96914 17750 99096 17818
rect 99304 17750 99338 19048
rect 96914 17716 99338 17750
rect 99680 19042 101916 19076
rect 99680 19014 99714 19042
rect 99680 17806 99748 19014
rect 99809 18974 100400 19021
rect 99856 18940 100400 18974
rect 100342 18893 100400 18940
rect 99758 18590 99764 18886
rect 99783 18881 99839 18892
rect 99794 17905 99839 18881
rect 99934 18356 100126 18408
rect 100354 18356 100399 18893
rect 99910 18288 100399 18356
rect 100354 17893 100399 18288
rect 100446 18108 100450 18893
rect 100420 17898 100450 18108
rect 100446 17893 100450 17898
rect 99809 17846 100400 17893
rect 99856 17812 100400 17846
rect 99680 17744 99714 17806
rect 100342 17796 100400 17812
rect 100385 17781 100400 17796
rect 100354 17744 100388 17778
rect 100468 17744 100502 19042
rect 101117 17744 101151 19042
rect 101172 18940 101189 18974
rect 101219 18940 101787 19021
rect 101882 19014 101916 19042
rect 101219 18893 101277 18940
rect 101231 17893 101276 18893
rect 101757 18881 101813 18892
rect 101768 17905 101813 18881
rect 101172 17812 101189 17846
rect 101219 17812 101787 17893
rect 101219 17796 101277 17812
rect 101882 17806 101950 19014
rect 101219 17781 101234 17796
rect 101231 17744 101265 17778
rect 101882 17744 101916 17806
rect 96714 16684 96720 17286
rect 96914 16874 99096 17716
rect 99680 17710 101916 17744
rect 99696 16874 99730 16908
rect 100354 16874 100388 16908
rect 100468 16874 100502 17710
rect 101117 17164 101151 17710
rect 101231 17164 101265 17710
rect 101889 17370 101923 17404
rect 102547 17370 102581 17404
rect 103863 17372 103897 17406
rect 104521 17372 104555 17406
rect 104635 17372 104669 19246
rect 101636 17336 103214 17370
rect 96914 16840 100922 16874
rect 96914 16772 99096 16840
rect 99518 16772 100400 16819
rect 96914 16738 99573 16772
rect 99616 16738 100231 16772
rect 100274 16738 100400 16772
rect 96914 16684 99096 16738
rect 99684 16732 99742 16738
rect 100342 16732 100400 16738
rect 99590 16690 99638 16732
rect 72370 16650 99096 16684
rect 99543 16679 99638 16690
rect 72382 16620 72416 16650
rect 73140 16620 73174 16650
rect 73898 16620 73932 16650
rect 74656 16620 74690 16650
rect 75414 16620 75448 16650
rect 76172 16620 76206 16650
rect 76930 16620 76964 16650
rect 77688 16620 77722 16650
rect 78446 16620 78480 16650
rect 79204 16620 79238 16650
rect 79962 16620 79996 16650
rect 80720 16620 80754 16650
rect 81478 16620 81512 16650
rect 82236 16620 82270 16650
rect 82994 16620 83028 16650
rect 83752 16620 83786 16650
rect 72382 16582 81636 16620
rect 82208 16616 82270 16620
rect 82208 16588 82276 16616
rect 82202 16582 82276 16588
rect 82286 16582 82304 16588
rect 82966 16582 83028 16620
rect 83724 16582 83786 16620
rect 83816 16620 83820 16650
rect 84510 16620 84544 16650
rect 84690 16620 84724 16650
rect 83816 16582 84728 16620
rect 84792 16582 84826 16650
rect 85268 16620 85302 16650
rect 86026 16620 86060 16650
rect 86784 16620 86818 16650
rect 87542 16620 87576 16650
rect 85240 16582 85302 16620
rect 85998 16582 86060 16620
rect 86756 16582 86818 16620
rect 87514 16582 87576 16620
rect 88250 16628 89170 16650
rect 88250 16620 88284 16628
rect 88300 16620 88334 16628
rect 89058 16620 89092 16628
rect 88250 16582 88334 16620
rect 89030 16582 89092 16620
rect 89136 16582 89170 16628
rect 89440 16628 90360 16650
rect 89440 16582 89474 16628
rect 89816 16620 89850 16628
rect 89788 16582 89850 16620
rect 89862 16582 89878 16598
rect 90326 16582 90360 16628
rect 90574 16620 90608 16650
rect 90546 16582 90608 16620
rect 90750 16636 91670 16650
rect 90750 16582 90784 16636
rect 91332 16620 91366 16636
rect 91304 16606 91366 16620
rect 91304 16582 91370 16606
rect 72382 15706 72416 16582
rect 72444 16548 73180 16582
rect 73106 16542 73124 16548
rect 73134 16514 73180 16548
rect 73190 16548 73932 16582
rect 73960 16548 74696 16582
rect 73190 16542 73208 16548
rect 72376 15682 72422 15706
rect 73140 15682 73174 16514
rect 73898 15682 73932 16548
rect 74622 16542 74640 16548
rect 74650 16514 74696 16548
rect 74706 16548 75448 16582
rect 75476 16548 76212 16582
rect 74706 16542 74724 16548
rect 74656 15682 74690 16514
rect 75414 15682 75448 16548
rect 76138 16542 76156 16548
rect 76166 16514 76212 16548
rect 76222 16548 76964 16582
rect 76992 16548 77728 16582
rect 76222 16542 76240 16548
rect 76172 15682 76206 16514
rect 76930 15706 76964 16548
rect 77654 16542 77672 16548
rect 77682 16514 77728 16548
rect 77738 16548 78480 16582
rect 78508 16548 79244 16582
rect 77738 16542 77756 16548
rect 76924 15682 76970 15706
rect 77688 15682 77722 16514
rect 78446 15706 78480 16548
rect 79170 16542 79188 16548
rect 79198 16514 79244 16548
rect 79254 16548 79996 16582
rect 80024 16548 80760 16582
rect 79254 16542 79272 16548
rect 72376 15644 74546 15682
rect 74628 15644 74690 15682
rect 75386 15678 75448 15682
rect 75386 15650 75454 15678
rect 75380 15644 75454 15650
rect 75464 15644 75482 15650
rect 76144 15644 76206 15682
rect 76902 15650 76970 15682
rect 76896 15644 76970 15650
rect 76980 15644 76998 15650
rect 77660 15644 77722 15682
rect 77808 15650 77824 15704
rect 78440 15682 78486 15706
rect 79204 15682 79238 16514
rect 79962 15706 79996 16548
rect 80686 16542 80704 16548
rect 80714 16514 80760 16548
rect 80770 16548 81512 16582
rect 81540 16548 82276 16582
rect 82282 16548 83028 16582
rect 83040 16548 83786 16582
rect 83798 16548 84544 16582
rect 84572 16548 85302 16582
rect 85314 16548 86060 16582
rect 86072 16548 86818 16582
rect 86830 16548 87576 16582
rect 87588 16566 88334 16582
rect 87588 16548 88288 16566
rect 80770 16542 80788 16548
rect 79956 15682 80002 15706
rect 80720 15682 80754 16514
rect 81478 15706 81512 16548
rect 82202 16542 82220 16548
rect 82230 16514 82276 16548
rect 82286 16542 82304 16548
rect 81472 15682 81518 15706
rect 82236 15682 82270 16514
rect 82994 15706 83028 16548
rect 82988 15682 83034 15706
rect 83752 15682 83786 16548
rect 78418 15650 78486 15682
rect 78412 15644 78486 15650
rect 78496 15644 78514 15650
rect 79176 15644 79238 15682
rect 79628 15644 80542 15682
rect 80692 15644 80754 15682
rect 81450 15650 81518 15682
rect 81444 15644 81518 15650
rect 81528 15644 81546 15650
rect 82208 15644 82270 15682
rect 82966 15650 83034 15682
rect 82960 15644 83034 15650
rect 83044 15644 83062 15650
rect 83724 15644 83786 15682
rect 83816 15682 83820 16548
rect 84510 15706 84544 16548
rect 84504 15682 84550 15706
rect 84690 15682 84724 16548
rect 84792 16464 84826 16548
rect 85256 16448 85257 16449
rect 85255 16447 85256 16448
rect 85268 16436 85302 16548
rect 85313 16448 85314 16449
rect 86014 16448 86015 16449
rect 85314 16447 85315 16448
rect 86013 16447 86014 16448
rect 86026 16436 86060 16548
rect 86071 16448 86072 16449
rect 86772 16448 86773 16449
rect 86072 16447 86073 16448
rect 86771 16447 86772 16448
rect 86784 16436 86818 16548
rect 86829 16448 86830 16449
rect 87530 16448 87531 16449
rect 86830 16447 86831 16448
rect 87529 16447 87530 16448
rect 87542 16436 87576 16548
rect 87587 16448 87588 16449
rect 87588 16447 87589 16448
rect 88250 16436 88284 16548
rect 88300 16516 88334 16566
rect 88346 16548 89092 16582
rect 89104 16560 89854 16582
rect 89862 16560 90608 16582
rect 89104 16548 90608 16560
rect 90620 16568 91370 16582
rect 91378 16582 91394 16606
rect 91636 16582 91670 16636
rect 91918 16644 92838 16650
rect 91918 16582 91952 16644
rect 92090 16620 92124 16644
rect 92062 16610 92124 16620
rect 92060 16598 92124 16610
rect 92136 16598 92152 16614
rect 92052 16582 92172 16598
rect 92804 16582 92838 16644
rect 91378 16568 92838 16582
rect 90620 16548 92838 16568
rect 88426 16526 89032 16548
rect 88300 16486 88340 16516
rect 88436 16510 88444 16514
rect 88364 16488 88368 16492
rect 88358 16487 88368 16488
rect 88288 16448 88289 16449
rect 88287 16447 88288 16448
rect 88300 16436 88334 16486
rect 88353 16476 88398 16487
rect 88345 16448 88346 16449
rect 88346 16447 88347 16448
rect 88364 16436 88398 16476
rect 88408 16482 88416 16486
rect 88408 16442 88418 16482
rect 88436 16442 88446 16510
rect 89024 16487 89056 16492
rect 89011 16476 89056 16487
rect 89022 16436 89056 16476
rect 89058 16436 89092 16548
rect 89103 16448 89104 16449
rect 89104 16447 89105 16448
rect 89136 16436 89170 16548
rect 89440 16436 89474 16548
rect 89616 16526 90222 16548
rect 89543 16476 89588 16487
rect 89554 16436 89588 16476
rect 89816 16436 89850 16526
rect 90201 16476 90246 16487
rect 90212 16436 90246 16476
rect 90326 16436 90360 16548
rect 90524 16442 90532 16520
rect 90562 16448 90563 16449
rect 90561 16447 90562 16448
rect 90574 16436 90608 16548
rect 90619 16448 90620 16449
rect 90620 16447 90621 16448
rect 90750 16436 90784 16548
rect 90926 16534 91532 16548
rect 90853 16484 90898 16495
rect 90864 16436 90898 16484
rect 91332 16436 91366 16534
rect 91462 16520 91472 16532
rect 91444 16476 91462 16520
rect 91472 16495 91518 16520
rect 91472 16484 91556 16495
rect 91472 16476 91518 16484
rect 91522 16436 91556 16484
rect 91636 16436 91670 16548
rect 91918 16520 92050 16548
rect 92052 16542 92700 16548
rect 91918 16476 91976 16520
rect 92026 16503 92050 16504
rect 92052 16503 92172 16542
rect 92021 16498 92172 16503
rect 91986 16476 92172 16498
rect 92679 16492 92724 16503
rect 91918 16436 91952 16476
rect 92002 16450 92172 16476
rect 92002 16436 92078 16450
rect 92090 16436 92124 16450
rect 92690 16436 92724 16492
rect 92804 16436 92838 16548
rect 92848 16582 92894 16650
rect 92902 16582 92936 16650
rect 92962 16588 92974 16650
rect 92990 16588 93002 16650
rect 93004 16582 93038 16650
rect 93078 16648 96630 16650
rect 93078 16582 93112 16648
rect 93578 16618 93616 16620
rect 93630 16618 93640 16620
rect 94336 16618 94374 16620
rect 94388 16618 94398 16620
rect 95094 16618 95132 16620
rect 95146 16618 95156 16620
rect 95298 16618 95890 16620
rect 95904 16618 96378 16620
rect 93578 16596 93644 16618
rect 93652 16596 93668 16618
rect 93578 16582 93668 16596
rect 94336 16596 94402 16618
rect 94410 16596 94426 16618
rect 94336 16582 94426 16596
rect 95094 16614 95160 16618
rect 95094 16582 95172 16614
rect 95298 16582 96378 16618
rect 96596 16582 96630 16648
rect 92848 16548 96630 16582
rect 92848 16448 92894 16548
rect 92902 16542 92936 16548
rect 92902 16520 92974 16542
rect 92896 16464 92942 16520
rect 92990 16496 93002 16542
rect 92896 16452 92916 16464
rect 92934 16452 92942 16464
rect 92902 16448 92916 16452
rect 92848 16436 92888 16448
rect 84876 16424 92888 16436
rect 84876 16414 92882 16424
rect 84876 16412 92888 16414
rect 84754 16374 84826 16412
rect 84876 16402 92936 16412
rect 85192 16396 85262 16402
rect 85255 16390 85256 16391
rect 85256 16389 85257 16390
rect 84792 15806 84826 16374
rect 85220 16368 85262 16384
rect 85256 15790 85257 15791
rect 85255 15789 85256 15790
rect 85268 15778 85302 16402
rect 85308 16396 85372 16402
rect 85314 16390 85315 16391
rect 86013 16390 86014 16391
rect 85313 16389 85314 16390
rect 86014 16389 86015 16390
rect 85308 16368 85344 16384
rect 85313 15790 85314 15791
rect 86014 15790 86015 15791
rect 85314 15789 85315 15790
rect 86013 15789 86014 15790
rect 86026 15778 86060 16402
rect 86710 16396 86778 16402
rect 86072 16390 86073 16391
rect 86071 16389 86072 16390
rect 86738 16368 86778 16394
rect 86071 15790 86072 15791
rect 86772 15790 86773 15791
rect 86072 15789 86073 15790
rect 86771 15789 86772 15790
rect 86784 15778 86818 16402
rect 86824 16396 86890 16402
rect 86824 16368 86862 16394
rect 87529 16390 87530 16391
rect 87530 16389 87531 16390
rect 86829 15790 86830 15791
rect 87530 15790 87531 15791
rect 86830 15789 86831 15790
rect 87529 15789 87530 15790
rect 87542 15778 87576 16402
rect 88218 16396 88294 16402
rect 87588 16390 87589 16391
rect 87587 16389 87588 16390
rect 88250 16378 88284 16396
rect 88287 16390 88288 16391
rect 88288 16389 88289 16390
rect 88246 16368 88294 16378
rect 87587 15790 87588 15791
rect 87588 15789 87589 15790
rect 88250 15778 88284 16368
rect 88288 15790 88289 15791
rect 88287 15789 88288 15790
rect 88300 15778 88334 16402
rect 88346 16390 88347 16391
rect 88345 16389 88346 16390
rect 88345 15790 88346 15791
rect 88346 15789 88347 15790
rect 88364 15778 88398 16402
rect 88408 16320 88418 16396
rect 88408 16304 88416 16320
rect 88436 16304 88446 16396
rect 88416 16292 88446 16304
rect 88558 16068 89006 16184
rect 88506 15972 89006 16068
rect 88506 15944 88934 15972
rect 89022 15778 89056 16402
rect 89058 15778 89092 16402
rect 89104 16390 89105 16391
rect 89103 16389 89104 16390
rect 89103 15790 89104 15791
rect 89104 15789 89105 15790
rect 89136 15778 89170 16402
rect 89440 15778 89474 16402
rect 89554 15778 89588 16402
rect 89816 15778 89850 16402
rect 90212 15778 90246 16402
rect 90326 15778 90360 16402
rect 90524 16304 90532 16396
rect 90561 16390 90562 16391
rect 90562 16389 90563 16390
rect 90562 15790 90563 15791
rect 90561 15789 90562 15790
rect 90574 15778 90608 16402
rect 90620 16390 90621 16391
rect 90619 16389 90620 16390
rect 90619 15790 90620 15791
rect 90620 15789 90621 15790
rect 90750 15778 90784 16402
rect 90864 15778 90898 16402
rect 91332 15778 91366 16402
rect 91462 16340 91472 16360
rect 91444 16304 91462 16340
rect 91472 16304 91518 16340
rect 91462 16284 91472 16304
rect 91444 15784 91462 15856
rect 91472 15784 91518 15856
rect 91522 15778 91556 16402
rect 91636 15778 91670 16402
rect 91918 16340 91952 16402
rect 92002 16340 92078 16402
rect 91918 16304 91976 16340
rect 91986 16304 92078 16340
rect 91918 15778 91952 16304
rect 92032 15856 92066 16304
rect 92090 15856 92124 16402
rect 92028 15784 92072 15856
rect 92084 15784 92124 15856
rect 92032 15778 92066 15784
rect 92090 15778 92124 15784
rect 92690 15778 92724 16402
rect 92776 16396 92842 16402
rect 92804 16384 92838 16396
rect 92848 16386 92936 16402
rect 92804 16368 92842 16384
rect 92848 16374 92942 16386
rect 92804 15778 92838 16368
rect 92848 15790 92894 16374
rect 92902 16304 92942 16374
rect 92902 15856 92962 16304
rect 92902 15806 92942 15856
rect 92902 15790 92916 15806
rect 92934 15794 92942 15806
rect 92848 15778 92882 15790
rect 84876 15754 92882 15778
rect 84754 15716 84826 15754
rect 84876 15744 92936 15754
rect 85255 15732 85256 15733
rect 85256 15731 85257 15732
rect 83816 15644 84728 15682
rect 84792 15644 84826 15716
rect 85158 15706 85220 15708
rect 85268 15682 85302 15744
rect 85314 15732 85315 15733
rect 86013 15732 86014 15733
rect 85313 15731 85314 15732
rect 86014 15731 86015 15732
rect 86026 15682 86060 15744
rect 86072 15732 86073 15733
rect 86771 15732 86772 15733
rect 86071 15731 86072 15732
rect 86772 15731 86773 15732
rect 86784 15682 86818 15744
rect 86830 15732 86831 15733
rect 87529 15732 87530 15733
rect 86829 15731 86830 15732
rect 87530 15731 87531 15732
rect 87542 15682 87576 15744
rect 87588 15732 87589 15733
rect 87587 15731 87588 15732
rect 85240 15644 85302 15682
rect 85998 15644 86060 15682
rect 86756 15644 86818 15682
rect 87514 15644 87576 15682
rect 88250 15644 88284 15744
rect 88287 15732 88288 15733
rect 88288 15731 88289 15732
rect 72376 15622 72422 15644
rect 72432 15622 73174 15644
rect 72382 15542 72416 15622
rect 72444 15610 73174 15622
rect 73202 15610 73938 15644
rect 73140 15542 73174 15610
rect 73864 15604 73882 15610
rect 73254 15542 73280 15604
rect 73282 15542 73336 15604
rect 73892 15576 73938 15610
rect 73948 15610 74690 15644
rect 74702 15610 75454 15644
rect 75460 15610 76206 15644
rect 76218 15622 76970 15644
rect 76218 15610 76964 15622
rect 76976 15610 77722 15644
rect 77734 15622 78486 15644
rect 77734 15610 78480 15622
rect 78492 15610 79238 15644
rect 79250 15622 80002 15644
rect 80012 15622 80754 15644
rect 79250 15610 79996 15622
rect 80024 15610 80754 15622
rect 80766 15622 81518 15644
rect 80766 15610 81512 15622
rect 81524 15610 82270 15644
rect 82282 15622 83034 15644
rect 82282 15610 83028 15622
rect 83040 15610 83786 15644
rect 83798 15622 84550 15644
rect 84560 15622 85302 15644
rect 83798 15610 84544 15622
rect 84572 15610 85302 15622
rect 85314 15610 86060 15644
rect 86072 15610 86818 15644
rect 86830 15610 87576 15644
rect 87588 15610 88288 15644
rect 73948 15604 73966 15610
rect 73898 15542 73932 15576
rect 74656 15542 74690 15610
rect 75380 15604 75398 15610
rect 75408 15576 75454 15610
rect 75464 15604 75482 15610
rect 75414 15542 75448 15576
rect 76172 15542 76206 15610
rect 76930 15542 76964 15610
rect 77688 15542 77722 15610
rect 78446 15542 78480 15610
rect 79204 15542 79238 15610
rect 79962 15542 79996 15610
rect 80720 15542 80754 15610
rect 81478 15542 81512 15610
rect 82236 15542 82270 15610
rect 82994 15542 83028 15610
rect 83752 15542 83786 15610
rect 83816 15542 83820 15610
rect 84510 15542 84544 15610
rect 84690 15542 84724 15610
rect 84792 15546 84826 15610
rect 84754 15542 84864 15546
rect 85268 15542 85302 15610
rect 86026 15542 86060 15610
rect 86784 15542 86818 15610
rect 87542 15542 87576 15610
rect 88250 15542 88284 15610
rect 88300 15542 88334 15744
rect 88346 15732 88347 15733
rect 88345 15731 88346 15732
rect 88364 15682 88398 15744
rect 89022 15682 89056 15744
rect 89058 15682 89092 15744
rect 89104 15732 89105 15733
rect 89103 15731 89104 15732
rect 88364 15644 88402 15682
rect 89022 15644 89092 15682
rect 89136 15644 89170 15744
rect 89440 15644 89474 15744
rect 89554 15682 89588 15744
rect 89816 15682 89850 15744
rect 89554 15644 89592 15682
rect 89788 15644 89850 15682
rect 90212 15682 90246 15744
rect 90212 15644 90250 15682
rect 90326 15644 90360 15744
rect 90561 15732 90562 15733
rect 90562 15731 90563 15732
rect 90574 15682 90608 15744
rect 90620 15732 90621 15733
rect 90619 15731 90620 15732
rect 90546 15644 90608 15682
rect 90750 15644 90784 15744
rect 90864 15682 90898 15744
rect 91332 15682 91366 15744
rect 90864 15644 90902 15682
rect 91304 15644 91366 15682
rect 91444 15652 91462 15738
rect 91472 15652 91518 15738
rect 91522 15682 91556 15744
rect 91522 15644 91560 15682
rect 91636 15644 91670 15744
rect 91918 15644 91952 15744
rect 92032 15738 92066 15744
rect 92090 15738 92124 15744
rect 92028 15678 92072 15738
rect 92084 15678 92124 15738
rect 92028 15652 92124 15678
rect 92032 15644 92124 15652
rect 92690 15682 92724 15744
rect 92690 15644 92728 15682
rect 92804 15644 92838 15744
rect 88346 15610 89092 15644
rect 89104 15610 89850 15644
rect 89862 15610 90608 15644
rect 90620 15610 91366 15644
rect 91378 15610 92124 15644
rect 92136 15610 92838 15644
rect 88364 15542 88398 15610
rect 89022 15542 89056 15610
rect 89058 15542 89092 15610
rect 89136 15542 89170 15610
rect 89440 15542 89474 15610
rect 89554 15542 89588 15610
rect 89816 15542 89850 15610
rect 90212 15542 90246 15610
rect 90326 15542 90360 15610
rect 90574 15542 90608 15610
rect 90750 15542 90784 15610
rect 90864 15542 90898 15610
rect 91332 15542 91366 15610
rect 91522 15542 91556 15610
rect 91636 15542 91670 15610
rect 91918 15542 91952 15610
rect 92032 15542 92066 15610
rect 92090 15542 92124 15610
rect 92690 15542 92724 15610
rect 92804 15542 92838 15610
rect 92848 15728 92936 15744
rect 92848 15716 92942 15728
rect 92848 15644 92894 15716
rect 92902 15652 92942 15716
rect 92902 15650 92968 15652
rect 92990 15650 92996 15680
rect 92902 15644 92936 15650
rect 93004 15644 93038 16548
rect 93078 15644 93112 16548
rect 93254 16546 93860 16548
rect 93912 16546 94518 16548
rect 94570 16546 95172 16548
rect 95228 16546 95834 16548
rect 93594 16508 93652 16546
rect 94352 16508 94410 16546
rect 95110 16508 95156 16546
rect 95846 16542 95864 16548
rect 95870 16546 96492 16548
rect 95870 16540 95926 16546
rect 93181 16496 93226 16507
rect 93192 15682 93226 16496
rect 93606 15682 93640 16508
rect 93839 16496 93884 16507
rect 93192 15644 93230 15682
rect 93578 15644 93640 15682
rect 93850 15682 93884 16496
rect 94364 15682 94398 16508
rect 94497 16496 94542 16507
rect 93850 15644 93888 15682
rect 94336 15644 94398 15682
rect 94508 15682 94542 16496
rect 95122 15682 95156 16508
rect 94508 15644 94546 15682
rect 95094 15678 95156 15682
rect 95166 16507 95190 16512
rect 95166 15678 95200 16507
rect 95760 16176 95786 16530
rect 95818 16507 95864 16508
rect 95813 16502 95868 16507
rect 95788 16204 95868 16502
rect 95762 15682 95786 16176
rect 95818 15682 95868 16204
rect 95094 15644 95200 15678
rect 95298 15678 95868 15682
rect 95870 16404 95948 16540
rect 96471 16496 96516 16507
rect 95870 15682 95925 16404
rect 96482 15682 96516 16496
rect 95870 15678 96378 15682
rect 95298 15644 96378 15678
rect 96482 15644 96520 15682
rect 96596 15644 96630 16548
rect 96638 15678 96672 16650
rect 96714 16588 96720 16650
rect 96914 16582 99096 16650
rect 96684 16548 99096 16582
rect 96714 15896 96720 16542
rect 96914 16510 99096 16548
rect 96914 16448 99370 16510
rect 96914 16144 99096 16448
rect 99554 16203 99638 16679
rect 99590 16191 99638 16203
rect 99646 16691 99742 16732
rect 99646 16191 99694 16691
rect 99696 16191 99741 16691
rect 100201 16679 100257 16690
rect 100212 16203 100257 16679
rect 100274 16191 100288 16732
rect 100302 16691 100400 16732
rect 100302 16191 100344 16691
rect 100354 16191 100399 16691
rect 100468 16510 100502 16840
rect 100418 16482 100594 16510
rect 100418 16464 100538 16482
rect 100418 16448 100594 16464
rect 99518 16144 100400 16191
rect 96914 16110 99573 16144
rect 99616 16110 100231 16144
rect 100274 16110 100400 16144
rect 96914 16042 99096 16110
rect 99684 16094 99742 16110
rect 100342 16094 100400 16110
rect 100385 16079 100400 16094
rect 99696 16042 99730 16076
rect 100354 16042 100388 16076
rect 100468 16042 100502 16448
rect 100538 16446 100594 16448
rect 96914 16008 100922 16042
rect 92848 15610 93640 15644
rect 93652 15610 94398 15644
rect 94410 15610 95156 15644
rect 92848 15546 92894 15610
rect 92902 15604 92936 15610
rect 92902 15546 92968 15604
rect 92848 15542 92974 15546
rect 92990 15542 92996 15604
rect 93004 15542 93038 15610
rect 93078 15542 93112 15610
rect 93192 15542 93226 15610
rect 93606 15542 93640 15610
rect 93850 15542 93884 15610
rect 94364 15542 94398 15610
rect 94508 15542 94542 15610
rect 95122 15542 95156 15610
rect 95166 15610 95925 15644
rect 95942 15610 96630 15644
rect 95166 15542 95200 15610
rect 95824 15604 95868 15610
rect 95762 15542 95786 15604
rect 95818 15542 95868 15604
rect 95870 15542 95925 15610
rect 96482 15542 96516 15610
rect 96596 15542 96630 15610
rect 96632 15576 96678 15678
rect 96688 15644 96706 15650
rect 96914 15644 99096 16008
rect 99100 15696 99107 15730
rect 100468 15690 100502 16008
rect 101081 15972 101308 17164
rect 101636 16038 101670 17336
rect 101744 17315 101796 17330
rect 102402 17315 102454 17330
rect 101744 17274 102840 17315
rect 101765 17268 102840 17274
rect 103038 17268 103085 17315
rect 101772 17200 101796 17268
rect 101800 17234 102427 17268
rect 101800 17228 101824 17234
rect 101792 17186 101796 17200
rect 101877 17187 101935 17234
rect 102430 17200 102454 17268
rect 102458 17234 103085 17268
rect 103180 17308 103214 17336
rect 103722 17338 105204 17372
rect 102458 17228 102510 17234
rect 101739 17184 101796 17186
rect 101739 17175 101814 17184
rect 101750 16944 101814 17175
rect 101750 16199 101796 16944
rect 101792 16187 101796 16199
rect 101889 16187 101934 17187
rect 102444 17186 102454 17200
rect 102397 17175 102454 17186
rect 102408 17154 102454 17175
rect 102408 16199 102442 17154
rect 102444 16460 102454 17154
rect 102500 16460 102510 17228
rect 102535 17187 102593 17234
rect 102547 17154 102592 17187
rect 103055 17175 103100 17186
rect 102444 16192 102470 16460
rect 101765 16140 101946 16187
rect 102380 16140 102427 16187
rect 102444 16174 102454 16192
rect 101772 16100 101796 16140
rect 101800 16106 102427 16140
rect 101800 16100 101824 16106
rect 101744 16044 101796 16100
rect 101877 16090 101935 16106
rect 102430 16100 102454 16174
rect 102500 16146 102526 16192
rect 102547 16187 102581 17154
rect 103066 16199 103100 17175
rect 102458 16140 102526 16146
rect 102535 16140 102594 16187
rect 103038 16140 103085 16187
rect 102458 16106 103085 16140
rect 102458 16100 102510 16106
rect 101889 16038 101923 16090
rect 102402 16044 102454 16100
rect 102535 16090 102593 16106
rect 103180 16100 103248 17308
rect 102547 16038 102581 16072
rect 103180 16038 103214 16100
rect 101636 16004 103214 16038
rect 103722 16040 103756 17338
rect 103863 17286 103897 17338
rect 103863 17270 103909 17286
rect 104466 17270 104513 17317
rect 103863 17236 104513 17270
rect 104521 17301 104555 17338
rect 104521 17270 104567 17301
rect 104521 17236 104593 17270
rect 103863 17189 103909 17236
rect 104521 17189 104567 17236
rect 103825 17177 103851 17188
rect 103863 17177 103897 17189
rect 104483 17177 104509 17188
rect 104521 17177 104555 17189
rect 103836 16201 103897 17177
rect 104494 16201 104555 17177
rect 103863 16189 103897 16201
rect 104521 16189 104555 16201
rect 104560 16189 104561 17189
rect 103863 16142 103909 16189
rect 104466 16142 104513 16189
rect 103863 16108 104513 16142
rect 104521 16142 104567 16189
rect 104588 16148 104589 17230
rect 104521 16108 104593 16142
rect 104635 16132 104669 17338
rect 105292 16596 105300 16650
rect 103863 16092 103909 16108
rect 103863 16040 103897 16092
rect 104521 16077 104567 16108
rect 104604 16106 104669 16132
rect 104521 16040 104555 16077
rect 104635 16040 104669 16106
rect 103722 16006 105204 16040
rect 105346 16030 105354 16596
rect 105790 16114 106026 16886
rect 106152 16114 109414 20162
rect 116282 20130 117312 20164
rect 117622 20126 117656 26762
rect 117736 20126 117770 20160
rect 118194 20126 118228 20160
rect 118308 20126 118342 26762
rect 128196 26334 128618 26954
rect 136564 26874 137562 26894
rect 129166 26845 129222 26873
rect 128762 26840 129222 26845
rect 136598 26840 137562 26860
rect 129022 26832 129222 26840
rect 141156 26820 141212 26830
rect 128762 26812 129222 26817
rect 128994 26804 129222 26812
rect 129166 26776 129222 26804
rect 142906 26778 144010 26802
rect 141156 26764 141212 26774
rect 142878 26750 144038 26774
rect 144742 26524 144776 26878
rect 141524 26490 149776 26524
rect 141524 26334 141558 26490
rect 144602 26410 144705 26422
rect 144742 26410 144776 26490
rect 141710 26407 144705 26410
rect 141588 26348 141660 26386
rect 141710 26376 144690 26407
rect 144708 26376 144776 26410
rect 144602 26364 144690 26376
rect 141524 26294 141620 26334
rect 123716 26136 127774 26159
rect 129166 26136 130058 26159
rect 131410 26136 131716 26159
rect 136524 26136 136570 26152
rect 136546 26106 136570 26136
rect 136812 26076 137790 26090
rect 138004 26076 138060 26090
rect 130002 26012 131466 26036
rect 141524 25544 141558 26294
rect 141614 26266 141620 26278
rect 141626 26214 141660 26348
rect 141666 26294 144634 26334
rect 141666 26266 144634 26278
rect 144640 26230 144674 26364
rect 144680 26294 144706 26334
rect 144680 26266 144734 26278
rect 141610 26206 141698 26214
rect 141588 26202 141698 26206
rect 144590 26202 144601 26213
rect 141588 26168 144601 26202
rect 141610 26156 141698 26168
rect 141626 25780 141660 26156
rect 144602 26140 144674 26178
rect 144640 25764 144674 26140
rect 144602 25752 144690 25764
rect 144742 25752 144776 26376
rect 213206 26006 213526 26448
rect 141588 25690 141660 25728
rect 141710 25718 144690 25752
rect 144708 25718 144776 25752
rect 214534 25750 215894 25764
rect 144602 25706 144690 25718
rect 141626 25556 141660 25690
rect 141670 25642 144634 25682
rect 141726 25586 144634 25626
rect 144640 25572 144674 25706
rect 144680 25642 144700 25682
rect 144742 25626 144776 25718
rect 144680 25586 144776 25626
rect 141610 25548 141698 25556
rect 141588 25544 141698 25548
rect 144590 25544 144601 25555
rect 136614 25510 144601 25544
rect 141524 25024 141558 25510
rect 141610 25498 141698 25510
rect 141626 25122 141660 25498
rect 144602 25482 144674 25520
rect 144640 25106 144674 25482
rect 144602 25094 144690 25106
rect 144742 25094 144776 25586
rect 141588 25032 141660 25070
rect 141710 25060 144690 25094
rect 144708 25060 144776 25094
rect 144602 25048 144690 25060
rect 141524 24978 141620 25024
rect 141524 24360 141558 24978
rect 141614 24950 141620 24968
rect 141626 24898 141660 25032
rect 141666 24978 144634 25024
rect 141666 24950 144634 24968
rect 141670 24922 144634 24950
rect 144640 24914 144674 25048
rect 144680 24978 144712 25024
rect 144742 24968 144776 25060
rect 144680 24922 144776 24968
rect 141610 24890 141698 24898
rect 141588 24886 141698 24890
rect 144590 24886 144601 24897
rect 141588 24852 144601 24886
rect 141610 24840 141698 24852
rect 141626 24464 141660 24840
rect 144602 24824 144674 24862
rect 144640 24448 144674 24824
rect 144602 24436 144690 24448
rect 144742 24436 144776 24922
rect 214400 24484 215914 24498
rect 214134 24446 214158 24468
rect 141588 24374 141660 24412
rect 141710 24402 144690 24436
rect 144708 24402 144776 24436
rect 214112 24422 214158 24446
rect 222222 24446 222246 24468
rect 222222 24422 222268 24446
rect 144602 24390 144690 24402
rect 141524 24320 141620 24360
rect 141524 23456 141558 24320
rect 141602 24264 141620 24304
rect 141626 24240 141660 24374
rect 141666 24320 144634 24360
rect 141666 24264 144634 24304
rect 144640 24256 144674 24390
rect 144680 24320 144716 24360
rect 144742 24304 144776 24402
rect 144680 24264 144776 24304
rect 141610 24232 141698 24240
rect 141588 24228 141698 24232
rect 144590 24228 144601 24239
rect 141588 24194 144601 24228
rect 141610 24182 141698 24194
rect 141626 23806 141660 24182
rect 144602 24166 144674 24204
rect 144640 23790 144674 24166
rect 144602 23778 144690 23790
rect 144742 23778 144776 24264
rect 141588 23716 141660 23754
rect 141710 23744 144690 23778
rect 144708 23744 144776 23778
rect 144602 23732 144690 23744
rect 141580 23668 141620 23680
rect 141608 23612 141620 23652
rect 141626 23582 141660 23716
rect 141666 23668 144634 23680
rect 141666 23612 144634 23652
rect 144640 23598 144674 23732
rect 144680 23668 144712 23680
rect 144742 23652 144776 23744
rect 144680 23612 144776 23652
rect 141610 23574 141698 23582
rect 141588 23570 141698 23574
rect 144590 23570 144601 23581
rect 141588 23536 144601 23570
rect 141595 23524 141698 23536
rect 144742 23456 144776 23612
rect 136524 23422 144776 23456
rect 141524 23068 141558 23422
rect 209034 23270 210214 23642
rect 145996 23170 146052 23182
rect 145996 23114 146052 23126
rect 214812 22994 214832 23052
rect 214840 22994 214860 23046
rect 140590 22918 140594 22952
rect 140624 22944 140628 22970
rect 141132 22748 141154 22754
rect 141132 22744 141150 22748
rect 141132 22688 141174 22698
rect 141229 22637 141282 22891
rect 214756 22754 215394 22994
rect 141483 22544 141536 22637
rect 142246 22588 142920 22601
rect 141615 22567 142920 22588
rect 141519 22386 141553 22505
rect 141630 22425 142250 22567
rect 142300 22533 142834 22552
rect 142334 22518 142832 22533
rect 142300 22493 142866 22499
rect 142300 22490 142334 22493
rect 142832 22490 142866 22493
rect 142266 22487 142368 22490
rect 142798 22487 142900 22490
rect 142266 22484 142900 22487
rect 142266 22453 142334 22484
rect 142457 22472 142709 22476
rect 142445 22453 142721 22472
rect 142798 22453 142900 22484
rect 141621 22386 142250 22425
rect 141519 22300 142250 22386
rect 126996 21940 127012 21970
rect 126962 21906 126978 21936
rect 141519 21903 141553 22300
rect 141621 22148 142250 22300
rect 142300 22412 142334 22453
rect 142671 22438 142682 22441
rect 142479 22423 142687 22438
rect 142355 22412 142436 22423
rect 142479 22419 142764 22423
rect 142300 22370 142340 22412
rect 142348 22376 142436 22412
rect 142495 22404 142682 22419
rect 142683 22376 142764 22419
rect 142348 22370 142368 22376
rect 142300 22196 142334 22370
rect 142402 22338 142436 22376
rect 142730 22338 142764 22376
rect 142671 22310 142682 22321
rect 142495 22276 142682 22310
rect 142832 22196 142866 22453
rect 214812 22422 214814 22598
rect 214840 22450 214842 22570
rect 142300 22162 142866 22196
rect 141621 22094 141655 22148
rect 141621 21903 142250 22094
rect 142300 22042 142866 22076
rect 142300 21903 142334 22042
rect 142671 21962 142682 21973
rect 142495 21937 142682 21962
rect 142348 21903 142350 21922
rect 142368 21916 142470 21934
rect 142479 21928 142687 21937
rect 142696 21916 142798 21934
rect 142355 21903 142470 21916
rect 142683 21903 142798 21916
rect 142832 21903 142866 22042
rect 215279 21926 215694 21957
rect 211726 21921 215694 21926
rect 220350 21926 220771 21957
rect 220350 21921 225710 21926
rect 136501 21870 144771 21903
rect 206655 21887 210491 21921
rect 211726 21892 225710 21921
rect 215279 21887 220771 21892
rect 136439 21869 144771 21870
rect 136439 21835 136474 21836
rect 123742 21706 131718 21740
rect 136473 21650 136474 21777
rect 136507 21650 136508 21743
rect 124988 20454 127954 21392
rect 128500 21126 130150 21396
rect 130586 21126 131940 21394
rect 134864 21218 134872 21244
rect 128500 21104 131940 21126
rect 116336 20096 119792 20126
rect 116432 20092 119792 20096
rect 109544 18256 109564 19360
rect 105790 16106 109414 16114
rect 105790 16086 106026 16106
rect 106152 16086 109414 16106
rect 105790 16078 109414 16086
rect 105790 16070 106026 16078
rect 105790 16044 106084 16070
rect 96684 15610 99096 15644
rect 96688 15604 96706 15610
rect 96638 15542 96672 15576
rect 96914 15558 99096 15610
rect 97396 15542 97430 15558
rect 98154 15542 98188 15558
rect 98912 15542 98946 15558
rect 72364 15508 98980 15542
rect 73140 13864 73174 15508
rect 73254 14434 73280 15508
rect 73282 14378 73336 15508
rect 73898 13864 73932 15508
rect 71264 13846 74832 13864
rect 71264 13844 71808 13846
rect 72146 13836 74832 13846
rect 72268 13808 72302 13836
rect 73140 13808 73174 13836
rect 73898 13808 73932 13836
rect 71264 13790 74832 13808
rect 71264 13788 71864 13790
rect 72090 13780 74832 13790
rect 72268 13158 72302 13780
rect 72382 13158 72416 13218
rect 73140 13180 73174 13780
rect 73898 13180 73932 13780
rect 79204 13189 79238 15508
rect 79962 13189 79996 15508
rect 72420 13158 73932 13180
rect 69768 13156 73932 13158
rect 69698 13124 73932 13156
rect 69620 12602 69644 12622
rect 69620 12574 69672 12594
rect 69698 12518 69816 13124
rect 69830 12518 70292 13124
rect 72268 13056 72302 13124
rect 72382 13094 72416 13124
rect 72420 13094 73932 13124
rect 72370 13056 73932 13094
rect 71884 13022 73932 13056
rect 69734 12372 69768 12518
rect 69724 12016 69768 12372
rect 55034 10368 56612 10402
rect 22762 9788 29349 9868
rect 29736 9788 29770 9868
rect 30394 9788 30428 9868
rect 30832 9788 30866 9868
rect 30946 9818 30980 9868
rect 31052 9818 31086 9868
rect 31604 9818 31638 9868
rect 31710 9818 31744 9868
rect 32262 9818 32296 9868
rect 32368 9818 32402 9868
rect 30946 9788 30991 9818
rect 31052 9788 31097 9818
rect 31604 9788 31649 9818
rect 31710 9788 31755 9818
rect 32262 9788 32307 9818
rect 32368 9788 32413 9818
rect 32482 9788 32516 9868
rect 32920 9788 32954 9868
rect 33578 9788 33612 9868
rect 34236 9788 34270 9868
rect 34350 9788 34384 9868
rect 51522 9872 54320 9906
rect 22762 9754 34998 9788
rect 22762 9718 29349 9754
rect 22762 9188 24790 9718
rect 22666 9154 24790 9188
rect 22762 9126 24790 9154
rect 18780 8636 22478 8670
rect 18780 8568 19201 8636
rect 19588 8584 19626 8606
rect 19576 8568 19634 8584
rect 19670 8568 19708 8606
rect 19714 8574 19738 8630
rect 20208 8606 20242 8636
rect 20246 8606 20276 8636
rect 20316 8606 20367 8636
rect 20124 8568 20367 8606
rect 18780 8534 19708 8568
rect 19760 8534 20367 8568
rect 18780 7240 19201 8534
rect 19576 8496 19634 8534
rect 20208 8528 20367 8534
rect 20208 8496 20292 8528
rect 20316 8496 20367 8528
rect 20372 8606 20390 8636
rect 20684 8606 20718 8636
rect 20798 8606 20843 8636
rect 20904 8606 20949 8636
rect 20980 8606 21025 8636
rect 21456 8606 21554 8636
rect 21556 8606 21610 8636
rect 21638 8606 21683 8636
rect 22114 8606 22212 8636
rect 22214 8606 22268 8636
rect 22296 8606 22330 8636
rect 22334 8606 22368 8636
rect 20372 8568 21025 8606
rect 21038 8568 21124 8606
rect 21322 8568 21683 8606
rect 21696 8568 22368 8606
rect 20372 8496 20390 8568
rect 20418 8534 21025 8568
rect 21076 8534 21683 8568
rect 21734 8534 22368 8568
rect 19588 7240 19622 8496
rect 19687 8484 19732 8495
rect 19698 7240 19732 8484
rect 20208 7268 20242 8496
rect 20246 7268 20291 8496
rect 20322 8495 20367 8496
rect 20322 8456 20401 8495
rect 20322 8168 20410 8456
rect 20306 8158 20410 8168
rect 20306 7514 20401 8158
rect 20208 7240 20291 7268
rect 18780 7214 20291 7240
rect 18780 7212 19201 7214
rect 19588 7212 19622 7214
rect 19698 7212 19732 7214
rect 20208 7212 20242 7214
rect 20246 7212 20291 7214
rect 18780 7158 20291 7212
rect 18780 6723 19201 7158
rect 15313 6689 19201 6723
rect 15613 6621 15647 6689
rect 15771 6676 15816 6683
rect 15821 6673 15879 6689
rect 16474 6683 16537 6689
rect 16429 6674 16537 6683
rect 16474 6673 16537 6674
rect 15827 6648 15844 6673
rect 16474 6627 16485 6673
rect 16514 6621 16525 6673
rect 16548 6621 16559 6689
rect 16562 6674 17554 6689
rect 17730 6682 18722 6689
rect 17778 6676 17806 6682
rect 17834 6676 17862 6682
rect 18486 6676 18514 6682
rect 17137 6673 17195 6674
rect 17180 6658 17195 6673
rect 17263 6621 17297 6674
rect 18655 6673 18689 6682
rect 18064 6651 18398 6668
rect 18655 6662 18666 6673
rect 18678 6662 18689 6673
rect 18780 6621 19201 6689
rect 15137 6587 19201 6621
rect 14032 6398 14422 6432
rect 13840 5864 13914 6352
rect 14032 5900 14066 6398
rect 14161 6330 14293 6377
rect 14208 6296 14293 6330
rect 14135 6237 14191 6248
rect 14263 6237 14319 6248
rect 14146 6061 14191 6237
rect 14274 6061 14319 6237
rect 14161 6002 14293 6049
rect 14208 5968 14293 6002
rect 14388 5900 14422 6398
rect 14032 5866 14422 5900
rect 14508 6398 14898 6432
rect 14508 5900 14551 6398
rect 14637 6330 14769 6377
rect 14684 6296 14769 6330
rect 14611 6237 14667 6248
rect 14739 6237 14795 6248
rect 14622 6061 14667 6237
rect 14750 6061 14795 6237
rect 14578 5900 14580 6048
rect 14637 6002 14769 6049
rect 14684 5968 14769 6002
rect 14864 5900 14898 6398
rect 14508 5866 14898 5900
rect 13648 5854 13684 5860
rect 13648 5826 13684 5832
rect 13786 5788 13914 5864
rect 14517 5816 14551 5866
rect 13840 5698 13914 5788
rect 13648 5454 13664 5460
rect 13648 5426 13664 5432
rect 14014 5196 14436 5816
rect 14490 5196 14912 5816
rect 14517 4982 14551 5196
rect 16514 5166 16525 6587
rect 16548 5166 16559 6587
rect 17149 4982 17183 6587
rect 17263 4883 17297 6587
rect 18780 6551 19201 6587
rect 18926 5156 18960 6551
rect 19040 5308 19074 6551
rect 19588 5296 19622 7158
rect 19698 5308 19732 7158
rect 20208 6644 20242 7158
rect 20246 7098 20291 7158
rect 20322 7098 20401 7514
rect 20246 7080 20280 7098
rect 20246 6728 20286 7080
rect 20322 6796 20390 7098
rect 20356 6780 20390 6796
rect 20350 6746 20390 6780
rect 20684 6746 20718 8534
rect 20798 7098 20843 8534
rect 20904 7098 20949 8534
rect 20980 8495 21025 8534
rect 20980 7098 21059 8495
rect 21456 7098 21501 8534
rect 21562 7098 21607 8534
rect 21638 8495 21683 8534
rect 21638 7098 21717 8495
rect 22114 7098 22159 8534
rect 22220 7098 22265 8534
rect 22296 8500 22330 8534
rect 22334 8518 22368 8534
rect 22334 8500 22398 8518
rect 20798 6796 20832 7098
rect 20904 6784 20938 7098
rect 20980 6796 21048 7098
rect 21456 6796 21490 7098
rect 21562 6812 21596 7098
rect 21638 6812 21706 7098
rect 21014 6784 21048 6796
rect 21562 6784 21606 6812
rect 21632 6796 21706 6812
rect 22114 6796 22148 7098
rect 21632 6784 21666 6796
rect 21672 6784 21706 6796
rect 22220 6784 22254 7098
rect 22296 6796 22398 8500
rect 22330 6784 22398 6796
rect 20892 6746 20950 6784
rect 21014 6746 21052 6784
rect 21550 6752 21608 6784
rect 21550 6746 21666 6752
rect 21672 6746 21710 6784
rect 22208 6746 22266 6784
rect 22318 6746 22398 6784
rect 22444 6746 22478 8636
rect 22762 7952 24273 9126
rect 24665 7952 24710 9126
rect 24886 8796 24931 9718
rect 24958 9478 28582 9718
rect 24958 9468 28610 9478
rect 24886 8142 24920 8796
rect 24886 8044 24931 8142
rect 24800 7962 24931 8044
rect 24886 7952 24931 7962
rect 24958 7952 28582 9468
rect 22762 7918 24570 7952
rect 22762 7777 24273 7918
rect 24309 7850 24441 7897
rect 24356 7816 24441 7850
rect 22762 7765 24272 7777
rect 24283 7765 24339 7768
rect 24411 7765 24467 7768
rect 24536 7765 24570 7918
rect 24656 7918 28582 7952
rect 24656 7890 24710 7918
rect 24886 7897 24920 7918
rect 24656 7765 24724 7890
rect 24782 7782 24800 7884
rect 24870 7850 24920 7897
rect 24816 7816 24920 7850
rect 24886 7795 24920 7816
rect 24886 7777 24932 7795
rect 24920 7773 24932 7777
rect 24759 7765 24804 7768
rect 24887 7765 24932 7768
rect 22762 7718 24817 7765
rect 24858 7718 24932 7765
rect 24958 7718 28582 7918
rect 22762 7616 24272 7718
rect 24290 7695 24943 7718
rect 24283 7684 24943 7695
rect 24948 7684 28582 7718
rect 24294 7616 24339 7684
rect 24422 7616 24467 7684
rect 24536 7616 24570 7684
rect 24653 7668 24724 7684
rect 24656 7616 24690 7668
rect 24699 7616 24724 7668
rect 24770 7616 24804 7684
rect 24898 7616 24932 7684
rect 24958 7616 28582 7684
rect 22762 7582 28582 7616
rect 22762 7546 24272 7582
rect 24294 7581 24339 7582
rect 24422 7581 24467 7582
rect 22772 7098 22817 7546
rect 22772 6796 22806 7098
rect 22848 6752 22876 7546
rect 22904 6752 22932 7546
rect 22936 7478 23010 7546
rect 22954 7098 22999 7478
rect 23430 7098 23475 7546
rect 22954 6796 22988 7098
rect 23430 6796 23464 7098
rect 23500 6872 23528 7546
rect 23556 6752 23584 7546
rect 23612 7098 23657 7546
rect 23612 6796 23646 7098
rect 23726 6746 23760 7546
rect 23857 7420 24272 7546
rect 24309 7522 24441 7569
rect 24356 7488 24441 7522
rect 24536 7420 24570 7582
rect 23857 7386 24570 7420
rect 24656 7420 24690 7582
rect 24699 7482 24724 7582
rect 24770 7581 24815 7582
rect 24898 7581 24943 7582
rect 24785 7522 24917 7569
rect 24958 7530 28582 7582
rect 24832 7488 24917 7522
rect 25012 7420 25046 7530
rect 24656 7386 25046 7420
rect 25132 7420 25166 7530
rect 25261 7522 25380 7530
rect 25266 7512 25380 7522
rect 25444 7513 25470 7530
rect 25282 7488 25380 7512
rect 25282 7448 25372 7488
rect 25266 7434 25282 7436
rect 25488 7420 25522 7530
rect 25132 7386 25522 7420
rect 23857 7336 24272 7386
rect 23857 6746 24584 7336
rect 20356 6744 24584 6746
rect 20246 6648 20280 6728
rect 20350 6723 24584 6744
rect 24638 6723 25060 7336
rect 25114 6723 25536 7336
rect 20350 6712 24637 6723
rect 24638 6716 25536 6723
rect 25761 6723 25795 7530
rect 25875 7098 25920 7530
rect 25947 7414 25950 7530
rect 25975 7522 26026 7530
rect 25975 7414 25978 7522
rect 25947 7106 25950 7214
rect 25875 6782 25909 7098
rect 25975 7078 25978 7214
rect 25981 7098 26026 7522
rect 26533 7098 26578 7530
rect 26639 7498 26684 7530
rect 26598 7224 26950 7498
rect 26639 7098 26684 7224
rect 27191 7098 27236 7530
rect 27291 7098 27342 7530
rect 25981 6782 26015 7098
rect 26533 7016 26573 7098
rect 26533 6782 26567 7016
rect 26639 6782 26673 7098
rect 27191 6782 27225 7098
rect 27291 7038 27331 7098
rect 27297 6782 27331 7038
rect 27411 6723 27445 7530
rect 20246 6644 20291 6648
rect 20294 6644 20312 6688
rect 20350 6648 20390 6712
rect 20350 6644 20401 6648
rect 20684 6644 20718 6712
rect 20892 6696 20950 6712
rect 20904 6648 20938 6696
rect 21014 6648 21048 6712
rect 21550 6708 21608 6712
rect 21672 6708 21706 6712
rect 21550 6706 21706 6708
rect 21550 6696 21608 6706
rect 21562 6648 21596 6696
rect 21606 6650 21634 6652
rect 20904 6644 20949 6648
rect 21014 6644 21059 6648
rect 21562 6644 21607 6648
rect 21610 6644 21634 6650
rect 21666 6648 21706 6706
rect 22208 6696 22266 6712
rect 22318 6696 22398 6712
rect 22220 6648 22254 6696
rect 21666 6644 21717 6648
rect 22220 6644 22265 6648
rect 22324 6644 22326 6696
rect 22334 6678 22398 6696
rect 22330 6644 22398 6678
rect 22444 6644 22478 6712
rect 22848 6694 22876 6706
rect 22904 6700 22932 6706
rect 23556 6694 23584 6706
rect 23726 6696 23760 6712
rect 23726 6685 23737 6696
rect 23749 6685 23760 6696
rect 23857 6689 24637 6712
rect 24727 6689 25295 6716
rect 25761 6689 27445 6723
rect 23857 6644 24272 6689
rect 25761 6673 25795 6689
rect 25761 6662 25772 6673
rect 25784 6662 25795 6673
rect 27411 6673 27445 6689
rect 27411 6662 27422 6673
rect 27434 6662 27445 6673
rect 20208 6621 24272 6644
rect 28928 6644 29349 9718
rect 30492 8230 30506 8430
rect 30520 8202 30534 8458
rect 30832 6746 30866 9754
rect 30946 8796 30991 9754
rect 31052 8796 31097 9754
rect 31604 8796 31649 9754
rect 31710 8796 31755 9754
rect 32262 8796 32307 9754
rect 32368 8796 32413 9754
rect 30946 6796 30980 8796
rect 31052 6796 31086 8796
rect 31604 8508 31638 8796
rect 31604 6994 31644 8508
rect 31604 6796 31638 6994
rect 31710 6796 31744 8796
rect 32262 7138 32296 8796
rect 32368 8544 32402 8796
rect 32362 7138 32402 8544
rect 32262 6796 32307 7138
rect 32368 6796 32413 7138
rect 32482 7012 32516 9754
rect 34350 9622 34384 9754
rect 41648 9660 42568 9694
rect 32920 7988 32954 9622
rect 33560 7988 33634 8132
rect 32900 7350 33362 7988
rect 33376 7350 33838 7988
rect 32920 7300 32954 7350
rect 33578 7300 33612 7334
rect 32920 7266 33304 7300
rect 32920 7012 32988 7266
rect 33074 7198 33184 7236
rect 33112 7164 33184 7198
rect 33057 7114 33113 7125
rect 33145 7114 33201 7125
rect 33068 7012 33113 7114
rect 33156 7012 33201 7114
rect 33270 7012 33304 7266
rect 33430 7266 33780 7300
rect 33430 7012 33464 7266
rect 33574 7232 33660 7236
rect 33554 7198 33660 7232
rect 33572 7194 33660 7198
rect 33572 7164 33664 7194
rect 33572 7148 33624 7164
rect 33650 7160 33664 7164
rect 33533 7114 33566 7125
rect 33578 7114 33620 7148
rect 33650 7132 33692 7138
rect 33544 7012 33620 7114
rect 33624 7125 33662 7126
rect 33624 7012 33677 7125
rect 33746 7012 33780 7266
rect 34236 7012 34270 9622
rect 41648 9468 41682 9660
rect 42392 9592 42430 9630
rect 41824 9558 42430 9592
rect 41751 9508 41796 9519
rect 42409 9508 42454 9519
rect 41762 9468 41796 9508
rect 41807 9480 41808 9481
rect 42408 9480 42409 9481
rect 41808 9479 41809 9480
rect 42407 9479 42408 9480
rect 42420 9468 42454 9508
rect 42534 9468 42568 9660
rect 41020 9428 41276 9450
rect 41614 9434 42568 9468
rect 41048 9400 41248 9422
rect 41048 8822 41248 8844
rect 41020 8794 41276 8816
rect 41648 8810 41682 9434
rect 41762 8810 41796 9434
rect 41808 9422 41809 9423
rect 42407 9422 42408 9423
rect 41807 9421 41808 9422
rect 42408 9421 42409 9422
rect 41814 9352 41816 9364
rect 41814 9324 41844 9336
rect 41956 9100 42404 9216
rect 41904 9004 42404 9100
rect 41904 8976 42332 9004
rect 41807 8822 41808 8823
rect 42408 8822 42409 8823
rect 41808 8821 41809 8822
rect 42407 8821 42408 8822
rect 42420 8810 42454 9434
rect 42534 8810 42568 9434
rect 42678 9272 42706 9770
rect 46422 9714 46436 9768
rect 42838 9660 43758 9694
rect 42838 9468 42872 9660
rect 43582 9592 43620 9630
rect 43014 9558 43620 9592
rect 42941 9508 42986 9519
rect 43599 9508 43644 9519
rect 42952 9468 42986 9508
rect 42997 9480 42998 9481
rect 43598 9480 43599 9481
rect 42998 9479 42999 9480
rect 43597 9479 43598 9480
rect 43610 9468 43644 9508
rect 43724 9468 43758 9660
rect 44148 9668 45068 9702
rect 44148 9468 44182 9668
rect 44892 9600 44930 9638
rect 44324 9566 44930 9600
rect 44228 9552 44330 9556
rect 44886 9552 44988 9556
rect 44256 9527 44302 9528
rect 44914 9527 44960 9528
rect 44251 9524 44302 9527
rect 44909 9524 44960 9527
rect 44251 9516 44296 9524
rect 44909 9516 44954 9524
rect 44262 9468 44296 9516
rect 44307 9480 44308 9481
rect 44908 9480 44909 9481
rect 44308 9479 44309 9480
rect 44907 9479 44908 9480
rect 44920 9468 44954 9516
rect 45034 9468 45068 9668
rect 45316 9676 46236 9710
rect 45316 9468 45350 9676
rect 46060 9608 46098 9646
rect 45492 9574 46098 9608
rect 45396 9558 45498 9564
rect 45356 9552 45516 9558
rect 46054 9552 46156 9564
rect 45424 9535 45470 9536
rect 46082 9535 46128 9536
rect 45419 9530 45470 9535
rect 45384 9524 45488 9530
rect 46077 9524 46128 9535
rect 45430 9468 45464 9524
rect 45475 9480 45476 9481
rect 46076 9480 46077 9481
rect 45476 9479 45477 9480
rect 46075 9479 46076 9480
rect 46088 9468 46122 9524
rect 46202 9468 46236 9676
rect 42804 9434 43758 9468
rect 44114 9434 45068 9468
rect 45282 9434 46236 9468
rect 46250 9434 46270 9468
rect 42650 9142 42678 9160
rect 42678 9104 42706 9142
rect 42650 9086 42678 9104
rect 42838 8810 42872 9434
rect 42952 8810 42986 9434
rect 42998 9422 42999 9423
rect 43597 9422 43598 9423
rect 42997 9421 42998 9422
rect 43598 9421 43599 9422
rect 42997 8822 42998 8823
rect 43598 8822 43599 8823
rect 42998 8821 42999 8822
rect 43597 8821 43598 8822
rect 43610 8810 43644 9434
rect 43724 8810 43758 9434
rect 44148 8810 44182 9434
rect 44262 8810 44296 9434
rect 44308 9422 44309 9423
rect 44907 9422 44908 9423
rect 44307 9421 44308 9422
rect 44908 9421 44909 9422
rect 44307 8822 44308 8823
rect 44908 8822 44909 8823
rect 44308 8821 44309 8822
rect 44907 8821 44908 8822
rect 44920 8810 44954 9434
rect 45034 8810 45068 9434
rect 45316 8810 45350 9434
rect 45430 8810 45464 9434
rect 45476 9422 45477 9423
rect 46075 9422 46076 9423
rect 45475 9421 45476 9422
rect 46076 9421 46077 9422
rect 45475 8822 45476 8823
rect 46076 8822 46077 8823
rect 45476 8821 45477 8822
rect 46075 8821 46076 8822
rect 46088 8810 46122 9434
rect 46202 8810 46236 9434
rect 41614 8776 42568 8810
rect 42804 8776 43758 8810
rect 44114 8776 45068 8810
rect 45282 8776 46236 8810
rect 46250 8776 46270 8810
rect 41648 8380 41682 8776
rect 41762 8532 41796 8776
rect 41808 8764 41809 8765
rect 42407 8764 42408 8765
rect 41807 8763 41808 8764
rect 42408 8763 42409 8764
rect 42420 8532 42454 8776
rect 42392 8482 42430 8520
rect 41824 8448 42430 8482
rect 42534 8380 42568 8776
rect 41648 8346 42568 8380
rect 42838 8380 42872 8776
rect 42952 8532 42986 8776
rect 42998 8764 42999 8765
rect 43597 8764 43598 8765
rect 42997 8763 42998 8764
rect 43598 8763 43599 8764
rect 43610 8532 43644 8776
rect 43582 8482 43620 8520
rect 43014 8448 43620 8482
rect 43724 8380 43758 8776
rect 42838 8346 43758 8380
rect 41020 8236 41276 8250
rect 43010 8236 43560 8238
rect 41048 8208 41248 8222
rect 43038 8208 43532 8210
rect 44148 8152 44182 8776
rect 44262 8152 44296 8776
rect 44308 8764 44309 8765
rect 44907 8764 44908 8765
rect 44307 8763 44308 8764
rect 44908 8763 44909 8764
rect 44920 8176 44954 8776
rect 45034 8176 45068 8776
rect 44307 8164 44308 8165
rect 44308 8163 44309 8164
rect 44822 8152 45280 8176
rect 45316 8152 45350 8776
rect 45430 8152 45464 8776
rect 45476 8764 45477 8765
rect 46075 8764 46076 8765
rect 45475 8763 45476 8764
rect 46076 8763 46077 8764
rect 45475 8164 45476 8165
rect 46076 8164 46077 8165
rect 45476 8163 45477 8164
rect 46075 8163 46076 8164
rect 46088 8152 46122 8776
rect 46202 8152 46236 8776
rect 41048 8118 45280 8152
rect 45282 8118 46236 8152
rect 46250 8118 46270 8152
rect 44148 8038 44182 8118
rect 44262 8038 44296 8118
rect 44822 8084 45280 8118
rect 44900 8038 44986 8084
rect 45034 8038 45068 8084
rect 45316 8038 45350 8118
rect 45430 8038 45464 8118
rect 46088 8038 46122 8118
rect 46202 8038 46236 8118
rect 41048 8004 46340 8038
rect 46476 8004 46490 9714
rect 47280 8010 47288 9540
rect 34928 7454 34968 7458
rect 35032 7454 35082 7458
rect 34928 7434 35082 7454
rect 34928 7430 34968 7434
rect 35032 7430 35082 7434
rect 35244 7436 35484 7988
rect 44148 7850 44182 8004
rect 44900 7936 44986 8004
rect 45034 7850 45068 8004
rect 45316 7858 45350 8004
rect 46202 7858 46236 8004
rect 35508 7436 35558 7446
rect 35244 7434 35558 7436
rect 34932 7406 35086 7426
rect 35244 7408 35484 7434
rect 35508 7430 35558 7434
rect 35244 7406 35562 7408
rect 35244 7350 35484 7406
rect 38884 7398 38904 7456
rect 38912 7398 38932 7450
rect 34420 7152 34620 7194
rect 38828 7158 39466 7398
rect 34392 7124 34648 7138
rect 32418 6746 34534 7012
rect 38884 6826 38886 7002
rect 38912 6854 38914 6974
rect 30456 6720 34534 6746
rect 30456 6712 34580 6720
rect 30832 6696 30866 6712
rect 30832 6685 30843 6696
rect 30855 6685 30866 6696
rect 32418 6644 34580 6712
rect 28928 6634 34580 6644
rect 28928 6621 34534 6634
rect 20208 6610 34534 6621
rect 20246 5736 20291 6610
rect 20350 6242 20401 6610
rect 20246 5296 20280 5736
rect 20284 5548 20314 5736
rect 20356 5548 20401 6242
rect 20904 6120 20949 6610
rect 21014 6120 21059 6610
rect 20904 5800 21354 6120
rect 21388 5800 21392 6120
rect 20904 5548 20949 5800
rect 21014 5548 21059 5800
rect 21562 5548 21607 6610
rect 21610 6242 21634 6610
rect 21666 6242 21717 6610
rect 21672 5548 21717 6242
rect 22220 5548 22265 6610
rect 22324 6242 22326 6610
rect 20356 5308 20390 5548
rect 20904 5296 20938 5548
rect 21014 5308 21048 5548
rect 21562 5296 21596 5548
rect 21672 5308 21706 5548
rect 22220 5296 22254 5548
rect 22334 5342 22398 6610
rect 22330 5308 22398 5342
rect 19576 5258 19634 5296
rect 19670 5258 19708 5296
rect 20234 5258 20292 5296
rect 20328 5258 20366 5296
rect 20892 5258 20950 5296
rect 20986 5258 21024 5296
rect 21550 5258 21608 5296
rect 21644 5258 21682 5296
rect 22208 5258 22266 5296
rect 19102 5224 19708 5258
rect 19760 5224 20366 5258
rect 20418 5224 21024 5258
rect 21076 5224 21682 5258
rect 21734 5224 22266 5258
rect 22300 5224 22318 5258
rect 19576 5208 19634 5224
rect 20234 5208 20292 5224
rect 20892 5208 20950 5224
rect 21550 5208 21608 5224
rect 22208 5208 22266 5224
rect 22251 5193 22266 5208
rect 22334 5156 22368 5308
rect 22444 5218 22478 6610
rect 23857 6587 29349 6610
rect 23857 6574 24272 6587
rect 28928 6574 29349 6587
rect 32418 6316 34534 6610
rect 47280 6606 47288 7226
rect 47906 7048 47940 9528
rect 48564 7048 48598 9528
rect 49186 9236 49212 9534
rect 49222 7048 49256 9528
rect 49880 7048 49914 9528
rect 51522 9074 51556 9872
rect 51778 9820 51825 9851
rect 51766 9804 51825 9820
rect 52266 9804 52313 9851
rect 52436 9820 52483 9851
rect 52424 9804 52483 9820
rect 52924 9804 52971 9851
rect 53094 9820 53141 9851
rect 53082 9804 53141 9820
rect 53582 9804 53629 9851
rect 53752 9820 53798 9851
rect 53740 9804 53798 9820
rect 51698 9770 52313 9804
rect 52356 9770 52971 9804
rect 53014 9770 53629 9804
rect 53672 9770 53798 9804
rect 51668 9722 51708 9764
rect 51625 9711 51708 9722
rect 51636 9235 51708 9711
rect 51668 9182 51708 9235
rect 51724 9182 51736 9764
rect 51766 9723 51824 9770
rect 51778 9223 51812 9723
rect 52283 9711 52328 9722
rect 52294 9235 52328 9711
rect 51766 9176 51825 9223
rect 52266 9176 52313 9223
rect 52330 9182 52364 9764
rect 52386 9182 52420 9764
rect 52424 9723 52482 9770
rect 53082 9764 53140 9770
rect 53740 9764 53798 9770
rect 52436 9223 52470 9723
rect 52941 9711 52986 9722
rect 52472 9480 52768 9542
rect 52952 9235 52986 9711
rect 52424 9176 52483 9223
rect 52924 9176 52971 9223
rect 52988 9182 53036 9764
rect 53044 9723 53140 9764
rect 53044 9223 53092 9723
rect 53094 9223 53128 9723
rect 53599 9711 53644 9722
rect 53610 9235 53644 9711
rect 53044 9182 53141 9223
rect 53082 9176 53141 9182
rect 53582 9176 53629 9223
rect 53672 9182 53686 9764
rect 53700 9723 53798 9764
rect 53700 9223 53742 9723
rect 53752 9223 53786 9723
rect 53866 9542 53900 9872
rect 53816 9514 53992 9542
rect 53816 9496 53936 9514
rect 53816 9480 53992 9496
rect 53700 9182 53798 9223
rect 53740 9176 53798 9182
rect 51698 9142 52313 9176
rect 52356 9142 52971 9176
rect 53014 9142 53629 9176
rect 53672 9142 53798 9176
rect 51766 9126 51824 9142
rect 52424 9126 52482 9142
rect 53082 9126 53140 9142
rect 53740 9126 53798 9142
rect 53783 9111 53798 9126
rect 51778 9074 51812 9108
rect 52436 9074 52470 9108
rect 53094 9074 53128 9108
rect 53752 9074 53786 9108
rect 53866 9074 53900 9480
rect 53936 9478 53992 9480
rect 51522 9040 54320 9074
rect 53866 8722 53900 9040
rect 54479 9004 54706 10196
rect 55034 9070 55068 10368
rect 55142 10347 55194 10362
rect 55800 10347 55852 10362
rect 55142 10306 56238 10347
rect 55163 10300 56238 10306
rect 56436 10300 56483 10347
rect 55170 10232 55194 10300
rect 55198 10266 55825 10300
rect 55198 10260 55222 10266
rect 55190 10218 55194 10232
rect 55275 10219 55333 10266
rect 55828 10232 55852 10300
rect 55856 10266 56483 10300
rect 56578 10340 56612 10368
rect 57120 10370 58602 10404
rect 55856 10260 55908 10266
rect 55137 10216 55194 10218
rect 55137 10207 55212 10216
rect 55148 10186 55212 10207
rect 55148 9231 55182 10186
rect 55190 9976 55212 10186
rect 55287 10186 55332 10219
rect 55842 10218 55852 10232
rect 55795 10207 55852 10218
rect 55806 10186 55852 10207
rect 55190 9206 55194 9976
rect 55287 9219 55321 10186
rect 55806 9231 55840 10186
rect 55842 9492 55852 10186
rect 55898 9492 55908 10260
rect 55933 10219 55991 10266
rect 55945 10186 55990 10219
rect 56453 10207 56498 10218
rect 55842 9224 55868 9492
rect 55170 9132 55194 9206
rect 55198 9172 55222 9178
rect 55275 9172 55334 9219
rect 55778 9172 55825 9219
rect 55842 9206 55852 9224
rect 55198 9138 55825 9172
rect 55198 9132 55222 9138
rect 55142 9076 55194 9132
rect 55275 9122 55333 9138
rect 55828 9132 55852 9206
rect 55898 9178 55924 9224
rect 55945 9219 55979 10186
rect 56464 9231 56498 10207
rect 55856 9172 55924 9178
rect 55933 9172 55992 9219
rect 56436 9172 56483 9219
rect 55856 9138 56483 9172
rect 55856 9132 55908 9138
rect 55287 9070 55321 9104
rect 55800 9076 55852 9132
rect 55933 9122 55991 9138
rect 56578 9132 56646 10340
rect 55945 9070 55979 9104
rect 56578 9070 56612 9132
rect 55034 9036 56612 9070
rect 57120 9072 57154 10370
rect 57261 10318 57295 10370
rect 57261 10302 57307 10318
rect 57864 10302 57911 10349
rect 57261 10268 57911 10302
rect 57919 10333 57953 10370
rect 57919 10302 57965 10333
rect 57919 10268 57991 10302
rect 57261 10221 57307 10268
rect 57919 10221 57965 10268
rect 57223 10209 57249 10220
rect 57261 10209 57295 10221
rect 57881 10209 57907 10220
rect 57919 10209 57953 10221
rect 57234 9233 57295 10209
rect 57892 9233 57953 10209
rect 57261 9221 57295 9233
rect 57919 9221 57953 9233
rect 57958 9221 57959 10221
rect 57261 9174 57307 9221
rect 57864 9174 57911 9221
rect 57261 9140 57911 9174
rect 57919 9174 57965 9221
rect 57986 9180 57987 10262
rect 57919 9140 57991 9174
rect 58033 9164 58067 10370
rect 58690 9628 58698 9682
rect 57261 9124 57307 9140
rect 57261 9072 57295 9124
rect 57919 9109 57965 9140
rect 58002 9138 58067 9164
rect 57919 9072 57953 9109
rect 58033 9072 58067 9138
rect 57120 9038 58602 9072
rect 58744 9062 58752 9628
rect 59188 9146 59424 9918
rect 59550 9146 62812 11719
rect 62942 11410 62962 11719
rect 66093 11288 66127 11742
rect 66093 10968 66564 11288
rect 65460 10682 65469 10904
rect 65494 10716 65503 10904
rect 66093 9622 66127 10968
rect 69734 9622 69768 12016
rect 69850 11960 69882 12502
rect 69884 12434 70234 12468
rect 69884 11954 69918 12434
rect 70076 12366 70114 12404
rect 70042 12332 70114 12366
rect 69987 12282 70032 12293
rect 70075 12282 70120 12293
rect 69998 12106 70032 12282
rect 70086 12106 70120 12282
rect 70076 12056 70114 12094
rect 70042 12022 70114 12056
rect 70200 11954 70234 12434
rect 69884 11920 70234 11954
rect 71898 11414 71918 12390
rect 72268 11798 72302 13022
rect 72370 12984 73932 13022
rect 72382 12860 73932 12984
rect 72344 12852 73932 12860
rect 72344 12712 73976 12852
rect 72382 12704 73976 12712
rect 72382 11950 73932 12704
rect 72420 11938 73902 11950
rect 72406 11900 73902 11938
rect 72420 11798 73902 11900
rect 76643 11798 80267 13189
rect 80720 11950 80754 15508
rect 84510 15112 84544 15508
rect 84690 15112 84724 15508
rect 84792 15148 84864 15508
rect 85268 15133 85313 15508
rect 86026 15133 86071 15508
rect 86784 15133 86829 15508
rect 87542 15133 87587 15508
rect 88250 15348 88284 15508
rect 88300 15348 88345 15508
rect 88364 15500 88409 15508
rect 89022 15500 89103 15508
rect 88388 15450 89032 15488
rect 88426 15416 89032 15450
rect 89058 15348 89103 15500
rect 89136 15348 89170 15508
rect 88250 15314 89170 15348
rect 89440 15348 89474 15508
rect 89554 15500 89599 15508
rect 89816 15488 89861 15508
rect 90212 15500 90257 15508
rect 89578 15450 90222 15488
rect 89616 15416 90222 15450
rect 89816 15348 89861 15416
rect 90326 15348 90360 15508
rect 89440 15314 90360 15348
rect 88300 15133 88345 15314
rect 89058 15133 89103 15314
rect 89706 15204 89764 15206
rect 89706 15148 89764 15178
rect 89816 15133 89861 15314
rect 89888 15204 89972 15206
rect 89888 15148 89972 15178
rect 90574 15133 90619 15508
rect 85256 15132 85257 15133
rect 85268 15132 85314 15133
rect 86014 15132 86015 15133
rect 86026 15132 86072 15133
rect 86772 15132 86773 15133
rect 86784 15132 86830 15133
rect 87530 15132 87531 15133
rect 87542 15132 87588 15133
rect 88288 15132 88289 15133
rect 88300 15132 88346 15133
rect 89046 15132 89047 15133
rect 89058 15132 89104 15133
rect 89804 15132 89805 15133
rect 89816 15132 89862 15133
rect 90562 15132 90563 15133
rect 90574 15132 90620 15133
rect 85255 15131 85256 15132
rect 84865 15120 85256 15131
rect 85268 15120 85302 15132
rect 85314 15131 85315 15132
rect 86013 15131 86014 15132
rect 85314 15120 86014 15131
rect 86026 15120 86060 15132
rect 86072 15131 86073 15132
rect 86771 15131 86772 15132
rect 86072 15120 86772 15131
rect 86784 15120 86818 15132
rect 86830 15131 86831 15132
rect 87529 15131 87530 15132
rect 86830 15120 87530 15131
rect 87542 15120 87576 15132
rect 87588 15131 87589 15132
rect 88287 15131 88288 15132
rect 87588 15120 88288 15131
rect 88300 15120 88334 15132
rect 88346 15131 88347 15132
rect 89045 15131 89046 15132
rect 88346 15120 89046 15131
rect 89058 15120 89092 15132
rect 89104 15131 89105 15132
rect 89803 15131 89804 15132
rect 89104 15120 89804 15131
rect 89816 15120 89850 15132
rect 89862 15131 89863 15132
rect 90561 15131 90562 15132
rect 89862 15120 90562 15131
rect 90574 15120 90608 15132
rect 90620 15131 90621 15132
rect 90750 15131 90784 15508
rect 90864 15131 90909 15508
rect 91332 15131 91377 15508
rect 91444 15168 91462 15204
rect 91472 15168 91518 15204
rect 91462 15148 91472 15168
rect 91522 15144 91567 15508
rect 91636 15144 91670 15508
rect 91424 15131 91882 15144
rect 91918 15131 91952 15508
rect 92032 15204 92077 15508
rect 92090 15204 92135 15508
rect 92028 15168 92077 15204
rect 92084 15168 92135 15204
rect 92032 15148 92084 15168
rect 92032 15131 92077 15148
rect 92090 15131 92135 15168
rect 92690 15164 92735 15508
rect 92690 15148 92778 15164
rect 92690 15131 92735 15148
rect 92776 15131 92778 15148
rect 92804 15131 92838 15508
rect 90620 15120 92838 15131
rect 92848 15132 92894 15508
rect 92902 15148 92974 15508
rect 92990 15176 92996 15508
rect 92934 15136 92942 15148
rect 92848 15120 92882 15132
rect 84876 15112 92882 15120
rect 84398 15086 92882 15112
rect 84398 15006 85112 15086
rect 85268 15006 85302 15086
rect 86026 15006 86060 15086
rect 86784 15006 86818 15086
rect 87542 15006 87576 15086
rect 88300 15006 88334 15086
rect 89058 15006 89092 15086
rect 89816 15006 89850 15086
rect 90574 15006 90608 15086
rect 90750 15006 90784 15086
rect 90864 15006 90909 15086
rect 91332 15006 91377 15086
rect 91424 15052 91882 15086
rect 91502 15032 91588 15052
rect 91444 15006 91462 15032
rect 91472 15006 91588 15032
rect 91636 15006 91670 15052
rect 91918 15006 91952 15086
rect 92032 15032 92077 15086
rect 92090 15032 92135 15086
rect 92028 15006 92077 15032
rect 92084 15006 92135 15032
rect 92690 15006 92735 15086
rect 92776 15006 92778 15080
rect 92804 15006 92838 15086
rect 92848 15006 92882 15086
rect 93004 15006 93038 15508
rect 84398 14972 93038 15006
rect 84398 14554 85112 14972
rect 86026 14884 86060 14972
rect 86026 14798 86124 14884
rect 85362 14698 85364 14700
rect 86026 14588 86060 14798
rect 84510 13158 84544 14554
rect 84832 14500 85380 14534
rect 84832 14218 84866 14500
rect 85202 14434 85234 14454
rect 85007 14426 85205 14431
rect 85007 14420 85206 14426
rect 85018 14414 85206 14420
rect 84896 14376 85006 14414
rect 85018 14410 85306 14414
rect 85018 14386 85312 14410
rect 85202 14380 85312 14386
rect 85206 14376 85312 14380
rect 84934 14342 85006 14376
rect 85007 14332 85205 14343
rect 85244 14342 85312 14376
rect 85018 14298 85205 14332
rect 85256 14326 85294 14342
rect 85346 14218 85380 14500
rect 84832 14184 85380 14218
rect 85430 14408 86068 14588
rect 85430 14322 86124 14408
rect 85430 14126 86068 14322
rect 85470 14112 85792 14126
rect 86026 14112 86060 14126
rect 84832 14024 85380 14058
rect 84832 13742 84866 14024
rect 85184 13978 85202 13986
rect 84968 13966 85244 13978
rect 85180 13955 85202 13966
rect 85180 13950 85205 13955
rect 85180 13944 85206 13950
rect 85002 13938 85210 13944
rect 84896 13900 84968 13938
rect 85002 13934 85306 13938
rect 85002 13932 85312 13934
rect 85018 13922 85312 13932
rect 85018 13910 85205 13922
rect 85206 13900 85312 13922
rect 84934 13866 84968 13900
rect 85194 13856 85205 13867
rect 85244 13866 85312 13900
rect 85018 13822 85205 13856
rect 85256 13850 85294 13866
rect 85346 13742 85380 14024
rect 84832 13708 85380 13742
rect 85430 13650 86068 14112
rect 81750 13124 85302 13158
rect 81416 11882 81462 11906
rect 81442 11860 81462 11882
rect 81750 11798 81784 13124
rect 83128 13094 83152 13124
rect 82236 13072 82274 13094
rect 82224 13056 82282 13072
rect 82494 13056 82532 13094
rect 82994 13072 83032 13094
rect 82982 13056 83040 13072
rect 83072 13062 83096 13094
rect 83128 13062 83190 13094
rect 83752 13072 83790 13094
rect 83152 13056 83190 13062
rect 83740 13056 83798 13072
rect 83810 13056 83848 13094
rect 84468 13056 84506 13094
rect 81926 13022 82532 13056
rect 82584 13022 83190 13056
rect 83242 13022 83848 13056
rect 83900 13022 84506 13056
rect 84510 13072 84544 13124
rect 82224 12984 82282 13022
rect 82982 12984 83040 13022
rect 81853 12972 81898 12983
rect 81864 11938 81898 12972
rect 82236 11950 82270 12984
rect 82511 12972 82556 12983
rect 82522 11938 82556 12972
rect 82994 11950 83028 12984
rect 81852 11900 81910 11938
rect 82208 11900 82246 11938
rect 82510 11900 82568 11938
rect 82966 11900 83004 11938
rect 83072 11906 83096 13016
rect 83128 11906 83152 13016
rect 83740 12984 83798 13022
rect 83169 12972 83214 12983
rect 83180 11938 83214 12972
rect 83752 12418 83786 12984
rect 83832 12983 83848 12984
rect 83862 12983 83878 12984
rect 83827 12972 83878 12983
rect 83752 11950 83792 12418
rect 83832 12390 83878 12972
rect 83890 12390 83906 13012
rect 84510 12984 84556 13072
rect 85126 13056 85164 13094
rect 84558 13022 85164 13056
rect 84485 12972 84498 12983
rect 84510 12972 84544 12984
rect 85143 12972 85188 12983
rect 83770 11938 83792 11950
rect 83798 11938 83872 12390
rect 84496 11950 84544 12972
rect 84496 11938 84530 11950
rect 85154 11938 85188 12972
rect 85268 12420 85302 13124
rect 86026 12856 86060 13650
rect 83168 11900 83226 11938
rect 83724 11900 83762 11938
rect 81852 11866 82246 11900
rect 82298 11866 83004 11900
rect 83056 11866 83762 11900
rect 83798 11900 83884 11938
rect 84482 11900 84530 11938
rect 83798 11882 84530 11900
rect 81852 11850 81910 11866
rect 82510 11850 82568 11866
rect 83168 11850 83226 11866
rect 83798 11860 83810 11882
rect 83814 11866 84530 11882
rect 83826 11850 83884 11866
rect 84484 11850 84530 11866
rect 81852 11835 81867 11850
rect 81864 11798 81898 11832
rect 82522 11798 82556 11832
rect 83180 11798 83214 11832
rect 83838 11798 83872 11832
rect 84496 11798 84530 11850
rect 84532 11832 84536 11934
rect 84560 11900 84564 11906
rect 85142 11900 85200 11938
rect 85234 11910 85242 12392
rect 85262 11938 85302 12420
rect 89816 11950 89850 14972
rect 90750 14756 90784 14972
rect 90864 14908 90909 14972
rect 91332 14896 91377 14972
rect 91444 14896 91462 14972
rect 91472 14904 91588 14972
rect 91472 14896 91518 14904
rect 90888 14858 91532 14896
rect 90926 14824 91532 14858
rect 91320 14808 91378 14824
rect 91332 14756 91366 14808
rect 91636 14756 91670 14972
rect 90750 14722 91670 14756
rect 91918 14764 91952 14972
rect 92028 14916 92077 14972
rect 92028 14904 92072 14916
rect 92084 14904 92135 14972
rect 92690 14916 92735 14972
rect 92776 14966 92778 14972
rect 92078 14900 92700 14904
rect 92060 14866 92700 14900
rect 92078 14832 92700 14866
rect 92078 14816 92136 14832
rect 92804 14764 92838 14972
rect 92848 14826 92872 14972
rect 91918 14730 92838 14764
rect 91332 11950 91366 14722
rect 92216 14534 92550 14680
rect 92216 14502 92638 14534
rect 93078 13168 93112 15508
rect 93192 13966 93237 15508
rect 93606 13966 93651 15508
rect 93850 13966 93895 15508
rect 93192 13320 93226 13966
rect 93606 13308 93640 13966
rect 93850 13320 93884 13966
rect 94364 13308 94409 15508
rect 94508 14016 94553 15508
rect 95122 14978 95156 15508
rect 95088 14194 95100 14978
rect 95116 14194 95156 14978
rect 94584 14024 94906 14028
rect 95122 14016 95156 14194
rect 95166 14016 95211 15508
rect 95762 14958 95786 15508
rect 95818 14978 95868 15508
rect 95824 14016 95868 14978
rect 95870 15014 95925 15508
rect 95870 14194 95948 15014
rect 95870 14016 95925 14194
rect 96482 14016 96527 15508
rect 96596 14016 96630 15508
rect 96638 14016 96672 15508
rect 96864 14024 97114 14028
rect 94508 13320 97102 14016
rect 98364 13980 98686 14488
rect 98424 13806 98576 13980
rect 94510 13308 97102 13320
rect 93594 13270 93652 13308
rect 93822 13270 93860 13308
rect 94114 13270 97102 13308
rect 93254 13236 93860 13270
rect 93912 13236 97102 13270
rect 93594 13220 93652 13236
rect 94352 13220 94410 13236
rect 94510 13168 97102 13236
rect 93078 13134 97102 13168
rect 99059 13153 99060 13207
rect 94510 13122 97102 13134
rect 95050 12770 95064 12974
rect 95078 12742 95092 12974
rect 95122 11950 95156 13122
rect 95880 11950 95914 13122
rect 96638 11950 96672 13122
rect 84556 11866 84564 11900
rect 84572 11866 85200 11900
rect 85234 11866 85256 11900
rect 84560 11860 84564 11866
rect 85142 11850 85200 11866
rect 85185 11835 85200 11850
rect 85154 11798 85188 11832
rect 85268 11798 85302 11938
rect 85314 11866 85349 11900
rect 72268 11764 80267 11798
rect 81368 11764 98964 11798
rect 72420 11604 73902 11764
rect 76643 11728 80267 11764
rect 72480 9622 72514 11604
rect 73138 9622 73172 11604
rect 73252 9622 73286 11604
rect 81750 9622 81784 11764
rect 83914 11286 83934 11482
rect 84496 9622 84530 11764
rect 85268 9622 85302 11764
rect 99077 11728 99096 13189
rect 101117 13180 101151 15972
rect 101231 13180 101265 15972
rect 99820 13153 101302 13180
rect 101889 13153 101923 16004
rect 99113 11764 99114 13153
rect 99209 13119 102665 13153
rect 99820 13098 101302 13119
rect 101889 13113 101923 13119
rect 101883 13098 101923 13113
rect 99820 13051 101946 13098
rect 102489 13057 102536 13098
rect 102478 13051 102536 13057
rect 99289 13017 101878 13051
rect 101889 13017 102536 13051
rect 99193 12622 99216 12822
rect 99221 12594 99244 12850
rect 99193 12222 99216 12422
rect 99221 12194 99244 12450
rect 99193 11822 99216 12022
rect 99221 11794 99244 12050
rect 99820 11938 101302 13017
rect 101889 12970 101935 13017
rect 102478 13011 102501 13017
rect 102506 12983 102529 13017
rect 101848 12958 101877 12969
rect 101889 12958 101934 12970
rect 102506 12958 102535 12969
rect 102547 12958 102581 13119
rect 101859 11950 101934 12958
rect 101859 11938 101893 11950
rect 99820 11857 101906 11938
rect 102446 11897 102454 12668
rect 102474 11897 102482 12640
rect 102517 11950 102581 12958
rect 102517 11938 102551 11950
rect 102505 11891 102563 11938
rect 101951 11857 102563 11891
rect 102593 11857 102610 11891
rect 99820 11789 101302 11857
rect 101847 11841 101893 11857
rect 102446 11828 102454 11851
rect 101859 11789 101893 11823
rect 102474 11800 102482 11851
rect 102505 11841 102551 11857
rect 102517 11789 102551 11823
rect 102631 11789 102665 13119
rect 103770 12184 103786 13698
rect 104635 13194 104669 16006
rect 105790 15994 106026 16044
rect 105332 15970 105336 15980
rect 106152 15968 109414 16078
rect 105506 15800 105582 15802
rect 105478 15772 105610 15774
rect 105488 15550 105598 15570
rect 105526 15512 105560 15532
rect 106188 14414 106222 15968
rect 107716 14434 107730 15622
rect 105352 14392 106444 14414
rect 105352 14388 106404 14392
rect 104148 13158 104705 13194
rect 106188 13158 106222 14388
rect 107744 14378 107786 15678
rect 111265 13410 111299 20025
rect 114018 16404 114045 19942
rect 114052 16438 114079 19976
rect 114702 18890 114853 19144
rect 114956 18432 115107 18890
rect 114740 18398 115218 18432
rect 114740 17944 114760 18398
rect 114956 18376 115107 18398
rect 114796 18342 115218 18376
rect 114796 17888 114816 18342
rect 114956 16568 115107 18342
rect 116300 16682 117394 18890
rect 115187 16648 117394 16682
rect 115440 16636 115938 16648
rect 115590 16568 115788 16596
rect 116300 16568 117394 16648
rect 114956 16534 117394 16568
rect 114956 16498 115107 16534
rect 116300 16498 117394 16534
rect 117622 16544 117656 20092
rect 117736 20055 117774 20062
rect 117724 19990 117774 20055
rect 118194 20055 118232 20062
rect 118194 20040 118240 20055
rect 118182 20024 118240 20040
rect 117828 19990 118240 20024
rect 117724 19952 117770 19990
rect 118182 19952 118240 19990
rect 117736 19940 117770 19952
rect 117782 19940 117800 19951
rect 117736 18478 117800 19940
rect 117730 17360 117800 18478
rect 117714 17292 117800 17360
rect 117714 17086 117811 17292
rect 118194 17240 118228 19952
rect 118308 17240 118342 20092
rect 119656 20042 119738 20058
rect 119656 20014 119724 20030
rect 119716 18948 119808 18970
rect 118920 18010 119924 18948
rect 123281 18916 123315 20025
rect 123520 19690 126869 20157
rect 128500 20126 130150 21104
rect 130586 20126 131940 21104
rect 134780 20966 134798 21188
rect 134808 21165 134872 21188
rect 134814 21162 134872 21165
rect 136098 21165 136170 21186
rect 136098 21162 136164 21165
rect 136098 20990 136120 21162
rect 128352 20092 131940 20126
rect 128352 19766 128386 20092
rect 128500 20024 130150 20092
rect 130412 20024 130450 20062
rect 130586 20024 131940 20092
rect 128500 19990 130450 20024
rect 130502 19990 131940 20024
rect 128500 19958 130150 19990
rect 130586 19956 131940 19990
rect 131729 19952 131730 19953
rect 131802 19952 131824 19956
rect 131730 19951 131731 19952
rect 128455 19940 128500 19951
rect 129113 19940 129158 19951
rect 129771 19940 129816 19951
rect 130429 19940 130474 19951
rect 131087 19940 131132 19951
rect 128466 19766 128500 19940
rect 128511 19778 128512 19779
rect 129112 19778 129113 19779
rect 128512 19777 128513 19778
rect 129111 19777 129112 19778
rect 129124 19766 129158 19940
rect 129169 19778 129170 19779
rect 129770 19778 129771 19779
rect 129170 19777 129171 19778
rect 129769 19777 129770 19778
rect 129782 19766 129816 19940
rect 129827 19778 129828 19779
rect 130428 19778 130429 19779
rect 129828 19777 129829 19778
rect 130427 19777 130428 19778
rect 130440 19766 130474 19940
rect 130485 19778 130486 19779
rect 131086 19778 131087 19779
rect 130486 19777 130487 19778
rect 131085 19777 131086 19778
rect 131098 19766 131132 19940
rect 131744 19794 131824 19952
rect 131143 19778 131144 19779
rect 131744 19778 131802 19794
rect 131144 19777 131145 19778
rect 131718 19772 131729 19777
rect 131718 19766 131730 19772
rect 128318 19738 131734 19766
rect 131750 19742 131768 19778
rect 131787 19763 131802 19778
rect 131750 19738 131802 19742
rect 128318 19732 131802 19738
rect 128352 19690 128386 19732
rect 128466 19690 128500 19732
rect 128512 19720 128513 19721
rect 129111 19720 129112 19721
rect 128511 19719 128512 19720
rect 129112 19719 129113 19720
rect 123520 19119 128852 19690
rect 129124 19392 129158 19732
rect 129170 19720 129171 19721
rect 129769 19720 129770 19721
rect 129169 19719 129170 19720
rect 129770 19719 129771 19720
rect 129782 19392 129816 19732
rect 129828 19720 129829 19721
rect 130427 19720 130428 19721
rect 129827 19719 129828 19720
rect 130428 19719 130429 19720
rect 129046 19186 129080 19192
rect 129080 19136 129102 19186
rect 129124 19121 129169 19392
rect 129216 19186 129298 19192
rect 129112 19120 129113 19121
rect 129124 19120 129170 19121
rect 129111 19119 129112 19120
rect 123520 19118 129112 19119
rect 129124 19118 129158 19120
rect 129170 19119 129171 19120
rect 129222 19119 129242 19136
rect 129250 19119 129298 19186
rect 129782 19121 129827 19392
rect 129770 19120 129771 19121
rect 129782 19120 129828 19121
rect 130428 19120 130429 19121
rect 129769 19119 129770 19120
rect 129170 19118 129770 19119
rect 123520 19108 129770 19118
rect 129782 19108 129816 19120
rect 129828 19119 129829 19120
rect 130427 19119 130428 19120
rect 129828 19108 130406 19119
rect 130440 19108 130474 19732
rect 130486 19720 130487 19721
rect 131085 19720 131086 19721
rect 130485 19719 130486 19720
rect 131086 19719 131087 19720
rect 130485 19120 130486 19121
rect 131086 19120 131087 19121
rect 130486 19119 130487 19120
rect 131085 19119 131086 19120
rect 131098 19108 131132 19732
rect 131722 19726 131730 19732
rect 131144 19720 131145 19721
rect 131143 19719 131144 19720
rect 131734 19704 131802 19732
rect 131744 19136 131824 19704
rect 131143 19120 131144 19121
rect 131744 19120 131802 19136
rect 131144 19119 131145 19120
rect 131718 19108 131729 19119
rect 123520 19080 131734 19108
rect 131756 19084 131768 19120
rect 131787 19105 131802 19120
rect 131752 19080 131802 19084
rect 123520 19074 131802 19080
rect 123520 18952 128852 19074
rect 129054 19068 129222 19074
rect 129054 18982 129242 19068
rect 129250 18982 129298 19068
rect 129769 19062 129770 19063
rect 129782 19062 129816 19074
rect 129828 19062 129829 19063
rect 130427 19062 130428 19063
rect 129770 19061 129771 19062
rect 129782 19061 129828 19062
rect 130428 19061 130429 19062
rect 129054 18952 129222 18982
rect 129782 18952 129827 19061
rect 123395 18916 123429 18950
rect 123520 18916 130246 18952
rect 122564 18882 130246 18916
rect 123281 18814 123315 18882
rect 123520 18861 130246 18882
rect 123184 18432 123194 18756
rect 123281 18755 123282 18787
rect 123286 18755 123315 18814
rect 123234 18728 123280 18733
rect 123281 18728 123315 18755
rect 123383 18780 130246 18861
rect 123383 18733 123441 18780
rect 123212 18721 123315 18728
rect 123212 18718 123274 18721
rect 123212 18460 123250 18718
rect 123234 18288 123250 18460
rect 123276 18460 123315 18721
rect 123234 17745 123274 18288
rect 123276 17745 123280 18460
rect 123234 17733 123280 17745
rect 123247 17729 123274 17733
rect 123281 17695 123315 18460
rect 123395 18288 123440 18733
rect 123520 18450 130246 18780
rect 130356 18534 130400 18554
rect 130400 18498 130412 18534
rect 130428 18462 130429 18463
rect 130427 18461 130428 18462
rect 130440 18450 130474 19074
rect 130486 19062 130487 19063
rect 131085 19062 131086 19063
rect 130485 19061 130486 19062
rect 131086 19061 131087 19062
rect 130485 18462 130486 18463
rect 131086 18462 131087 18463
rect 130486 18461 130487 18462
rect 131085 18461 131086 18462
rect 131098 18450 131132 19074
rect 131144 19062 131145 19063
rect 131143 19061 131144 19062
rect 131734 19046 131802 19074
rect 131744 18478 131824 19046
rect 131143 18462 131144 18463
rect 131744 18462 131802 18478
rect 131144 18461 131145 18462
rect 131718 18450 131729 18461
rect 123520 18416 131734 18450
rect 123520 18336 130246 18416
rect 130400 18336 130412 18362
rect 130440 18336 130474 18416
rect 131098 18336 131132 18416
rect 131756 18382 131768 18462
rect 131787 18447 131802 18462
rect 123520 18302 131802 18336
rect 123395 17733 123429 18288
rect 123520 18266 130246 18302
rect 123898 18228 123943 18266
rect 123898 17900 123932 18228
rect 124012 18098 124046 18266
rect 124053 18098 124093 18266
rect 124098 18252 124166 18266
rect 124098 18098 124149 18252
rect 124554 18098 124588 18266
rect 124668 18098 124702 18266
rect 124711 18098 124745 18266
rect 124866 18248 125088 18266
rect 125264 18230 125280 18266
rect 125326 18098 125360 18266
rect 125369 18098 125409 18266
rect 125420 18098 125437 18266
rect 125978 18230 126018 18266
rect 125984 18098 126018 18230
rect 126027 18098 126056 18266
rect 126098 18098 126132 18266
rect 126658 18106 126726 18266
rect 126760 18106 126785 18266
rect 126799 18106 126833 18266
rect 128316 18114 130246 18266
rect 130400 18254 130412 18302
rect 123990 17900 124982 18098
rect 123662 17733 124982 17900
rect 123286 17686 123315 17695
rect 123383 17686 123442 17733
rect 123520 17731 124982 17733
rect 123520 17686 125088 17731
rect 123286 17684 125088 17686
rect 125180 17684 126172 18098
rect 123286 17652 126172 17684
rect 123281 17584 123315 17652
rect 123383 17636 123441 17652
rect 123662 17650 126172 17652
rect 123383 17621 123398 17636
rect 123395 17584 123429 17618
rect 123662 17584 124996 17650
rect 122564 17582 124996 17584
rect 125018 17582 125056 17642
rect 125110 17594 125134 17640
rect 125124 17582 125134 17594
rect 125180 17582 126172 17650
rect 122564 17550 126172 17582
rect 117736 17068 117811 17086
rect 117710 16840 117856 17068
rect 117676 16800 117682 16830
rect 117704 16828 117710 16830
rect 117736 16726 117811 16840
rect 117838 16828 117862 16830
rect 117866 16800 117890 16830
rect 117702 16656 117708 16698
rect 117730 16696 117811 16726
rect 117730 16684 117736 16696
rect 117766 16684 117811 16696
rect 117898 16684 119924 17240
rect 121910 17083 121926 17114
rect 121880 17068 121926 17083
rect 120002 17006 120014 17018
rect 119998 16818 120014 17006
rect 120002 16810 120014 16818
rect 117762 16646 119924 16684
rect 117766 16612 119924 16646
rect 117766 16596 117812 16612
rect 117898 16544 119924 16612
rect 117622 16510 119924 16544
rect 116336 14414 116370 16498
rect 117898 15802 119924 16510
rect 121844 15986 121880 16780
rect 121900 15986 121908 16724
rect 118008 15652 118220 15802
rect 118424 15618 118458 15652
rect 119320 15634 119532 15802
rect 119740 15618 119774 15652
rect 119854 15618 119888 15802
rect 123281 15674 123315 17550
rect 123662 17548 126172 17550
rect 123662 17478 124996 17548
rect 123990 17424 124996 17478
rect 123662 17070 124996 17424
rect 125018 17130 125056 17548
rect 125124 17536 125134 17548
rect 123662 17002 124982 17070
rect 123990 16678 124982 17002
rect 125180 16678 126172 17548
rect 123399 15674 123429 16661
rect 126490 16627 127482 18106
rect 127658 18082 130246 18114
rect 130440 18082 130474 18116
rect 131098 18082 131132 18116
rect 131756 18082 131790 18116
rect 131870 18082 131904 19956
rect 134816 18198 134854 20966
rect 134872 18254 134882 20966
rect 136369 18315 136568 21650
rect 141519 19083 141553 21869
rect 141621 21857 142250 21869
rect 141630 21827 142250 21857
rect 142300 21829 142334 21869
rect 142348 21835 142350 21869
rect 142402 21846 142436 21869
rect 142730 21863 142764 21869
rect 142722 21854 142774 21863
rect 142724 21850 142770 21854
rect 142730 21846 142764 21850
rect 142484 21841 142682 21845
rect 142495 21829 142671 21834
rect 142694 21829 142802 21835
rect 142832 21829 142866 21869
rect 144737 21841 144771 21869
rect 142266 21827 142900 21829
rect 141630 21823 144614 21827
rect 141630 21801 144626 21823
rect 141574 21795 144626 21801
rect 144703 21795 144805 21841
rect 207035 21835 207046 21846
rect 207058 21835 207069 21846
rect 207035 21819 207069 21835
rect 208530 21825 208558 21838
rect 209200 21825 209228 21838
rect 209256 21825 209284 21838
rect 209908 21825 209936 21838
rect 210077 21819 210111 21857
rect 141574 21789 142250 21795
rect 142300 21789 142334 21795
rect 142832 21789 142866 21795
rect 141574 21774 144592 21789
rect 141574 21761 144669 21774
rect 141574 21755 144587 21761
rect 141605 21743 142250 21755
rect 141621 21672 142250 21743
rect 142300 21749 142356 21755
rect 142300 21720 142334 21749
rect 142832 21720 142866 21755
rect 144588 21727 144669 21761
rect 142300 21686 142866 21720
rect 141621 21199 141655 21672
rect 141998 21224 142128 21240
rect 142328 21224 143456 21240
rect 142026 21196 142128 21212
rect 142328 21196 143428 21212
rect 142850 21177 143428 21196
rect 144635 21183 144669 21727
rect 142850 21171 144314 21177
rect 144588 21171 144685 21183
rect 144737 21171 144771 21795
rect 207035 21785 210111 21819
rect 141714 21165 149690 21171
rect 141574 21143 141655 21144
rect 141574 21131 141689 21143
rect 141698 21137 149690 21165
rect 141574 21125 141655 21131
rect 141664 21125 144592 21131
rect 141574 21116 144592 21125
rect 141574 21103 144669 21116
rect 141574 21097 144587 21103
rect 141605 21085 141702 21097
rect 141621 20541 141655 21085
rect 142128 21068 142328 21078
rect 144588 21069 144669 21103
rect 142100 21040 142356 21050
rect 144635 20525 144669 21069
rect 144588 20513 144685 20525
rect 144737 20513 144771 21137
rect 141714 20507 144685 20513
rect 141574 20485 141655 20486
rect 141698 20485 144685 20507
rect 141574 20473 141689 20485
rect 141698 20479 144626 20485
rect 144703 20479 144805 20513
rect 141574 20467 141655 20473
rect 141664 20467 144592 20473
rect 141574 20458 144592 20467
rect 141574 20445 144669 20458
rect 141574 20439 144587 20445
rect 141605 20427 141702 20439
rect 141621 19883 141655 20427
rect 144588 20411 144669 20445
rect 142936 20390 144288 20408
rect 142908 20362 144316 20380
rect 141976 19902 143434 19920
rect 142004 19874 143406 19892
rect 144635 19867 144669 20411
rect 144588 19855 144685 19867
rect 144737 19855 144771 20479
rect 141714 19849 144685 19855
rect 141574 19827 141655 19828
rect 141698 19827 144685 19849
rect 141574 19815 141689 19827
rect 141698 19821 144626 19827
rect 144703 19821 144805 19855
rect 141574 19809 141655 19815
rect 141664 19809 144592 19815
rect 141574 19800 144592 19809
rect 141574 19787 144669 19800
rect 141574 19781 144587 19787
rect 141605 19769 141702 19781
rect 141621 19225 141655 19769
rect 144588 19753 144669 19787
rect 144635 19209 144669 19753
rect 144588 19197 144685 19209
rect 144737 19197 144771 19821
rect 141714 19191 144685 19197
rect 141698 19169 144685 19191
rect 141698 19163 144626 19169
rect 144703 19163 144805 19197
rect 149715 19175 149722 19248
rect 149749 19209 149756 19282
rect 141664 19129 144592 19157
rect 141676 19125 144576 19129
rect 144635 19083 144669 19111
rect 144737 19083 144771 19163
rect 141519 19049 149789 19083
rect 144737 18447 144771 19049
rect 192758 18820 192792 19552
rect 193530 18914 193564 18948
rect 194188 18914 194222 18948
rect 195360 18916 195370 18970
rect 195476 18916 195484 18950
rect 196108 18916 196142 18950
rect 196766 18916 196800 18950
rect 197424 18916 197458 18950
rect 197538 18916 197572 19558
rect 193310 18880 194888 18914
rect 192758 18378 192802 18820
rect 144152 18354 144410 18366
rect 192768 18098 192802 18378
rect 193310 18316 193344 18880
rect 193446 18744 193470 18846
rect 193530 18828 193577 18859
rect 193474 18812 193498 18818
rect 193518 18812 193577 18828
rect 194054 18812 194101 18859
rect 193474 18778 194101 18812
rect 193474 18772 193498 18778
rect 193518 18731 193576 18778
rect 194104 18744 194122 18846
rect 194188 18828 194235 18859
rect 194132 18812 194150 18818
rect 194176 18812 194235 18828
rect 194712 18812 194759 18859
rect 194854 18852 194888 18880
rect 194820 18818 194888 18852
rect 195414 18860 195424 18916
rect 195438 18882 198870 18916
rect 195438 18860 195448 18882
rect 194132 18778 194759 18812
rect 194132 18776 194150 18778
rect 194176 18776 194234 18778
rect 194132 18772 194234 18776
rect 194176 18748 194234 18772
rect 194152 18744 194234 18748
rect 193413 18719 193458 18730
rect 193424 18465 193458 18719
rect 193530 18477 193564 18731
rect 194071 18719 194116 18730
rect 194082 18465 194116 18719
rect 194124 18550 194146 18726
rect 194152 18522 194174 18744
rect 194176 18731 194234 18744
rect 194188 18477 194222 18731
rect 194729 18719 194774 18730
rect 194740 18465 194774 18719
rect 194854 18511 194914 18818
rect 194846 18477 194914 18511
rect 193412 18418 193471 18465
rect 193502 18424 193549 18465
rect 193494 18418 193549 18424
rect 194070 18418 194129 18465
rect 194160 18424 194207 18465
rect 194148 18418 194207 18424
rect 194728 18418 194786 18465
rect 193412 18384 193549 18418
rect 193592 18384 194207 18418
rect 194250 18384 194786 18418
rect 194820 18384 194834 18418
rect 193412 18368 193470 18384
rect 193494 18378 193514 18384
rect 193412 18353 193427 18368
rect 193522 18350 193542 18384
rect 194070 18368 194128 18384
rect 194148 18378 194172 18384
rect 194176 18350 194200 18384
rect 194728 18368 194786 18384
rect 194771 18353 194786 18368
rect 194854 18316 194888 18477
rect 195414 18322 195448 18860
rect 195450 18467 195482 18860
rect 196108 18830 196155 18861
rect 196096 18814 196155 18830
rect 196158 18814 196205 18861
rect 196766 18830 196813 18861
rect 196754 18814 196813 18830
rect 196816 18814 196863 18861
rect 197424 18830 197470 18861
rect 197412 18814 197470 18830
rect 197538 18814 197572 18882
rect 195590 18780 196205 18814
rect 196248 18780 196863 18814
rect 196906 18780 197470 18814
rect 197474 18780 197492 18814
rect 195494 18732 195518 18761
rect 196096 18733 196154 18780
rect 196754 18774 196828 18780
rect 196754 18754 196812 18774
rect 196754 18746 196838 18754
rect 196754 18733 196812 18746
rect 197412 18744 197470 18780
rect 197538 18755 197544 18787
rect 197548 18755 197572 18814
rect 197412 18733 197492 18744
rect 195522 18732 195546 18733
rect 195494 18721 195562 18732
rect 195494 18478 195518 18721
rect 195522 18471 195562 18721
rect 196108 18514 196148 18733
rect 196175 18728 196220 18732
rect 196158 18721 196220 18728
rect 196158 18542 196176 18721
rect 196108 18483 196142 18514
rect 196186 18471 196220 18721
rect 196766 18483 196800 18733
rect 196833 18721 196878 18732
rect 196844 18471 196878 18721
rect 197424 18494 197464 18733
rect 197468 18522 197492 18733
rect 197424 18483 197458 18494
rect 195516 18424 195575 18471
rect 196080 18424 196127 18471
rect 196174 18424 196233 18471
rect 196738 18424 196785 18471
rect 196832 18424 196891 18471
rect 197396 18424 197443 18471
rect 195516 18390 196127 18424
rect 196170 18390 196785 18424
rect 196828 18390 197443 18424
rect 195516 18374 195574 18390
rect 196174 18374 196232 18390
rect 196832 18374 196890 18390
rect 195516 18359 195531 18374
rect 197502 18322 197510 18356
rect 197538 18322 197572 18755
rect 192854 18282 194898 18316
rect 195414 18288 197572 18322
rect 193310 18178 193344 18282
rect 193204 18158 193866 18178
rect 193246 18138 193812 18158
rect 193310 18134 193344 18138
rect 193274 18110 193812 18134
rect 193310 18098 193344 18110
rect 194854 18098 194888 18282
rect 195414 18106 195448 18288
rect 127658 18048 132310 18082
rect 127658 17980 130246 18048
rect 130256 17980 130294 18018
rect 130440 17996 130478 18018
rect 130428 17980 130486 17996
rect 130914 17980 130952 18018
rect 131098 17996 131136 18018
rect 131086 17980 131144 17996
rect 131572 17980 131610 18018
rect 131756 18011 131794 18018
rect 131756 17996 131802 18011
rect 131744 17980 131802 17996
rect 127658 17946 130294 17980
rect 130346 17946 130952 17980
rect 131004 17946 131610 17980
rect 131662 17946 131802 17980
rect 127658 16663 130246 17946
rect 130273 17896 130318 17907
rect 130284 16663 130318 17896
rect 130322 16663 130356 17940
rect 130378 16663 130412 17940
rect 130428 17908 130486 17946
rect 130440 16663 130474 17908
rect 130931 17896 130976 17907
rect 130942 16663 130976 17896
rect 130980 16663 131020 17940
rect 131036 16663 131076 17940
rect 131086 17908 131144 17946
rect 131098 16663 131132 17908
rect 131589 17896 131634 17907
rect 131600 16663 131634 17896
rect 131700 16663 131728 17940
rect 131744 17908 131802 17946
rect 131756 16663 131790 17908
rect 127658 16627 131835 16663
rect 123433 16593 131835 16627
rect 123433 15674 123467 16593
rect 123984 16513 124041 16524
rect 124053 16513 124087 16593
rect 124677 16546 124682 16548
rect 124705 16546 124710 16576
rect 124099 16518 124699 16524
rect 124711 16518 124745 16593
rect 125369 16574 125409 16593
rect 125335 16524 125354 16546
rect 124757 16518 124984 16524
rect 124099 16513 124998 16518
rect 125182 16513 125357 16524
rect 125363 16519 125409 16574
rect 125416 16524 125437 16578
rect 125369 16513 125403 16519
rect 125415 16513 126015 16524
rect 126027 16513 126061 16593
rect 126490 16534 127482 16593
rect 127510 16562 131835 16593
rect 127510 16534 127544 16562
rect 126073 16513 126182 16524
rect 126490 16513 127578 16534
rect 127658 16528 131835 16562
rect 127652 16526 131835 16528
rect 127639 16513 131835 16526
rect 123488 16451 123569 16498
rect 123628 16479 131835 16513
rect 124040 16467 124041 16468
rect 124053 16467 124087 16479
rect 124099 16467 124100 16468
rect 124041 16466 124042 16467
rect 124053 16466 124099 16467
rect 123535 15883 123569 16451
rect 124053 15868 124098 16466
rect 124296 16458 124998 16479
rect 125369 16473 125403 16479
rect 124160 16398 124170 16424
rect 124132 16370 124170 16396
rect 124296 16246 124654 16458
rect 124677 16396 124682 16438
rect 124705 16396 124710 16438
rect 124711 15868 124756 16458
rect 125335 16438 125354 16473
rect 125356 16467 125357 16468
rect 125363 16467 125409 16473
rect 125416 16468 125437 16473
rect 125415 16467 125437 16468
rect 126014 16467 126015 16468
rect 126027 16467 126061 16479
rect 126073 16467 126074 16468
rect 125357 16466 125358 16467
rect 125363 16466 125415 16467
rect 125363 16410 125414 16466
rect 125369 15868 125414 16410
rect 125416 16396 125437 16467
rect 126015 16466 126016 16467
rect 126027 16466 126073 16467
rect 126027 15868 126072 16466
rect 126490 16294 127482 16479
rect 127510 16294 127544 16479
rect 127658 16412 131835 16479
rect 127613 16401 131835 16412
rect 127624 16294 131835 16401
rect 126490 16094 131835 16294
rect 126490 16086 127806 16094
rect 124041 15867 124042 15868
rect 124053 15867 124099 15868
rect 124699 15867 124700 15868
rect 124711 15867 124757 15868
rect 125357 15867 125358 15868
rect 125369 15867 125415 15868
rect 126015 15867 126016 15868
rect 126027 15867 126073 15868
rect 126658 15867 126730 16086
rect 126772 15948 126833 16086
rect 126848 15958 127118 16086
rect 127358 16082 127806 16086
rect 126772 15944 126840 15948
rect 124040 15866 124041 15867
rect 123984 15855 124041 15866
rect 124053 15855 124087 15867
rect 124099 15866 124100 15867
rect 124698 15866 124699 15867
rect 124099 15855 124699 15866
rect 124711 15855 124745 15867
rect 124757 15866 124758 15867
rect 125356 15866 125357 15867
rect 124757 15855 124984 15866
rect 125182 15855 125357 15866
rect 125369 15855 125403 15867
rect 125415 15866 125416 15867
rect 126014 15866 126015 15867
rect 125415 15855 126015 15866
rect 126027 15855 126061 15867
rect 126073 15866 126074 15867
rect 126658 15866 126726 15867
rect 126073 15855 126182 15866
rect 126476 15855 126726 15866
rect 126772 15866 126833 15944
rect 127430 15868 127475 16082
rect 127476 15996 127488 16082
rect 127510 16064 127544 16082
rect 127866 16064 127900 16094
rect 128088 16080 128133 16094
rect 128316 16080 131835 16094
rect 127510 16030 127900 16064
rect 127418 15867 127419 15868
rect 127430 15867 127476 15868
rect 127417 15866 127418 15867
rect 126772 15855 127418 15866
rect 127430 15855 127464 15867
rect 127476 15866 127477 15867
rect 127496 15866 127918 15980
rect 127992 15902 131835 16080
rect 128018 15876 128082 15889
rect 127992 15866 128018 15876
rect 128048 15870 128082 15876
rect 128088 15870 128178 15902
rect 128088 15868 128133 15870
rect 128076 15867 128077 15868
rect 128088 15867 128134 15868
rect 128075 15866 128076 15867
rect 127476 15855 127488 15866
rect 127496 15861 128076 15866
rect 128088 15861 128128 15867
rect 128134 15866 128135 15867
rect 128316 15866 131835 15902
rect 128134 15861 131835 15866
rect 127496 15855 128082 15861
rect 128088 15855 128122 15861
rect 128128 15855 131835 15861
rect 123488 15793 123569 15840
rect 123628 15821 131835 15855
rect 124040 15809 124041 15810
rect 124053 15809 124087 15821
rect 124099 15809 124100 15810
rect 124698 15809 124699 15810
rect 124711 15809 124745 15821
rect 124757 15809 124758 15810
rect 125356 15809 125357 15810
rect 125369 15809 125403 15821
rect 125415 15809 125416 15810
rect 126014 15809 126015 15810
rect 126027 15809 126061 15821
rect 126073 15809 126074 15810
rect 126658 15809 126726 15821
rect 124041 15808 124042 15809
rect 124053 15808 124099 15809
rect 124699 15808 124700 15809
rect 124711 15808 124757 15809
rect 125357 15808 125358 15809
rect 125369 15808 125415 15809
rect 126015 15808 126016 15809
rect 126027 15808 126073 15809
rect 123535 15674 123569 15793
rect 124053 15674 124098 15808
rect 124614 15738 124618 15788
rect 124642 15738 124646 15760
rect 124711 15674 124756 15808
rect 125369 15674 125414 15808
rect 126027 15674 126072 15808
rect 117958 15584 118878 15618
rect 115500 14392 116592 14414
rect 115500 14388 116552 14392
rect 111229 13254 111316 13410
rect 111360 13254 111434 13320
rect 111196 13178 111434 13254
rect 104148 13124 107736 13158
rect 110600 13140 110840 13156
rect 111229 13140 111316 13178
rect 103876 11938 103903 12240
rect 104148 11789 104705 13124
rect 104912 11844 104934 12408
rect 99820 11755 104705 11789
rect 106188 11812 106222 13124
rect 106238 13016 106256 13062
rect 106266 12988 106284 13090
rect 106300 13072 106302 13090
rect 106300 13056 106348 13072
rect 106902 13056 106940 13094
rect 107560 13090 107598 13094
rect 106958 13072 106960 13090
rect 106958 13056 107006 13072
rect 107560 13062 107600 13090
rect 107548 13056 107600 13062
rect 106302 13022 106940 13056
rect 106960 13022 107600 13056
rect 106302 12984 106348 13022
rect 106960 12984 107006 13022
rect 107548 13016 107572 13022
rect 107576 12988 107600 13022
rect 106302 12972 106336 12984
rect 106919 12972 106948 12983
rect 106960 12972 106994 12984
rect 107577 12972 107606 12983
rect 107618 12972 107652 13124
rect 106272 11964 106336 12972
rect 106930 11964 106994 12972
rect 107512 11980 107534 12420
rect 106272 11846 106306 11964
rect 106930 11952 106964 11964
rect 107540 11952 107562 12392
rect 107588 11964 107652 12972
rect 107588 11952 107622 11964
rect 106918 11914 106968 11952
rect 107576 11914 107626 11952
rect 106364 11880 106968 11914
rect 107022 11880 107626 11914
rect 107664 11880 107680 11914
rect 106918 11864 106964 11880
rect 107576 11864 107622 11880
rect 106250 11812 106306 11846
rect 106930 11812 106964 11864
rect 107588 11812 107622 11846
rect 107702 11812 107736 13124
rect 110256 13104 110454 13120
rect 110732 13104 110930 13120
rect 111265 13104 111299 13140
rect 111360 13104 111434 13178
rect 110234 13070 112458 13104
rect 110286 13040 110424 13052
rect 110762 13040 110900 13052
rect 110160 13008 110194 13024
rect 110138 12650 110194 13008
rect 110320 13006 110390 13018
rect 110336 13002 110374 13006
rect 110516 13002 110550 13040
rect 110314 12975 110550 13002
rect 110298 12968 110550 12975
rect 110438 12962 110470 12965
rect 110476 12962 110550 12968
rect 110274 12937 110308 12941
rect 110402 12937 110436 12941
rect 110274 12934 110320 12937
rect 110283 12925 110320 12934
rect 110274 12921 110320 12925
rect 110390 12921 110448 12937
rect 110138 12504 110172 12650
rect 110240 12622 110248 12921
rect 110274 12909 110308 12921
rect 110252 12749 110308 12909
rect 110402 12749 110436 12921
rect 110252 12726 110286 12749
rect 110252 12622 110292 12726
rect 110222 12594 110292 12622
rect 110294 12622 110320 12698
rect 110374 12690 110421 12737
rect 110336 12656 110421 12690
rect 110294 12602 110414 12622
rect 110222 12588 110442 12594
rect 110476 12588 110488 12594
rect 110516 12588 110550 12962
rect 110240 12554 110550 12588
rect 110636 13002 110670 13040
rect 110796 13006 110866 13018
rect 110812 13002 110850 13006
rect 110992 13002 111026 13040
rect 110636 12968 111026 13002
rect 110636 12588 110670 12968
rect 110750 12937 110784 12941
rect 110878 12937 110912 12941
rect 110738 12921 110796 12937
rect 110866 12921 110924 12937
rect 110750 12749 110784 12921
rect 110878 12749 110912 12921
rect 110850 12690 110897 12737
rect 110812 12656 110897 12690
rect 110992 12588 111026 12968
rect 110636 12554 111026 12588
rect 110476 12536 110488 12554
rect 110476 12504 110490 12536
rect 110138 11884 110564 12504
rect 110618 11884 111040 12504
rect 106188 11778 109644 11812
rect 99193 11422 99216 11622
rect 99221 11394 99244 11650
rect 99820 11604 101302 11755
rect 99193 11022 99216 11222
rect 99221 10994 99244 11250
rect 99193 10622 99216 10822
rect 99221 10594 99244 10850
rect 99193 10222 99216 10422
rect 99221 10194 99244 10450
rect 99885 9436 99919 11604
rect 100543 9436 100577 11604
rect 101112 11414 101152 11466
rect 101112 11358 101152 11410
rect 101201 9436 101235 11604
rect 101280 11414 101334 11466
rect 101280 11358 101334 11410
rect 102631 9622 102665 11755
rect 104148 11719 104705 11755
rect 106930 9622 106964 11778
rect 107702 9622 107736 11778
rect 110138 10834 110172 11884
rect 111265 11789 111299 13070
rect 111360 13002 111434 13070
rect 112031 13049 112077 13070
rect 112003 13018 112026 13020
rect 112031 13018 112084 13049
rect 112003 13008 112084 13018
rect 112025 13002 112084 13008
rect 112282 13002 112329 13049
rect 111360 12968 112329 13002
rect 111360 12666 111434 12968
rect 112025 12962 112083 12968
rect 112003 12921 112083 12962
rect 111379 11950 111413 12666
rect 112003 11938 112026 12921
rect 112031 11938 112077 12921
rect 112299 12909 112344 12920
rect 112310 11938 112344 12909
rect 112003 11910 112056 11938
rect 112009 11891 112056 11910
rect 112298 11891 112356 11938
rect 111441 11857 112056 11891
rect 112099 11857 112356 11891
rect 112298 11841 112356 11857
rect 112341 11826 112356 11841
rect 112310 11789 112344 11823
rect 112424 11789 112458 13070
rect 113999 11968 114057 11986
rect 114657 11968 114715 11986
rect 113698 11932 114853 11968
rect 116336 11932 116370 14388
rect 117958 14304 117992 15584
rect 118394 15516 118740 15554
rect 118134 15482 118740 15516
rect 118412 15444 118470 15482
rect 118061 15432 118106 15443
rect 118072 14456 118106 15432
rect 118424 14444 118469 15444
rect 118719 15432 118775 15443
rect 118730 14456 118775 15432
rect 118394 14406 118740 14444
rect 118134 14372 118740 14406
rect 118412 14356 118470 14372
rect 118424 14304 118458 14356
rect 118844 14304 118878 15584
rect 119148 15584 119972 15618
rect 119114 15522 119116 15556
rect 118960 15090 118970 15196
rect 119056 15092 119066 15196
rect 117958 14270 118878 14304
rect 119148 14304 119182 15584
rect 119740 15547 119778 15554
rect 119740 15532 119786 15547
rect 119728 15516 119786 15532
rect 119324 15482 119786 15516
rect 119728 15444 119786 15482
rect 119251 15432 119307 15443
rect 119262 14456 119307 15432
rect 119740 14444 119774 15444
rect 119854 14778 119888 15584
rect 121770 15454 121780 15460
rect 119854 14468 119910 14778
rect 119728 14406 119786 14444
rect 119324 14372 119786 14406
rect 119728 14356 119786 14372
rect 119740 14341 119786 14356
rect 119740 14304 119774 14341
rect 119854 14304 119888 14468
rect 119920 14440 119922 15448
rect 121770 15240 121798 15454
rect 119148 14270 119972 14304
rect 117696 12822 117708 13022
rect 117724 12794 117736 13050
rect 117696 12422 117708 12622
rect 117724 12394 117736 12650
rect 118424 11986 118458 14270
rect 116438 11952 116496 11986
rect 117096 11952 117154 11986
rect 117754 11952 117812 11986
rect 118412 11952 118470 11986
rect 119740 11964 119774 14270
rect 116450 11948 116484 11952
rect 117108 11948 117142 11952
rect 113698 11914 119054 11932
rect 113698 11909 117096 11914
rect 117154 11909 117754 11914
rect 117812 11909 118412 11914
rect 118470 11909 119054 11914
rect 113698 11898 117107 11909
rect 117143 11898 117765 11909
rect 117801 11898 118423 11909
rect 118459 11898 119054 11909
rect 113698 11789 114853 11898
rect 111265 11755 114853 11789
rect 116336 11812 116370 11898
rect 116500 11888 117092 11898
rect 117158 11888 117536 11898
rect 116496 11864 117096 11888
rect 117154 11864 117754 11888
rect 117812 11864 118412 11888
rect 118470 11864 118936 11888
rect 119020 11864 119054 11898
rect 119854 11874 119888 14270
rect 121770 13860 121780 15240
rect 123245 15197 126374 15674
rect 126658 15209 126730 15809
rect 126658 15208 126726 15209
rect 126476 15197 126726 15208
rect 126772 15208 126833 15821
rect 127417 15809 127418 15810
rect 127430 15809 127464 15821
rect 127476 15809 127477 15810
rect 127418 15808 127419 15809
rect 127430 15808 127476 15809
rect 127430 15210 127475 15808
rect 127496 15360 127918 15821
rect 127992 15815 128082 15821
rect 128088 15815 128122 15821
rect 128128 15815 128178 15821
rect 128075 15809 128076 15810
rect 128088 15809 128128 15815
rect 128134 15809 128135 15810
rect 128076 15808 128077 15809
rect 128088 15808 128134 15809
rect 128088 15766 128133 15808
rect 128088 15759 128178 15766
rect 128088 15364 128133 15759
rect 128088 15278 128160 15364
rect 127528 15218 127648 15231
rect 128060 15218 128082 15231
rect 128088 15210 128133 15278
rect 127418 15209 127419 15210
rect 127430 15209 127476 15210
rect 128076 15209 128077 15210
rect 128088 15209 128134 15210
rect 127417 15208 127418 15209
rect 126772 15197 127418 15208
rect 127430 15197 127464 15209
rect 127476 15208 127477 15209
rect 128075 15208 128076 15209
rect 127476 15197 127488 15208
rect 127648 15203 128076 15208
rect 127648 15197 128082 15203
rect 128088 15197 128122 15209
rect 128134 15208 128135 15209
rect 128316 15208 131835 15821
rect 128134 15197 131835 15208
rect 123245 15163 131835 15197
rect 123245 14550 126374 15163
rect 126658 15157 126766 15163
rect 126772 15157 126864 15163
rect 126658 15151 126726 15157
rect 126658 15138 126730 15151
rect 126772 15138 126833 15157
rect 127417 15151 127418 15152
rect 127430 15151 127464 15163
rect 127476 15151 127477 15152
rect 128075 15151 128076 15152
rect 128088 15151 128122 15163
rect 128134 15151 128135 15152
rect 127418 15150 127419 15151
rect 127430 15150 127476 15151
rect 128076 15150 128077 15151
rect 128088 15150 128134 15151
rect 126658 15129 126766 15138
rect 126772 15129 126836 15138
rect 126658 15076 126753 15129
rect 126658 14584 126730 15076
rect 126772 14745 126833 15129
rect 127430 14745 127475 15150
rect 128088 14745 128133 15150
rect 126799 14733 126833 14745
rect 128316 14733 131835 15163
rect 126787 14686 127449 14733
rect 127648 14686 131835 14733
rect 126799 14584 126833 14686
rect 126834 14652 127449 14686
rect 127492 14674 128107 14686
rect 128150 14674 131835 14686
rect 127492 14652 131835 14674
rect 128028 14650 131835 14652
rect 128316 14646 131835 14650
rect 127498 14628 127754 14644
rect 127526 14600 127726 14616
rect 128028 14594 131835 14646
rect 128316 14584 131835 14594
rect 126658 14568 131835 14584
rect 131870 14568 131904 18048
rect 192746 17514 192838 18098
rect 193274 17702 193738 18098
rect 193274 17512 193752 17702
rect 193756 17650 193812 17668
rect 193866 17650 193918 17668
rect 141542 15862 141576 17434
rect 149720 16758 149722 17382
rect 149754 16770 149756 17370
rect 193714 17070 193752 17512
rect 193774 17130 193812 17642
rect 193866 17622 193890 17640
rect 193936 17512 194924 18098
rect 142324 16118 142676 16204
rect 142324 16100 143072 16118
rect 149720 16100 149722 16724
rect 149754 16112 149756 16712
rect 141848 16066 149704 16100
rect 195378 16086 196238 18106
rect 196414 16094 197406 18114
rect 197574 17884 199002 18118
rect 197574 17556 199024 17884
rect 142324 16044 143072 16066
rect 142324 15930 142676 16044
rect 140816 15828 144272 15862
rect 141542 15760 141576 15828
rect 141644 15760 141678 15828
rect 142122 15760 142160 15798
rect 142780 15760 142818 15798
rect 143438 15760 143476 15798
rect 144096 15760 144134 15798
rect 141542 15726 142160 15760
rect 142212 15726 142818 15760
rect 142870 15726 143476 15760
rect 143528 15726 144134 15760
rect 141524 15684 141532 15688
rect 141542 15684 141576 15726
rect 141458 15622 141484 15684
rect 141524 15622 141576 15684
rect 126658 14550 132310 14568
rect 123245 14539 126673 14550
rect 126685 14539 126719 14550
rect 126799 14539 126833 14550
rect 123245 14505 126867 14539
rect 128316 14534 132310 14550
rect 123245 13881 126374 14505
rect 126672 14493 126673 14494
rect 126685 14493 126719 14505
rect 126673 14492 126674 14493
rect 126685 14066 126730 14493
rect 126673 13893 126674 13894
rect 126672 13892 126673 13893
rect 126685 13881 126719 14066
rect 126799 13881 126833 14505
rect 127526 14416 127726 14434
rect 127498 14388 127754 14406
rect 123245 13847 126833 13881
rect 123245 13223 126374 13847
rect 126672 13835 126673 13836
rect 126673 13834 126674 13835
rect 126673 13235 126674 13236
rect 126672 13234 126673 13235
rect 126685 13223 126719 13847
rect 126799 13223 126833 13847
rect 128316 13278 131835 14534
rect 123245 13189 126833 13223
rect 120442 12602 120562 12622
rect 120748 12604 120988 13156
rect 123245 13109 126374 13189
rect 126685 13109 126719 13189
rect 126799 13109 126833 13189
rect 127724 13109 131835 13278
rect 123245 13075 131835 13109
rect 120748 12602 121038 12604
rect 120436 12574 120590 12594
rect 120748 12576 120988 12602
rect 120748 12574 121066 12576
rect 120748 12518 120988 12574
rect 123245 12054 126374 13075
rect 124711 11950 124745 12054
rect 118556 11856 118918 11864
rect 119020 11853 119031 11864
rect 119043 11853 119054 11864
rect 124115 11857 124683 11891
rect 116398 11836 118878 11846
rect 116398 11830 118890 11836
rect 118528 11828 118890 11830
rect 119020 11812 119054 11836
rect 124170 11828 124362 11834
rect 124735 11819 124742 11929
rect 124773 11857 124780 11891
rect 126799 11851 126833 13075
rect 127724 13039 131835 13075
rect 131870 13028 131904 14534
rect 139844 14226 139902 14256
rect 139878 14192 139902 14222
rect 137346 14020 137728 14120
rect 136560 13648 137740 14020
rect 141542 14012 141576 15622
rect 141644 15470 141678 15726
rect 141716 15688 141717 15689
rect 141715 15687 141716 15688
rect 142139 15676 142184 15687
rect 142797 15676 142842 15687
rect 143455 15676 143500 15687
rect 144113 15676 144158 15687
rect 142138 15454 142139 15455
rect 142137 15453 142138 15454
rect 142150 15442 142184 15676
rect 142195 15454 142196 15455
rect 142796 15454 142797 15455
rect 142196 15453 142197 15454
rect 142795 15453 142796 15454
rect 142808 15442 142842 15676
rect 142853 15454 142854 15455
rect 143454 15454 143455 15455
rect 142854 15453 142855 15454
rect 143453 15453 143454 15454
rect 143466 15442 143500 15676
rect 143511 15454 143512 15455
rect 144112 15454 144113 15455
rect 143512 15453 143513 15454
rect 144111 15453 144112 15454
rect 144124 15442 144158 15676
rect 144238 15442 144272 15828
rect 148500 15526 148556 15538
rect 149720 15442 149722 16066
rect 149754 15454 149756 16054
rect 195554 15916 195568 16086
rect 195582 15944 195596 16086
rect 141606 15380 141678 15418
rect 141728 15408 144272 15442
rect 142137 15396 142138 15397
rect 142138 15395 142139 15396
rect 141644 14968 141678 15380
rect 142150 14968 142184 15408
rect 142196 15396 142197 15397
rect 142795 15396 142796 15397
rect 142195 15395 142196 15396
rect 142796 15395 142797 15396
rect 142808 14968 142842 15408
rect 142854 15396 142855 15397
rect 143453 15396 143454 15397
rect 142853 15395 142854 15396
rect 143454 15395 143455 15396
rect 143466 14968 143500 15408
rect 143512 15396 143513 15397
rect 144111 15396 144112 15397
rect 143511 15395 143512 15396
rect 144112 15395 144113 15396
rect 141644 14812 141716 14968
rect 142150 14797 142195 14968
rect 142808 14797 142853 14968
rect 143466 14797 143511 14968
rect 142138 14796 142139 14797
rect 142150 14796 142196 14797
rect 142796 14796 142797 14797
rect 142808 14796 142854 14797
rect 143454 14796 143455 14797
rect 143466 14796 143512 14797
rect 144112 14796 144113 14797
rect 142137 14795 142138 14796
rect 141717 14784 142138 14795
rect 142150 14784 142184 14796
rect 142196 14795 142197 14796
rect 142795 14795 142796 14796
rect 142196 14784 142796 14795
rect 142808 14784 142842 14796
rect 142854 14795 142855 14796
rect 143453 14795 143454 14796
rect 142854 14784 143454 14795
rect 143466 14784 143500 14796
rect 143512 14795 143513 14796
rect 144111 14795 144112 14796
rect 143512 14784 143580 14795
rect 144124 14784 144158 15408
rect 144238 14784 144272 15408
rect 148500 15346 148556 15366
rect 148500 15290 148556 15310
rect 149720 14784 149722 15408
rect 149754 14846 149756 15396
rect 149748 14824 149772 14846
rect 149748 14800 149794 14824
rect 149754 14796 149756 14800
rect 141606 14722 141716 14760
rect 141728 14750 144272 14784
rect 142137 14738 142138 14739
rect 142150 14738 142184 14750
rect 142196 14738 142197 14739
rect 142795 14738 142796 14739
rect 142808 14738 142842 14750
rect 142854 14738 142855 14739
rect 143453 14738 143454 14739
rect 143466 14738 143500 14750
rect 143512 14738 143513 14739
rect 144111 14738 144112 14739
rect 142138 14737 142139 14738
rect 142150 14737 142196 14738
rect 142796 14737 142797 14738
rect 142808 14737 142854 14738
rect 143454 14737 143455 14738
rect 143466 14737 143512 14738
rect 144112 14737 144113 14738
rect 141644 14154 141716 14722
rect 142150 14139 142195 14737
rect 142808 14139 142853 14737
rect 143466 14139 143511 14737
rect 142138 14138 142139 14139
rect 142150 14138 142196 14139
rect 142796 14138 142797 14139
rect 142808 14138 142854 14139
rect 143454 14138 143455 14139
rect 143466 14138 143512 14139
rect 144112 14138 144113 14139
rect 142137 14137 142138 14138
rect 141717 14126 142138 14137
rect 142150 14126 142184 14138
rect 142196 14137 142197 14138
rect 142795 14137 142796 14138
rect 142196 14126 142796 14137
rect 142808 14126 142842 14138
rect 142854 14137 142855 14138
rect 143453 14137 143454 14138
rect 142854 14126 143454 14137
rect 143466 14126 143500 14138
rect 143512 14137 143513 14138
rect 144111 14137 144112 14138
rect 143512 14126 143638 14137
rect 144124 14126 144158 14750
rect 144238 14126 144272 14750
rect 149720 14126 149722 14750
rect 149754 14138 149756 14738
rect 194912 14578 194938 15502
rect 194946 14578 194972 15468
rect 196844 14745 196878 16094
rect 197548 14652 197564 14686
rect 197574 14514 199002 17556
rect 141728 14092 144306 14126
rect 142150 14012 142184 14092
rect 142808 14012 142842 14092
rect 143466 14012 143500 14092
rect 144124 14012 144158 14092
rect 144238 14012 144272 14092
rect 141542 13978 149794 14012
rect 138356 13684 139348 13696
rect 139524 13678 140516 13696
rect 132764 13028 133004 13156
rect 139278 13028 139312 13046
rect 127562 12836 127716 12990
rect 128014 12556 128048 12892
rect 128014 12456 128080 12556
rect 128102 12456 128108 12584
rect 128014 12398 128048 12456
rect 128128 12398 128162 12432
rect 127804 12364 128274 12398
rect 128014 12294 128048 12364
rect 128116 12318 128145 12350
rect 128080 12305 128145 12318
rect 128080 12294 128119 12305
rect 128014 12290 128080 12294
rect 128014 12244 128091 12290
rect 128014 12156 128048 12244
rect 128102 12216 128119 12294
rect 128140 12194 128172 12238
rect 128174 12224 128210 12258
rect 128074 12156 128091 12162
rect 128014 12122 128091 12156
rect 128074 12116 128091 12122
rect 128102 12156 128119 12190
rect 128138 12168 128172 12194
rect 128240 12156 128274 12364
rect 128316 12156 130944 13024
rect 131490 12992 131940 13028
rect 132324 12992 132358 13024
rect 132680 12992 132714 13024
rect 132800 12992 132834 13024
rect 133024 12993 133026 13024
rect 132980 12992 133026 12993
rect 131490 12991 133052 12992
rect 131490 12958 133084 12991
rect 131062 12218 131076 12892
rect 128102 12122 130944 12156
rect 116336 11778 119792 11812
rect 128074 11810 128086 12116
rect 128102 12088 128119 12122
rect 128240 12104 128274 12122
rect 128102 11810 128114 12088
rect 128316 12086 130944 12122
rect 128432 11914 128464 12086
rect 128466 11948 128498 12086
rect 124142 11800 124362 11806
rect 112424 10834 112458 11755
rect 113698 11719 114853 11755
rect 117508 11622 117536 11778
rect 118894 11753 118952 11758
rect 119020 10880 119054 11778
rect 131490 11742 131940 12958
rect 132324 12831 132358 12958
rect 132426 12856 132612 12937
rect 132324 12650 132366 12831
rect 132426 12809 132484 12856
rect 132554 12809 132612 12856
rect 132438 12749 132472 12809
rect 132566 12749 132600 12809
rect 132538 12690 132585 12737
rect 132500 12656 132585 12690
rect 132324 12598 132358 12650
rect 132680 12598 132714 12958
rect 132800 12598 132834 12958
rect 133070 12937 133084 12958
rect 132902 12933 132961 12937
rect 133030 12933 133088 12937
rect 132914 12924 132961 12933
rect 132914 12921 132962 12924
rect 132902 12856 132962 12921
rect 132902 12847 132944 12856
rect 132902 12809 132948 12847
rect 132914 12749 132948 12809
rect 132922 12733 132948 12749
rect 132956 12808 132982 12813
rect 132956 12737 132990 12808
rect 133070 12749 133088 12933
rect 132950 12724 133002 12737
rect 132942 12699 133002 12724
rect 132942 12690 132956 12699
rect 132960 12698 133002 12699
rect 132960 12681 133054 12698
rect 132960 12640 133002 12681
rect 133014 12656 133054 12681
rect 132987 12625 133002 12640
rect 132934 12602 132950 12604
rect 132956 12598 132990 12622
rect 133024 12604 133054 12656
rect 132996 12602 133054 12604
rect 132020 12588 132286 12598
rect 132324 12588 132488 12598
rect 132552 12588 132990 12598
rect 133070 12588 133104 12749
rect 133156 12588 133158 13024
rect 134360 12626 134378 12802
rect 132324 12570 132714 12588
rect 132800 12570 133104 12588
rect 132048 12560 132286 12570
rect 132324 12560 133104 12570
rect 132324 12554 132714 12560
rect 132800 12554 133104 12560
rect 133070 12504 133104 12554
rect 132306 12452 132728 12504
rect 132782 12452 133140 12504
rect 132306 12434 133140 12452
rect 132306 12306 133158 12434
rect 132306 11884 132728 12306
rect 132782 11954 133158 12306
rect 135156 12299 135190 12894
rect 135716 12299 135750 12896
rect 135856 12299 136848 13028
rect 137046 12299 138038 13028
rect 138356 12360 139312 13028
rect 139704 12712 139714 13580
rect 142150 13540 142170 13574
rect 141684 13506 142232 13540
rect 141684 13224 141718 13506
rect 142164 13444 142184 13478
rect 141859 13426 142057 13437
rect 142064 13432 142078 13440
rect 141748 13382 141858 13420
rect 141870 13392 142057 13426
rect 142060 13420 142078 13432
rect 142058 13382 142168 13420
rect 141786 13348 141858 13382
rect 141859 13338 142057 13349
rect 141870 13304 142057 13338
rect 142060 13300 142078 13382
rect 142088 13348 142168 13382
rect 142088 13328 142106 13348
rect 142138 13332 142146 13348
rect 142092 13306 142106 13328
rect 142150 13310 142168 13348
rect 142064 13278 142078 13300
rect 142150 13224 142170 13258
rect 142186 13224 142190 13230
rect 142198 13224 142232 13506
rect 141684 13190 142232 13224
rect 142282 13189 142920 13594
rect 139704 12498 139732 12712
rect 139704 12492 139714 12498
rect 138356 12358 139304 12360
rect 138356 12326 139312 12358
rect 139560 12352 139594 12358
rect 139847 12352 140516 13189
rect 140684 12998 143471 13189
rect 140621 12976 143471 12998
rect 140684 12970 143471 12976
rect 140649 12920 143471 12970
rect 140612 12414 140618 12664
rect 139560 12340 140516 12352
rect 140684 12348 143471 12920
rect 144238 12410 144272 13978
rect 207035 13691 207069 21785
rect 207138 21726 207183 21737
rect 207149 13750 207183 21726
rect 207210 13697 207238 21779
rect 207320 21726 207365 21737
rect 207796 21726 207841 21737
rect 207331 13750 207365 21726
rect 207368 17920 207580 17928
rect 207368 17480 207780 17920
rect 207568 17472 207780 17480
rect 207807 13750 207841 21726
rect 207868 13697 207896 21779
rect 207924 13697 207952 21779
rect 207978 21726 208023 21737
rect 208454 21726 208499 21737
rect 207989 13750 208023 21726
rect 208214 17920 208426 17928
rect 208044 17480 208426 17920
rect 208044 17472 208256 17480
rect 208465 13750 208499 21726
rect 208530 13697 208558 21779
rect 208586 13697 208614 21779
rect 208636 21726 208681 21737
rect 209112 21726 209157 21737
rect 208647 13750 208681 21726
rect 208898 17920 208902 17928
rect 208910 17480 208914 17920
rect 209123 13750 209157 21726
rect 209200 13697 209228 21779
rect 209256 13697 209284 21779
rect 209294 21726 209339 21737
rect 209770 21726 209815 21737
rect 209305 13750 209339 21726
rect 209386 17472 209768 17920
rect 209781 13750 209815 21726
rect 209908 13697 209936 21779
rect 209952 21726 209997 21737
rect 209963 13750 209997 21726
rect 210077 17920 210111 21785
rect 212106 21840 212117 21851
rect 212129 21840 212140 21851
rect 212106 21824 212140 21840
rect 212296 21830 212324 21862
rect 212948 21830 212976 21862
rect 213004 21830 213032 21862
rect 213606 21830 213634 21850
rect 213662 21830 213690 21862
rect 214270 21830 214298 21850
rect 214326 21830 214354 21850
rect 214978 21830 215006 21850
rect 215148 21824 215182 21871
rect 212106 21790 215182 21824
rect 210498 18432 210623 18686
rect 210032 17828 210244 17920
rect 210032 17696 210330 17828
rect 210752 17794 210877 18432
rect 211228 17898 211468 18432
rect 210924 17878 211044 17880
rect 211228 17878 211520 17898
rect 211228 17870 211468 17878
rect 210896 17850 211072 17852
rect 211228 17850 211526 17870
rect 211228 17794 211468 17850
rect 211594 17794 211690 18432
rect 211774 17840 211784 17898
rect 210032 17472 210244 17696
rect 211630 17648 211664 17794
rect 211772 17698 211784 17840
rect 211802 17812 211812 17870
rect 211800 17726 211812 17812
rect 210077 13691 210111 17472
rect 211602 17292 211664 17648
rect 211774 17642 211784 17698
rect 211802 17670 211812 17726
rect 206523 13519 206610 13690
rect 207035 13657 210111 13691
rect 211630 13674 211664 17292
rect 212106 13714 212140 21790
rect 212209 21740 212254 21751
rect 212220 13764 212254 21740
rect 212296 17796 212324 21784
rect 212391 21740 212436 21751
rect 212867 21740 212912 21751
rect 212296 17396 212324 17596
rect 212296 13764 212324 17196
rect 212402 13764 212436 21740
rect 212464 17896 212676 17900
rect 212464 17452 212866 17896
rect 212654 17448 212866 17452
rect 212878 13764 212912 21740
rect 212948 13780 212976 21784
rect 213004 13780 213032 21784
rect 213049 21740 213094 21751
rect 213525 21740 213570 21751
rect 213060 13764 213094 21740
rect 213302 17896 213514 17900
rect 213130 17452 213514 17896
rect 213130 17448 213342 17452
rect 213536 13764 213570 21740
rect 213606 13720 213634 21784
rect 213662 13764 213690 21784
rect 213707 21740 213752 21751
rect 214183 21740 214228 21751
rect 213718 13764 213752 21740
rect 213778 17894 213990 17900
rect 213778 17452 214182 17894
rect 213970 17446 214182 17452
rect 214194 13764 214228 21740
rect 214270 13720 214298 21784
rect 214326 13720 214354 21784
rect 214365 21740 214410 21751
rect 214841 21740 214886 21751
rect 214376 13764 214410 21740
rect 214446 17882 214658 17894
rect 214446 17446 214826 17882
rect 214614 17434 214826 17446
rect 214852 13764 214886 21740
rect 214922 20000 214950 21216
rect 214922 13840 214950 15532
rect 214978 13720 215006 21784
rect 215023 21740 215068 21751
rect 215034 13764 215068 21740
rect 215148 13714 215182 21790
rect 215279 14920 215694 21887
rect 217183 21835 217194 21846
rect 217206 21835 217217 21846
rect 217183 21819 217217 21835
rect 218833 21819 218867 21857
rect 217183 21785 218867 21819
rect 216044 20080 216050 21216
rect 216724 14920 216798 15120
rect 215279 14886 215992 14920
rect 215279 14388 215694 14886
rect 215816 14818 215863 14865
rect 215778 14784 215863 14818
rect 215705 14725 215750 14736
rect 215833 14725 215878 14736
rect 215716 14549 215750 14725
rect 215844 14549 215878 14725
rect 215816 14490 215863 14537
rect 215778 14456 215863 14490
rect 215958 14388 215992 14886
rect 215279 14354 215992 14388
rect 216078 14886 216468 14920
rect 216078 14388 216112 14886
rect 216121 14450 216146 14858
rect 216292 14818 216339 14865
rect 216254 14784 216339 14818
rect 216181 14725 216226 14736
rect 216309 14725 216354 14736
rect 216192 14549 216226 14725
rect 216320 14549 216354 14725
rect 216292 14490 216339 14537
rect 216254 14456 216339 14490
rect 216434 14388 216468 14886
rect 216078 14354 216468 14388
rect 216554 14886 216944 14920
rect 216554 14388 216588 14886
rect 216724 14852 216798 14886
rect 216724 14784 216802 14852
rect 216634 14732 216652 14765
rect 216724 14741 216798 14784
rect 216724 14737 216813 14741
rect 216662 14736 216680 14737
rect 216724 14736 216826 14737
rect 216657 14725 216702 14736
rect 216668 14549 216702 14725
rect 216724 14549 216830 14736
rect 216724 14537 216826 14549
rect 216676 14536 216702 14537
rect 216704 14533 216813 14537
rect 216704 14524 216798 14533
rect 216704 14508 216802 14524
rect 216724 14480 216802 14508
rect 216704 14456 216802 14480
rect 216704 14416 216794 14456
rect 216688 14402 216704 14404
rect 216910 14388 216944 14886
rect 216554 14354 216944 14388
rect 215279 14304 215694 14354
rect 215279 13714 216006 14304
rect 211806 13691 216006 13714
rect 216060 13691 216482 14304
rect 216536 13691 216958 14304
rect 211806 13680 216059 13691
rect 216060 13684 216958 13691
rect 217183 13691 217217 21785
rect 217286 21726 217331 21737
rect 217392 21726 217437 21737
rect 217944 21726 217989 21737
rect 218050 21726 218095 21737
rect 218602 21726 218647 21737
rect 218708 21726 218753 21737
rect 217297 21494 217331 21726
rect 217297 20030 217337 21494
rect 217354 20086 217365 21438
rect 217297 13750 217331 20030
rect 217369 14382 217372 15476
rect 217397 14382 217400 15504
rect 217369 14074 217372 14182
rect 217397 14046 217400 14182
rect 217403 13750 217437 21726
rect 217516 17920 217728 17928
rect 217516 17480 217878 17920
rect 217666 17472 217878 17480
rect 217955 15498 217989 21726
rect 218061 21488 218095 21726
rect 218027 20080 218040 21432
rect 218055 20024 218096 21488
rect 217955 13984 217995 15498
rect 217955 13750 217989 13984
rect 218061 13750 218095 20024
rect 218192 17472 218524 17920
rect 218613 13750 218647 21726
rect 218648 20028 218653 21436
rect 218676 20056 218681 21408
rect 218719 15520 218753 21726
rect 218713 14006 218753 15520
rect 218719 13750 218753 14006
rect 218833 17928 218867 21785
rect 219544 18362 219934 18396
rect 218833 17828 219050 17928
rect 219544 17920 219578 18362
rect 219758 18294 219805 18341
rect 219720 18260 219805 18294
rect 219900 18334 219934 18362
rect 219647 18201 219692 18212
rect 219775 18201 219820 18212
rect 219658 18025 219692 18201
rect 219786 18025 219820 18201
rect 219758 17966 219805 18013
rect 219720 17956 219805 17966
rect 219694 17932 219805 17956
rect 219694 17920 219784 17932
rect 219534 17892 219784 17920
rect 219900 17926 219968 18334
rect 219534 17864 219746 17892
rect 219900 17864 219934 17926
rect 220350 17920 220771 21887
rect 222254 21840 222265 21851
rect 222277 21840 222288 21851
rect 222254 21824 222288 21840
rect 223904 21824 223938 21871
rect 222254 21790 223938 21824
rect 219534 17830 219934 17864
rect 220180 17900 220771 17920
rect 218833 17696 219086 17828
rect 219534 17780 219746 17830
rect 220180 17828 220956 17900
rect 218833 17480 219050 17696
rect 218833 13691 218867 17480
rect 219530 17160 219952 17780
rect 220108 17752 220956 17828
rect 221376 17794 221838 18432
rect 220180 17472 220956 17752
rect 220350 17452 220956 17472
rect 221410 17744 221622 17794
rect 221410 17710 221784 17744
rect 221410 17674 221622 17710
rect 221626 17674 221664 17680
rect 221410 17608 221664 17674
rect 207035 13641 207069 13657
rect 207210 13644 207238 13651
rect 207868 13644 207896 13651
rect 207924 13644 207952 13651
rect 208530 13644 208558 13651
rect 208586 13644 208614 13651
rect 209200 13644 209228 13651
rect 209256 13644 209284 13651
rect 209908 13644 209936 13651
rect 207035 13630 207046 13641
rect 207058 13630 207069 13641
rect 210077 13641 210111 13657
rect 212106 13664 212140 13680
rect 213606 13668 213634 13674
rect 212106 13653 212117 13664
rect 212129 13653 212140 13664
rect 214270 13662 214298 13674
rect 214326 13668 214354 13674
rect 214978 13662 215006 13674
rect 215148 13664 215182 13680
rect 215148 13653 215159 13664
rect 215171 13653 215182 13664
rect 215279 13657 216059 13680
rect 216149 13657 216717 13684
rect 217183 13657 218867 13691
rect 210077 13630 210088 13641
rect 210100 13630 210111 13641
rect 215279 13612 215694 13657
rect 217183 13641 217217 13657
rect 217183 13630 217194 13641
rect 217206 13630 217217 13641
rect 218833 13641 218867 13657
rect 218833 13630 218844 13641
rect 218856 13630 218867 13641
rect 211726 13589 215694 13612
rect 220350 13612 220771 17452
rect 221410 17448 221622 17608
rect 221625 17558 221670 17569
rect 221434 17230 221468 17448
rect 221548 17382 221582 17448
rect 221636 17382 221670 17558
rect 221626 17332 221664 17370
rect 221592 17298 221664 17332
rect 221750 17230 221784 17710
rect 221816 17236 221818 17778
rect 222058 17752 222060 17840
rect 221434 17196 221784 17230
rect 222254 13714 222288 21790
rect 222357 21740 222402 21751
rect 222463 21740 222508 21751
rect 223015 21740 223060 21751
rect 223121 21740 223166 21751
rect 223673 21740 223718 21751
rect 223779 21740 223824 21751
rect 222368 21214 222402 21740
rect 222368 19998 222408 21214
rect 222434 20054 222436 21158
rect 222368 13764 222402 19998
rect 222474 13764 222508 21740
rect 222612 17894 222824 17900
rect 222612 17452 222938 17894
rect 222726 17446 222938 17452
rect 223026 15476 223060 21740
rect 223132 21232 223166 21740
rect 223098 20072 223118 21176
rect 223126 20016 223174 21232
rect 223684 21188 223718 21740
rect 223684 20028 223724 21188
rect 223742 20056 223752 21160
rect 223026 13962 223066 15476
rect 223026 13764 223060 13962
rect 223132 13764 223166 20016
rect 223278 17882 223490 17896
rect 223278 17448 223582 17882
rect 223370 17434 223582 17448
rect 223684 13764 223718 20028
rect 223790 15512 223824 21740
rect 223784 13998 223824 15512
rect 223790 13764 223824 13998
rect 223904 13714 223938 21790
rect 224982 14956 225056 15100
rect 224322 14318 224784 14956
rect 224798 14318 225260 14956
rect 226360 14402 226474 14422
rect 226354 14374 226474 14394
rect 225000 14268 225034 14302
rect 224376 14234 224726 14268
rect 224376 14206 224410 14234
rect 224342 14172 224410 14206
rect 224376 13754 224410 14172
rect 224568 14166 224606 14204
rect 224534 14132 224606 14166
rect 224479 14082 224524 14093
rect 224567 14082 224612 14093
rect 224490 13906 224524 14082
rect 224578 13906 224612 14082
rect 224568 13856 224606 13894
rect 224534 13822 224606 13856
rect 224692 13754 224726 14234
rect 224376 13720 224726 13754
rect 224852 14234 225202 14268
rect 224852 13754 224886 14234
rect 224976 14182 225000 14200
rect 225044 14182 225082 14204
rect 224976 14166 225082 14182
rect 224994 14132 225082 14166
rect 224994 14116 225046 14132
rect 225000 14094 225042 14116
rect 225054 14094 225068 14098
rect 224955 14082 224988 14093
rect 225000 14082 225034 14094
rect 224966 14018 225034 14082
rect 225046 14093 225084 14094
rect 224966 13906 225040 14018
rect 225000 13894 225040 13906
rect 225046 13906 225088 14093
rect 225046 13894 225084 13906
rect 225000 13890 225042 13894
rect 224976 13872 225042 13890
rect 225044 13872 225082 13894
rect 224976 13856 225082 13872
rect 224994 13822 225082 13856
rect 224994 13806 225046 13822
rect 225000 13764 225034 13788
rect 225168 13754 225202 14234
rect 224852 13720 225202 13754
rect 222254 13680 224314 13714
rect 224404 13680 224972 13714
rect 222254 13664 222288 13680
rect 222254 13653 222265 13664
rect 222277 13653 222288 13664
rect 223904 13664 223938 13680
rect 223904 13653 223915 13664
rect 223927 13653 223938 13664
rect 220350 13589 225710 13612
rect 206655 13555 210491 13589
rect 211726 13578 225710 13589
rect 215279 13555 220771 13578
rect 215279 13542 215694 13555
rect 220350 13542 220771 13555
rect 144238 12348 144272 12353
rect 140684 12340 144272 12348
rect 139560 12335 144272 12340
rect 138356 12304 139304 12326
rect 139560 12318 144308 12335
rect 139847 12304 144308 12318
rect 138356 12299 144308 12304
rect 144592 12299 144626 13306
rect 144918 12335 148180 13194
rect 144918 12304 148297 12335
rect 148310 12304 148330 12392
rect 148472 12304 148506 13062
rect 205588 12882 205708 12902
rect 205894 12884 206134 13436
rect 205894 12882 206184 12884
rect 205582 12854 205736 12874
rect 205894 12856 206134 12882
rect 205894 12854 206212 12856
rect 205894 12798 206134 12854
rect 212772 12768 212776 13088
rect 212810 12768 212814 13088
rect 149995 12304 153368 12340
rect 144918 12299 153368 12304
rect 134085 12265 138113 12299
rect 138356 12290 153368 12299
rect 132782 11884 133140 11954
rect 133024 11836 133028 11884
rect 132292 11809 132338 11836
rect 132920 11812 133028 11836
rect 132950 11809 132996 11812
rect 132264 11781 132366 11808
rect 132892 11784 133056 11808
rect 132922 11781 133024 11784
rect 134085 11658 134119 12265
rect 134561 12244 134595 12265
rect 134214 12213 135042 12244
rect 135076 12228 135088 12244
rect 135073 12213 135088 12228
rect 134214 12197 135088 12213
rect 135122 12197 135144 12262
rect 135156 12197 135190 12265
rect 135716 12197 135750 12265
rect 137603 12244 137637 12265
rect 137908 12244 137938 12265
rect 135818 12213 135833 12228
rect 135818 12197 135876 12213
rect 136476 12197 136534 12213
rect 137134 12197 137192 12213
rect 137603 12197 137650 12244
rect 137804 12213 137851 12244
rect 137792 12197 137851 12213
rect 137880 12203 137882 12216
rect 137908 12203 137984 12244
rect 137937 12197 137984 12203
rect 134261 12163 137984 12197
rect 134372 12116 134430 12163
rect 134188 12104 134244 12115
rect 134199 11807 134244 12104
rect 134384 11819 134429 12116
rect 134561 11807 134595 12163
rect 135030 12116 135088 12163
rect 134664 12104 134720 12115
rect 134846 12104 134902 12115
rect 134675 11807 134720 12104
rect 134857 11807 134902 12104
rect 135042 11819 135087 12116
rect 134187 11760 135061 11807
rect 134187 11726 134403 11760
rect 134446 11726 135061 11760
rect 134187 11710 134245 11726
rect 134187 11695 134202 11710
rect 134199 11658 134233 11692
rect 134316 11658 134324 11720
rect 134561 11658 134595 11726
rect 134675 11658 134720 11726
rect 134736 11658 134764 11720
rect 134845 11710 134903 11726
rect 134857 11658 134902 11710
rect 135122 11658 135144 12163
rect 135156 11658 135190 12163
rect 135322 12104 135367 12115
rect 122564 11622 122600 11634
rect 133708 11624 135190 11658
rect 122564 11592 122566 11600
rect 122406 11480 122428 11498
rect 122548 11480 122566 11592
rect 131490 11590 131840 11592
rect 122582 11480 122600 11558
rect 122390 11180 122404 11208
rect 122390 10888 122404 11078
rect 122390 10814 122414 10888
rect 123932 10154 125334 10168
rect 118378 9930 118962 9944
rect 126956 9878 129264 11316
rect 129534 9884 131840 11322
rect 131854 10944 131856 11160
rect 131854 10908 131864 10920
rect 131858 10896 131884 10908
rect 131860 10886 131884 10896
rect 127016 9660 127936 9694
rect 127016 9468 127050 9660
rect 127760 9592 127798 9630
rect 127192 9558 127798 9592
rect 127119 9508 127164 9519
rect 127777 9508 127822 9519
rect 127130 9468 127164 9508
rect 127175 9480 127176 9481
rect 127776 9480 127777 9481
rect 127176 9479 127177 9480
rect 127775 9479 127776 9480
rect 127788 9468 127822 9508
rect 127902 9468 127936 9660
rect 59188 9138 62812 9146
rect 59188 9118 59424 9138
rect 59550 9118 62812 9138
rect 59188 9110 62812 9118
rect 59188 9102 59424 9110
rect 59188 9076 59482 9102
rect 47280 6344 47306 6606
rect 47906 6352 50500 7048
rect 47280 6340 47288 6344
rect 47870 6268 47878 6302
rect 22914 5736 23052 5756
rect 22948 5702 23018 5722
rect 23228 5550 23468 6188
rect 47908 6154 50500 6352
rect 18926 5122 22382 5156
rect 20866 4958 20882 5054
rect 20904 4996 20920 5092
rect 20308 4912 20876 4946
rect 22334 4906 22368 5122
rect 22886 5088 22898 5166
rect 22920 5122 22932 5200
rect 58033 4883 58067 9038
rect 59188 9026 59424 9076
rect 58730 9002 58734 9012
rect 59550 9000 62812 9110
rect 58904 8832 58980 8834
rect 58876 8804 59008 8806
rect 58886 8582 58996 8602
rect 58924 8544 58958 8564
rect 99820 7860 101302 9436
rect 127016 9434 127936 9468
rect 127016 8810 127050 9434
rect 127130 8810 127164 9434
rect 127176 9422 127177 9423
rect 127775 9422 127776 9423
rect 127175 9421 127176 9422
rect 127776 9421 127777 9422
rect 127182 9352 127184 9364
rect 127182 9324 127212 9336
rect 127324 9100 127772 9216
rect 127272 9004 127772 9100
rect 127272 8976 127700 9004
rect 127175 8822 127176 8823
rect 127776 8822 127777 8823
rect 127176 8821 127177 8822
rect 127775 8821 127776 8822
rect 127788 8810 127822 9434
rect 127902 8810 127936 9434
rect 128046 9272 128074 9770
rect 131790 9714 131804 9768
rect 134085 9750 134119 11624
rect 134316 9750 134324 11624
rect 134561 9750 134595 11624
rect 134675 9750 134720 11624
rect 134736 9750 134764 11624
rect 134857 9750 134902 11624
rect 135333 9750 135367 12104
rect 135394 11510 135422 12157
rect 135386 11454 135422 11510
rect 135450 11454 135478 12157
rect 135504 12104 135560 12115
rect 135414 11254 135422 11454
rect 135442 11254 135478 11454
rect 135386 11198 135422 11254
rect 135394 9750 135422 11198
rect 128206 9660 129126 9694
rect 128206 9468 128240 9660
rect 128950 9592 128988 9630
rect 128382 9558 128988 9592
rect 128309 9508 128354 9519
rect 128967 9508 129012 9519
rect 128320 9468 128354 9508
rect 128365 9480 128366 9481
rect 128966 9480 128967 9481
rect 128366 9479 128367 9480
rect 128965 9479 128966 9480
rect 128978 9468 129012 9508
rect 129092 9468 129126 9660
rect 128206 9434 129126 9468
rect 128018 9142 128046 9160
rect 128046 9104 128074 9142
rect 128018 9086 128046 9104
rect 127016 8776 127936 8810
rect 127016 8380 127050 8776
rect 127130 8532 127164 8776
rect 127176 8764 127177 8765
rect 127775 8764 127776 8765
rect 127175 8763 127176 8764
rect 127776 8763 127777 8764
rect 127788 8532 127822 8776
rect 127760 8482 127798 8520
rect 127192 8448 127798 8482
rect 127902 8380 127936 8776
rect 127016 8346 127936 8380
rect 128206 8810 128240 9434
rect 128320 8810 128354 9434
rect 128366 9422 128367 9423
rect 128965 9422 128966 9423
rect 128365 9421 128366 9422
rect 128966 9421 128967 9422
rect 128365 8822 128366 8823
rect 128966 8822 128967 8823
rect 128366 8821 128367 8822
rect 128965 8821 128966 8822
rect 128978 8810 129012 9434
rect 129092 8810 129126 9434
rect 128206 8776 129126 8810
rect 128206 8380 128240 8776
rect 128320 8532 128354 8776
rect 128366 8764 128367 8765
rect 128965 8764 128966 8765
rect 128365 8763 128366 8764
rect 128966 8763 128967 8764
rect 128978 8532 129012 8776
rect 128950 8482 128988 8520
rect 128382 8448 128988 8482
rect 129092 8380 129126 8776
rect 128206 8346 129126 8380
rect 129516 9668 130436 9702
rect 129516 9468 129550 9668
rect 130260 9600 130298 9638
rect 129692 9566 130298 9600
rect 129596 9552 129698 9556
rect 130254 9552 130356 9556
rect 129624 9527 129670 9528
rect 130282 9527 130328 9528
rect 129619 9524 129670 9527
rect 130277 9524 130328 9527
rect 129619 9516 129664 9524
rect 130277 9516 130322 9524
rect 129630 9468 129664 9516
rect 129675 9480 129676 9481
rect 130276 9480 130277 9481
rect 129676 9479 129677 9480
rect 130275 9479 130276 9480
rect 130288 9468 130322 9516
rect 130402 9468 130436 9668
rect 129516 9434 130436 9468
rect 129516 8810 129550 9434
rect 129630 8810 129664 9434
rect 129676 9422 129677 9423
rect 130275 9422 130276 9423
rect 129675 9421 129676 9422
rect 130276 9421 130277 9422
rect 129675 8822 129676 8823
rect 130276 8822 130277 8823
rect 129676 8821 129677 8822
rect 130275 8821 130276 8822
rect 130288 8810 130322 9434
rect 130402 8810 130436 9434
rect 129516 8776 130436 8810
rect 128378 8236 128928 8238
rect 128406 8208 128900 8210
rect 129516 8152 129550 8776
rect 129630 8152 129664 8776
rect 129676 8764 129677 8765
rect 130275 8764 130276 8765
rect 129675 8763 129676 8764
rect 130276 8763 130277 8764
rect 130288 8176 130322 8776
rect 130402 8176 130436 8776
rect 130684 9676 131604 9710
rect 130684 9468 130718 9676
rect 131428 9608 131466 9646
rect 130860 9574 131466 9608
rect 130764 9558 130866 9564
rect 130724 9552 130884 9558
rect 131422 9552 131524 9564
rect 130792 9535 130838 9536
rect 131450 9535 131496 9536
rect 130787 9530 130838 9535
rect 130752 9524 130856 9530
rect 131445 9524 131496 9535
rect 130798 9468 130832 9524
rect 130843 9480 130844 9481
rect 131444 9480 131445 9481
rect 130844 9479 130845 9480
rect 131443 9479 131444 9480
rect 131456 9468 131490 9524
rect 131570 9468 131604 9676
rect 130684 9434 131604 9468
rect 130684 8810 130718 9434
rect 130798 8810 130832 9434
rect 130844 9422 130845 9423
rect 131443 9422 131444 9423
rect 130843 9421 130844 9422
rect 131444 9421 131445 9422
rect 130843 8822 130844 8823
rect 131444 8822 131445 8823
rect 130844 8821 130845 8822
rect 131443 8821 131444 8822
rect 131456 8810 131490 9434
rect 131570 8810 131604 9434
rect 130684 8776 131604 8810
rect 129675 8164 129676 8165
rect 129676 8163 129677 8164
rect 130190 8152 130648 8176
rect 123642 8118 130648 8152
rect 129516 8038 129550 8118
rect 129630 8038 129664 8118
rect 130190 8084 130648 8118
rect 130684 8152 130718 8776
rect 130798 8152 130832 8776
rect 130844 8764 130845 8765
rect 131443 8764 131444 8765
rect 130843 8763 130844 8764
rect 131444 8763 131445 8764
rect 130843 8164 130844 8165
rect 131444 8164 131445 8165
rect 130844 8163 130845 8164
rect 131443 8163 131444 8164
rect 131456 8152 131490 8776
rect 131570 8152 131604 8776
rect 130684 8118 131604 8152
rect 130268 8038 130354 8084
rect 130402 8038 130436 8084
rect 130684 8038 130718 8118
rect 130798 8038 130832 8118
rect 131456 8038 131490 8118
rect 131570 8038 131604 8118
rect 123552 8004 131708 8038
rect 131844 8004 131858 9714
rect 132648 8010 132656 9540
rect 58750 7424 59842 7446
rect 68898 7424 69990 7446
rect 58750 7420 59802 7424
rect 68898 7420 69950 7424
rect 63692 5634 63812 5654
rect 63998 5636 64238 6188
rect 63998 5634 64288 5636
rect 63686 5606 63840 5626
rect 63998 5608 64238 5634
rect 63998 5606 64316 5608
rect 63998 5550 64238 5606
rect 64627 5550 64714 6442
rect 73840 5634 73960 5654
rect 74146 5636 74386 6188
rect 74146 5634 74436 5636
rect 85856 5634 85976 5654
rect 86162 5636 86402 6188
rect 86162 5634 86452 5636
rect 73834 5606 73988 5626
rect 74146 5608 74386 5634
rect 74146 5606 74464 5608
rect 85850 5606 86004 5626
rect 86162 5608 86402 5634
rect 86162 5606 86480 5608
rect 74146 5550 74386 5606
rect 86162 5550 86402 5606
rect 99885 4982 99919 7860
rect 100543 4982 100577 7860
rect 101201 4982 101235 7860
rect 129516 7850 129550 8004
rect 130268 7936 130354 8004
rect 130402 7850 130436 8004
rect 130684 7858 130718 8004
rect 131570 7858 131604 8004
rect 124252 7398 124272 7456
rect 124280 7398 124300 7450
rect 124196 7158 124834 7398
rect 124252 6826 124254 7002
rect 124280 6854 124282 6974
rect 132648 6606 132656 7226
rect 133274 7048 133308 9528
rect 133932 7048 133966 9528
rect 133970 7226 133972 8010
rect 134049 7048 135432 9750
rect 135450 7226 135478 11254
rect 135515 10660 135560 12104
rect 135716 11140 135750 12163
rect 135818 12116 135876 12163
rect 135830 12114 135875 12116
rect 135957 12114 136059 12138
rect 136139 12114 136241 12138
rect 136476 12116 136534 12163
rect 136488 12114 136522 12116
rect 136615 12114 136717 12138
rect 136797 12114 136899 12138
rect 137134 12116 137192 12163
rect 137146 12114 137180 12116
rect 137273 12114 137375 12138
rect 137455 12114 137557 12138
rect 137603 12114 137637 12163
rect 137792 12116 137850 12163
rect 137804 12114 137838 12116
rect 137880 12114 137882 12157
rect 137908 12138 137938 12157
rect 137908 12114 138033 12138
rect 138079 12114 138113 12265
rect 135830 12080 138113 12114
rect 139120 12270 153368 12290
rect 139120 12144 139304 12270
rect 139847 12265 148297 12270
rect 139847 12240 143220 12265
rect 139632 12218 139643 12229
rect 139655 12218 139666 12229
rect 139632 12202 139666 12218
rect 139822 12208 143220 12240
rect 143244 12216 143260 12234
rect 143287 12213 143333 12244
rect 139847 12202 143220 12208
rect 139632 12197 143220 12202
rect 143275 12197 143333 12213
rect 139632 12168 143333 12197
rect 139632 12144 139666 12168
rect 139847 12163 143333 12168
rect 139847 12162 143220 12163
rect 139822 12144 143220 12162
rect 139120 12108 143220 12144
rect 143275 12116 143333 12163
rect 135644 11014 135752 11140
rect 135515 7226 135549 10660
rect 135716 8660 135750 11014
rect 135830 10782 135902 12080
rect 135991 11930 136025 12080
rect 136173 12059 136207 12080
rect 136488 12059 136522 12080
rect 136649 12059 136683 12080
rect 136173 12012 136220 12059
rect 136488 12028 136535 12059
rect 136476 12012 136535 12028
rect 136612 12012 136683 12059
rect 136831 12059 136865 12080
rect 137146 12059 137180 12080
rect 137307 12059 137341 12080
rect 136831 12012 136878 12059
rect 137146 12028 137193 12059
rect 137134 12012 137193 12028
rect 137270 12012 137341 12059
rect 137489 12059 137523 12080
rect 137489 12012 137536 12059
rect 137603 12012 137637 12080
rect 137804 12059 137838 12080
rect 137804 12028 137851 12059
rect 137792 12012 137851 12028
rect 137880 12018 137882 12080
rect 137908 12059 137938 12080
rect 137965 12059 137999 12080
rect 137908 12018 137999 12059
rect 137928 12012 137999 12018
rect 136028 11978 136683 12012
rect 136686 11978 137341 12012
rect 137344 11978 137999 12012
rect 135971 11919 136025 11930
rect 135982 11466 136025 11919
rect 136173 11466 136207 11978
rect 136476 11931 136534 11978
rect 135982 11408 136374 11466
rect 136488 11408 136522 11931
rect 136649 11930 136683 11978
rect 136629 11919 136683 11930
rect 135982 11304 136548 11408
rect 135982 11302 136374 11304
rect 135982 10943 136025 11302
rect 135991 10782 136025 10943
rect 136173 10931 136207 11302
rect 136488 10931 136522 11304
rect 136640 11272 136683 11919
rect 136831 11450 136865 11978
rect 137134 11931 137192 11978
rect 136760 11408 136952 11450
rect 137146 11408 137180 11931
rect 137307 11930 137341 11978
rect 137287 11919 137341 11930
rect 136760 11336 137180 11408
rect 136628 11202 136698 11272
rect 136620 10938 136698 11202
rect 136628 10931 136698 10938
rect 136173 10884 136220 10931
rect 136476 10884 136535 10931
rect 136612 10884 136698 10931
rect 136831 10931 136865 11336
rect 136870 11302 137180 11336
rect 137146 10931 137180 11302
rect 137298 10943 137341 11919
rect 137489 11456 137523 11978
rect 137404 11406 137596 11456
rect 137603 11406 137637 11978
rect 137792 11931 137850 11978
rect 137804 11406 137838 11931
rect 137404 11342 137838 11406
rect 137307 10931 137341 10943
rect 136831 10884 136878 10931
rect 137134 10884 137193 10931
rect 137270 10884 137341 10931
rect 137489 10931 137523 11342
rect 137528 11300 137838 11342
rect 137489 10884 137536 10931
rect 137603 10884 137637 11300
rect 137804 10931 137838 11300
rect 137792 10884 137851 10931
rect 137880 10890 137892 11972
rect 137908 11930 137948 11972
rect 137965 11930 137999 11978
rect 137908 11919 137999 11930
rect 137908 11134 137948 11919
rect 137956 11250 137999 11919
rect 137950 11134 138020 11250
rect 137908 10946 138020 11134
rect 137908 10931 137948 10946
rect 137950 10931 138020 10946
rect 137908 10890 138020 10931
rect 137928 10884 138020 10890
rect 136028 10850 137341 10884
rect 137344 10850 138020 10884
rect 136173 10782 136207 10850
rect 136476 10834 136534 10850
rect 136488 10782 136522 10834
rect 136628 10816 136698 10850
rect 136649 10782 136683 10816
rect 136831 10782 136865 10850
rect 137134 10834 137192 10850
rect 137146 10782 137180 10834
rect 137307 10782 137341 10850
rect 137489 10782 137523 10850
rect 137603 10782 137637 10850
rect 137792 10834 137850 10850
rect 137804 10782 137838 10834
rect 137880 10782 137882 10844
rect 137908 10782 137938 10844
rect 137950 10794 138020 10850
rect 137965 10782 137999 10794
rect 138070 10782 138113 12080
rect 135830 10748 138113 10782
rect 135830 10660 135875 10748
rect 135830 8821 135864 10660
rect 135991 8809 136025 10748
rect 136173 8809 136207 10748
rect 136488 8821 136522 10748
rect 136649 8809 136683 10748
rect 136831 9092 136865 10748
rect 137146 9906 137180 10748
rect 137307 9906 137341 10748
rect 137489 9906 137523 10748
rect 137603 9906 137637 10748
rect 137804 9906 137838 10748
rect 137880 9906 137882 10748
rect 137908 9906 137938 10748
rect 137965 9906 137999 10748
rect 138079 9906 138113 10748
rect 138446 12074 143220 12108
rect 138446 12046 138480 12074
rect 138446 10838 138514 12046
rect 139120 12022 143220 12074
rect 139108 12006 143220 12022
rect 138622 11972 143220 12006
rect 139108 11925 143220 11972
rect 138524 11622 138530 11918
rect 138549 11913 138594 11924
rect 138560 10937 138594 11913
rect 138700 11388 138892 11440
rect 139120 11388 143220 11925
rect 138676 11320 143220 11388
rect 139120 10925 143220 11320
rect 139108 10878 143220 10925
rect 138622 10844 143220 10878
rect 138446 10776 138480 10838
rect 139108 10828 143220 10844
rect 139120 10776 143220 10828
rect 138446 10742 143220 10776
rect 139120 10706 143220 10742
rect 139120 9942 139304 10706
rect 139632 9942 139666 10706
rect 139746 10328 139791 10706
rect 139822 10404 143220 10706
rect 143287 10404 143321 12116
rect 143401 10404 143435 12265
rect 144178 12157 144255 12180
rect 144321 12157 144330 12180
rect 144178 12129 144283 12152
rect 144293 12129 144302 12152
rect 143570 10458 143576 11810
rect 143613 10404 143647 10438
rect 139822 10370 144066 10404
rect 139746 9942 139780 10328
rect 139822 10302 143220 10370
rect 143232 10302 143279 10349
rect 139822 10268 143279 10302
rect 143287 10318 143321 10370
rect 143287 10302 143333 10318
rect 143401 10302 143435 10370
rect 143613 10318 143660 10349
rect 143601 10302 143660 10318
rect 143890 10302 143937 10349
rect 143287 10268 143937 10302
rect 138462 9906 138496 9940
rect 139120 9906 139820 9942
rect 136890 9872 139820 9906
rect 136708 8809 136717 9092
rect 136831 8809 136876 9092
rect 136890 9074 136924 9872
rect 137146 9851 137180 9872
rect 137307 9851 137341 9872
rect 137489 9851 137523 9872
rect 137146 9820 137193 9851
rect 137134 9804 137193 9820
rect 137307 9804 137354 9851
rect 137489 9804 137536 9851
rect 137603 9804 137637 9872
rect 137804 9851 137838 9872
rect 137804 9820 137851 9851
rect 137792 9804 137851 9820
rect 137880 9810 137882 9872
rect 137908 9810 137938 9872
rect 137965 9851 137999 9872
rect 137965 9804 138012 9851
rect 138079 9804 138113 9872
rect 138292 9804 138339 9851
rect 138462 9820 138509 9851
rect 138450 9804 138509 9820
rect 138950 9804 138997 9851
rect 139120 9820 139820 9872
rect 139108 9804 139820 9820
rect 137066 9770 137637 9804
rect 137724 9770 138339 9804
rect 138382 9770 138997 9804
rect 139040 9770 139820 9804
rect 137134 9723 137192 9770
rect 136993 9711 137038 9722
rect 137004 9235 137038 9711
rect 137146 9223 137180 9723
rect 137307 9223 137341 9770
rect 137489 9223 137523 9770
rect 137134 9176 137193 9223
rect 137307 9176 137354 9223
rect 137489 9176 137536 9223
rect 137603 9176 137637 9770
rect 137662 9722 137671 9727
rect 137792 9723 137850 9770
rect 137651 9711 137696 9722
rect 137662 9235 137696 9711
rect 137662 9219 137671 9235
rect 137804 9223 137838 9723
rect 137965 9542 137999 9770
rect 138079 9542 138113 9770
rect 138450 9764 138508 9770
rect 139108 9764 139820 9770
rect 138309 9711 138354 9722
rect 137840 9480 138136 9542
rect 137965 9223 137999 9480
rect 137792 9176 137851 9223
rect 137965 9176 138012 9223
rect 138079 9176 138113 9480
rect 138320 9235 138354 9711
rect 138292 9176 138339 9223
rect 138356 9182 138404 9764
rect 138412 9723 138508 9764
rect 138412 9223 138460 9723
rect 138462 9223 138496 9723
rect 139012 9722 139054 9764
rect 138967 9711 139054 9722
rect 138978 9235 139054 9711
rect 138412 9182 138509 9223
rect 138450 9176 138509 9182
rect 138950 9176 138997 9223
rect 139012 9182 139054 9235
rect 139068 9723 139820 9764
rect 139068 9223 139110 9723
rect 139120 9223 139820 9723
rect 139068 9182 139820 9223
rect 139108 9176 139820 9182
rect 137066 9142 137637 9176
rect 137724 9142 138339 9176
rect 138382 9142 138997 9176
rect 139040 9142 139820 9176
rect 137134 9126 137192 9142
rect 137146 9092 137180 9126
rect 137307 9092 137341 9142
rect 137489 9092 137523 9142
rect 137146 9074 137191 9092
rect 137307 9074 137352 9092
rect 137489 9074 137534 9092
rect 137603 9074 137637 9142
rect 137792 9126 137850 9142
rect 137804 9092 137838 9126
rect 137804 9074 137849 9092
rect 137880 9074 137882 9136
rect 137908 9074 137938 9136
rect 137965 9092 137999 9142
rect 137965 9074 138010 9092
rect 138079 9074 138113 9142
rect 138450 9126 138508 9142
rect 139108 9126 139820 9142
rect 138462 9074 138496 9108
rect 139120 9074 139820 9126
rect 136890 9040 139820 9074
rect 137146 8821 137191 9040
rect 137307 8809 137352 9040
rect 137489 8809 137534 9040
rect 137603 8809 137637 9040
rect 137804 8821 137849 9040
rect 137880 8809 137882 9040
rect 137908 8809 137938 9040
rect 137965 8809 138010 9040
rect 135991 8762 136038 8809
rect 136161 8762 136220 8809
rect 136460 8762 136507 8809
rect 136649 8762 136696 8809
rect 136708 8762 138011 8809
rect 135892 8728 136507 8762
rect 136550 8728 137165 8762
rect 137208 8728 137823 8762
rect 137866 8728 138011 8762
rect 135991 8660 136025 8728
rect 136056 8660 136084 8722
rect 136112 8660 136140 8722
rect 136161 8712 136219 8728
rect 136173 8660 136207 8712
rect 136649 8660 136683 8728
rect 136708 8660 136717 8728
rect 136726 8660 136754 8722
rect 136782 8660 136810 8722
rect 136819 8712 136877 8728
rect 136831 8660 136876 8712
rect 137307 8660 137352 8728
rect 137434 8660 137462 8722
rect 137477 8712 137535 8728
rect 137489 8660 137534 8712
rect 137603 8660 137637 8728
rect 137953 8712 138011 8728
rect 137996 8697 138011 8712
rect 137965 8660 137999 8694
rect 138079 8660 138113 9040
rect 139120 9004 139820 9040
rect 139822 9174 143220 10268
rect 143287 10221 143333 10268
rect 143287 10220 143321 10221
rect 143249 10209 143321 10220
rect 143260 9233 143321 10209
rect 143287 9221 143321 9233
rect 143232 9174 143279 9221
rect 139822 9140 143279 9174
rect 143287 9174 143333 9221
rect 143401 9174 143435 10268
rect 143601 10221 143659 10268
rect 143613 9221 143647 10221
rect 143907 10209 143952 10220
rect 143918 9233 143952 10209
rect 143601 9174 143660 9221
rect 143890 9174 143937 9221
rect 143287 9140 143937 9174
rect 139822 9072 143220 9140
rect 143287 9124 143333 9140
rect 143370 9138 143435 9140
rect 143287 9092 143321 9124
rect 143287 9072 143332 9092
rect 143401 9072 143435 9138
rect 143520 9134 143576 9140
rect 143601 9124 143659 9140
rect 143520 9078 143607 9090
rect 143613 9072 143647 9106
rect 143653 9084 143694 9090
rect 143653 9078 143730 9084
rect 144032 9072 144066 10370
rect 144271 9628 144305 9662
rect 139822 9038 144066 9072
rect 144112 9594 144502 9628
rect 144112 9096 144146 9594
rect 144254 9526 144271 9560
rect 144272 9526 144317 9542
rect 144326 9526 144373 9573
rect 144272 9492 144373 9526
rect 144272 9483 144317 9492
rect 144336 9484 144352 9492
rect 144220 9444 144234 9445
rect 144237 9444 144260 9449
rect 144215 9433 144260 9444
rect 144226 9257 144260 9433
rect 144220 9245 144234 9254
rect 144237 9241 144260 9257
rect 144271 9445 144317 9483
rect 144271 9245 144305 9445
rect 144343 9433 144388 9444
rect 144354 9257 144388 9433
rect 144271 9232 144317 9245
rect 144254 9207 144317 9232
rect 144254 9198 144271 9207
rect 144272 9206 144317 9207
rect 144326 9206 144373 9245
rect 144272 9164 144373 9206
rect 144272 9148 144317 9164
rect 144271 9096 144305 9130
rect 144336 9110 144368 9164
rect 144392 9096 144396 9231
rect 144468 9096 144502 9594
rect 144112 9062 144502 9096
rect 144592 9146 144626 12265
rect 144709 12244 144743 12265
rect 144706 12228 144753 12244
rect 144694 12197 144753 12228
rect 144918 12240 148297 12265
rect 148310 12240 148330 12270
rect 144918 12197 148404 12240
rect 144694 12168 148404 12197
rect 144694 12163 148297 12168
rect 144694 12116 144752 12163
rect 144706 9231 144743 12116
rect 144812 12104 144857 12115
rect 144823 9818 144857 12104
rect 144823 9720 144868 9818
rect 144748 9638 144868 9720
rect 144709 9146 144743 9231
rect 144823 9596 144868 9638
rect 144823 9219 144857 9596
rect 144918 9219 148297 12163
rect 148346 12130 148404 12168
rect 144823 9172 144870 9219
rect 144917 9172 148297 9219
rect 144752 9146 148297 9172
rect 144592 9138 148297 9146
rect 144592 9070 144626 9138
rect 144709 9118 144743 9138
rect 144823 9118 144857 9138
rect 144917 9122 148297 9138
rect 144918 9118 148297 9122
rect 144644 9110 148297 9118
rect 144709 9070 144743 9110
rect 144823 9092 144857 9110
rect 144823 9070 144868 9092
rect 144918 9070 148297 9110
rect 138450 8809 138508 8828
rect 138950 8784 139036 8800
rect 139086 8784 139088 8964
rect 139114 8828 139116 8992
rect 139120 8828 139304 9004
rect 139108 8809 139304 8828
rect 139120 8774 139304 8809
rect 138314 8763 138461 8774
rect 138497 8763 138704 8774
rect 138314 8751 138450 8763
rect 138508 8751 138704 8763
rect 138314 8740 138461 8751
rect 138497 8740 138704 8751
rect 138314 8712 138348 8740
rect 138432 8712 138450 8728
rect 138508 8712 138586 8730
rect 138670 8712 138704 8740
rect 138314 8701 138325 8712
rect 138337 8701 138348 8712
rect 138670 8701 138681 8712
rect 138693 8701 138704 8712
rect 138790 8740 139304 8774
rect 138790 8712 138824 8740
rect 138908 8712 139062 8730
rect 138790 8701 138801 8712
rect 138813 8701 138824 8712
rect 138314 8660 138348 8678
rect 138490 8672 138528 8694
rect 138670 8660 138704 8678
rect 138790 8660 138824 8678
rect 138966 8672 139004 8694
rect 139120 8660 139304 8740
rect 135716 8626 139304 8660
rect 135740 8298 135952 8306
rect 135570 7858 135952 8298
rect 135570 7850 135782 7858
rect 135991 7226 136025 8626
rect 136056 7226 136084 8626
rect 136112 7282 136140 8626
rect 135515 7048 135560 7226
rect 132648 6344 132674 6606
rect 133274 6352 135868 7048
rect 132648 6340 132656 6344
rect 133238 6268 133246 6302
rect 108290 5634 108410 5654
rect 108596 5636 108836 6188
rect 133276 6154 135868 6352
rect 134049 6130 135432 6154
rect 108596 5634 108886 5636
rect 108284 5606 108438 5626
rect 108596 5608 108836 5634
rect 108596 5606 108914 5608
rect 108596 5550 108836 5606
rect 13648 4454 13848 4498
rect 13648 4426 13876 4442
rect 134199 4128 134233 6130
rect 134561 4069 134595 6130
rect 134675 5698 134720 6130
rect 134675 4128 134709 5698
rect 134736 4075 134764 6006
rect 134857 5698 134902 6130
rect 135333 5698 135378 6130
rect 134857 4128 134891 5698
rect 135333 4128 135367 5698
rect 135394 4075 135422 6006
rect 135450 4075 135478 6006
rect 135515 5698 135560 6154
rect 135991 6006 136036 7226
rect 136056 6006 136100 7226
rect 135515 4128 135549 5698
rect 135991 4128 136025 6006
rect 136056 4075 136084 6006
rect 136112 5950 136156 7282
rect 136112 4075 136140 5950
rect 136173 4128 136207 8626
rect 136424 8298 136428 8306
rect 136436 7858 136440 8298
rect 136649 4128 136683 8626
rect 136708 8560 136717 8626
rect 136726 4075 136754 8626
rect 136782 4075 136810 8626
rect 136831 8560 136876 8626
rect 137307 8560 137352 8626
rect 136831 4128 136865 8560
rect 136912 7850 137294 8298
rect 137307 4128 137341 8560
rect 137434 4075 137462 8626
rect 137489 8560 137534 8626
rect 137489 4128 137523 8560
rect 137603 8298 137637 8626
rect 137558 8206 137770 8298
rect 137558 8074 137856 8206
rect 137558 7850 137770 8074
rect 137603 4069 137637 7850
rect 134049 3897 134136 4068
rect 134561 4035 137637 4069
rect 134561 4019 134595 4035
rect 134736 4022 134764 4029
rect 135394 4022 135422 4029
rect 135450 4022 135478 4029
rect 136056 4022 136084 4029
rect 136112 4022 136140 4029
rect 136726 4022 136754 4029
rect 136782 4022 136810 4029
rect 137434 4022 137462 4029
rect 134561 4008 134572 4019
rect 134584 4008 134595 4019
rect 137603 4019 137637 4035
rect 138079 4029 138113 8626
rect 138314 8590 138348 8626
rect 138278 8172 138403 8590
rect 138670 8304 138704 8626
rect 138790 8590 138824 8626
rect 139120 8590 139304 8626
rect 138754 8276 138994 8590
rect 138450 8256 138570 8258
rect 138754 8256 139046 8276
rect 138754 8248 138994 8256
rect 138422 8228 138598 8230
rect 138754 8228 139052 8248
rect 138754 8172 138994 8228
rect 139120 8172 139216 8590
rect 139300 8218 139310 8276
rect 139156 8026 139190 8172
rect 139298 8076 139310 8218
rect 139328 8190 139338 8248
rect 139326 8104 139338 8190
rect 139128 7670 139190 8026
rect 139300 8020 139310 8076
rect 139328 8048 139338 8104
rect 139156 4052 139190 7670
rect 139632 4092 139666 9004
rect 139746 8560 139791 9004
rect 139746 4142 139780 8560
rect 139822 8174 143220 9038
rect 139847 7974 143220 8174
rect 139822 7774 143220 7974
rect 139847 7574 143220 7774
rect 139822 5298 143220 7574
rect 143287 8560 143332 9038
rect 143287 5488 143321 8560
rect 143287 5298 143332 5488
rect 143401 5298 143435 9038
rect 144592 9036 148297 9070
rect 144098 8392 144520 9012
rect 144709 7446 144743 9036
rect 144823 8798 144868 9036
rect 144823 8560 144870 8798
rect 144823 8468 144857 8560
rect 144867 8468 144870 8560
rect 144785 8310 144812 8396
rect 144823 8250 144870 8468
rect 144918 8278 148297 9036
rect 148358 8524 148403 12130
rect 148358 8278 148392 8524
rect 148472 8278 148506 12270
rect 149780 12218 149791 12229
rect 149803 12218 149814 12229
rect 149780 12202 149814 12218
rect 149995 12202 153368 12270
rect 149780 12168 153368 12202
rect 148640 10450 148662 11554
rect 144823 7446 144857 8250
rect 144918 7830 148506 8278
rect 144918 7446 148297 7830
rect 144118 7420 148297 7446
rect 144709 7390 144743 7420
rect 144823 7390 144857 7420
rect 144918 7390 148297 7420
rect 144062 7364 148297 7390
rect 144202 5848 144265 5870
rect 144311 5848 144338 5870
rect 144230 5820 144265 5842
rect 144311 5820 144338 5842
rect 144250 5298 144324 5498
rect 139822 5264 143518 5298
rect 139822 4923 143220 5264
rect 143287 5230 143321 5264
rect 143270 5212 143321 5230
rect 143270 5196 143333 5212
rect 143342 5196 143389 5243
rect 143287 5162 143389 5196
rect 143253 5114 143276 5119
rect 143231 5103 143276 5114
rect 143242 4970 143276 5103
rect 143287 5115 143333 5162
rect 143401 5137 143435 5264
rect 143287 4982 143321 5115
rect 143401 5114 143438 5137
rect 143359 5103 143438 5114
rect 143287 4970 143310 4982
rect 143230 4966 143310 4970
rect 143230 4923 143306 4966
rect 143370 4927 143438 5103
rect 139822 4889 143306 4923
rect 139822 4821 143220 4889
rect 143342 4868 143389 4915
rect 143288 4834 143389 4868
rect 143401 4821 143435 4927
rect 139822 4787 143435 4821
rect 139822 4766 143220 4787
rect 143484 4766 143518 5264
rect 139822 4751 143518 4766
rect 139822 4442 139850 4751
rect 139928 4142 139962 4751
rect 140404 4142 140438 4751
rect 140474 4442 140502 4751
rect 140530 4442 140558 4751
rect 140586 4142 140620 4751
rect 141062 4142 141096 4751
rect 141132 4442 141160 4751
rect 141188 4442 141216 4751
rect 141244 4142 141278 4751
rect 141720 4142 141754 4751
rect 141796 4442 141824 4751
rect 141852 4442 141880 4751
rect 141902 4142 141936 4751
rect 142378 4142 142412 4751
rect 142448 4442 142476 4751
rect 142504 4442 142532 4751
rect 142560 4142 142594 4751
rect 142674 4092 142708 4751
rect 142805 4732 143518 4751
rect 143604 5264 143994 5298
rect 143604 4766 143638 5264
rect 143647 4828 143672 5236
rect 143818 5196 143865 5243
rect 143780 5162 143865 5196
rect 143707 5103 143752 5114
rect 143835 5103 143880 5114
rect 143718 4927 143752 5103
rect 143846 4927 143880 5103
rect 143818 4868 143865 4915
rect 143780 4834 143865 4868
rect 143960 4766 143994 5264
rect 143604 4732 143994 4766
rect 144080 5264 144470 5298
rect 144080 4766 144114 5264
rect 144250 5230 144324 5264
rect 144250 5162 144328 5230
rect 144160 5110 144178 5143
rect 144250 5119 144324 5162
rect 144250 5115 144339 5119
rect 144188 5114 144206 5115
rect 144250 5114 144352 5115
rect 144183 5103 144228 5114
rect 144194 4927 144228 5103
rect 144250 4927 144356 5114
rect 144250 4915 144352 4927
rect 144202 4914 144228 4915
rect 144230 4911 144339 4915
rect 144230 4902 144324 4911
rect 144230 4886 144328 4902
rect 144250 4858 144328 4886
rect 144230 4834 144328 4858
rect 144230 4794 144320 4834
rect 144214 4780 144230 4782
rect 144436 4766 144470 5264
rect 144080 4732 144470 4766
rect 142805 4682 143220 4732
rect 142805 4092 143532 4682
rect 139632 4069 143532 4092
rect 143586 4069 144008 4682
rect 144062 4069 144484 4682
rect 144709 4069 144743 7364
rect 144823 4128 144857 7364
rect 144867 4844 144898 5854
rect 144895 4760 144898 4844
rect 144918 4946 148297 7364
rect 148358 4996 148392 7830
rect 148330 4946 148368 4984
rect 144918 4912 148368 4946
rect 144918 4844 148297 4912
rect 148472 4844 148506 7830
rect 148646 6162 148680 6244
rect 148606 5296 148662 5322
rect 148684 4920 148718 9622
rect 148902 8172 149364 8810
rect 148936 8122 149148 8172
rect 148936 8088 149310 8122
rect 148936 8052 149148 8088
rect 149152 8052 149190 8058
rect 148936 7986 149190 8052
rect 148936 7826 149148 7986
rect 149151 7936 149196 7947
rect 148960 7608 148994 7826
rect 149074 7760 149108 7826
rect 149162 7760 149196 7936
rect 149152 7710 149190 7748
rect 149118 7676 149190 7710
rect 149276 7608 149310 8088
rect 149342 7614 149344 8156
rect 149584 8130 149586 8218
rect 148960 7574 149310 7608
rect 149780 6188 149814 12168
rect 149938 12162 153368 12168
rect 149995 12129 153368 12162
rect 149883 12118 149928 12129
rect 149989 12118 153368 12129
rect 149894 11592 149928 12118
rect 149894 10376 149934 11592
rect 149960 10432 149962 11536
rect 148890 5550 149352 6188
rect 149366 5550 149828 6188
rect 149244 5500 149258 5550
rect 148944 5466 149294 5500
rect 148944 4986 148978 5466
rect 149136 5398 149174 5436
rect 149102 5364 149174 5398
rect 149047 5314 149092 5325
rect 149135 5314 149180 5325
rect 149244 5322 149258 5466
rect 149058 5138 149092 5314
rect 149146 5138 149180 5314
rect 149136 5088 149174 5126
rect 149102 5054 149174 5088
rect 149260 4986 149294 5466
rect 148944 4952 149294 4986
rect 149420 5466 149770 5500
rect 149420 4986 149454 5466
rect 149612 5398 149650 5436
rect 149578 5364 149650 5398
rect 149523 5314 149568 5325
rect 149611 5314 149656 5325
rect 149534 5138 149568 5314
rect 149622 5138 149656 5314
rect 149612 5088 149650 5126
rect 149578 5054 149650 5088
rect 149736 4992 149770 5466
rect 149736 4986 149774 4992
rect 149420 4952 149774 4986
rect 144918 4810 148506 4844
rect 148616 4834 148718 4920
rect 144918 4774 148297 4810
rect 144923 4760 144926 4774
rect 144895 4498 144898 4560
rect 144863 4452 144898 4498
rect 144923 4442 144926 4560
rect 144863 4424 144926 4442
rect 144929 4128 144974 4774
rect 145481 4128 145526 4774
rect 145587 4128 145632 4774
rect 145658 4090 145659 4320
rect 146139 4128 146184 4774
rect 146239 4442 146290 4774
rect 146245 4128 146290 4442
rect 146359 4069 146393 4774
rect 139632 4058 143585 4069
rect 143586 4062 146769 4069
rect 139632 4042 139666 4058
rect 139632 4031 139643 4042
rect 139655 4031 139666 4042
rect 142674 4042 142708 4058
rect 142674 4031 142685 4042
rect 142697 4031 142708 4042
rect 142805 4035 143585 4058
rect 143675 4035 144243 4062
rect 144333 4035 146769 4062
rect 137603 4008 137614 4019
rect 137626 4008 137637 4019
rect 142805 3990 143220 4035
rect 144709 4019 144743 4035
rect 144709 4008 144720 4019
rect 144732 4008 144743 4019
rect 146359 4019 146393 4035
rect 146359 4008 146370 4019
rect 146382 4008 146393 4019
rect 139252 3967 143220 3990
rect 147876 3990 148297 4774
rect 148684 4142 148718 4834
rect 149746 4774 149774 4952
rect 149780 4092 149814 5550
rect 149894 4154 149928 10376
rect 149932 8174 149934 8230
rect 149932 7918 149934 7974
rect 149932 7774 149934 7830
rect 149932 7518 149934 7574
rect 149995 6014 153368 12118
rect 153392 11288 153408 12234
rect 149938 5828 149950 5958
rect 149938 5608 149966 5828
rect 149994 5608 153368 6014
rect 149995 5488 153368 5608
rect 153435 5588 153469 9622
rect 154266 7424 155358 7446
rect 154266 7420 155318 7424
rect 159208 5634 159328 5654
rect 159514 5636 159754 6188
rect 159514 5634 159804 5636
rect 159202 5606 159356 5626
rect 159514 5608 159754 5634
rect 159514 5606 159832 5608
rect 149995 5422 153408 5488
rect 149938 4820 149966 5422
rect 149994 5072 153408 5422
rect 149995 4929 153408 5072
rect 153435 5334 153619 5588
rect 159514 5550 159754 5606
rect 153435 4982 153469 5334
rect 149995 4751 153368 4929
rect 153716 4751 153873 5334
rect 153886 4780 154006 4800
rect 154192 4782 154432 5334
rect 154192 4780 154482 4782
rect 153880 4752 154034 4772
rect 154192 4754 154432 4780
rect 154192 4752 154510 4754
rect 149894 4142 149934 4154
rect 150000 4142 150034 4751
rect 150552 4442 150592 4751
rect 150552 4142 150586 4442
rect 150658 4142 150692 4751
rect 151210 4142 151244 4751
rect 151254 4442 151276 4524
rect 151310 4442 151350 4751
rect 151316 4142 151350 4442
rect 149916 4130 149934 4142
rect 149878 4098 149916 4130
rect 149934 4098 149944 4130
rect 151430 4092 151464 4751
rect 151848 4696 152310 4751
rect 152324 4696 152786 4751
rect 154192 4696 154432 4752
rect 152526 4646 152560 4680
rect 151902 4612 152252 4646
rect 151902 4584 151936 4612
rect 151868 4550 151936 4584
rect 151902 4132 151936 4550
rect 152094 4544 152132 4582
rect 152060 4510 152132 4544
rect 152005 4460 152050 4471
rect 152093 4460 152138 4471
rect 152016 4284 152050 4460
rect 152104 4284 152138 4460
rect 152094 4234 152132 4272
rect 152060 4200 152132 4234
rect 152218 4132 152252 4612
rect 151902 4098 152252 4132
rect 152378 4612 152728 4646
rect 152378 4132 152412 4612
rect 152502 4560 152526 4578
rect 152570 4560 152608 4582
rect 152502 4544 152608 4560
rect 152520 4510 152608 4544
rect 152520 4494 152572 4510
rect 152526 4472 152568 4494
rect 152580 4472 152594 4476
rect 152481 4460 152514 4471
rect 152526 4460 152560 4472
rect 152492 4284 152560 4460
rect 152526 4272 152560 4284
rect 152572 4471 152610 4472
rect 152572 4284 152614 4471
rect 152652 4462 152676 4528
rect 152572 4272 152610 4284
rect 152526 4268 152568 4272
rect 152502 4250 152568 4268
rect 152570 4250 152608 4272
rect 152502 4234 152608 4250
rect 152520 4200 152608 4234
rect 152520 4184 152572 4200
rect 152526 4142 152560 4166
rect 152694 4132 152728 4612
rect 153368 4498 153568 4524
rect 153924 4502 153966 4524
rect 154442 4442 154456 4468
rect 152378 4098 152728 4132
rect 149404 4058 151840 4092
rect 151930 4058 152498 4092
rect 149780 4042 149814 4058
rect 149878 4046 149916 4052
rect 149780 4031 149791 4042
rect 149803 4031 149814 4042
rect 149934 4018 149944 4052
rect 151430 4042 151464 4058
rect 151430 4031 151441 4042
rect 151453 4031 151464 4042
rect 147876 3967 153236 3990
rect 134181 3933 138017 3967
rect 139252 3956 153236 3967
rect 142805 3933 148297 3956
rect 142805 3920 143220 3933
rect 147876 3920 148297 3933
rect 133114 3260 133234 3280
rect 133420 3262 133660 3814
rect 133420 3260 133710 3262
rect 133420 3256 133660 3260
rect 132676 3254 133144 3256
rect 133208 3254 133660 3256
rect 133108 3232 133262 3252
rect 133420 3234 133660 3254
rect 133420 3232 133738 3234
rect 133420 3228 133660 3232
rect 132704 3198 133144 3228
rect 133208 3198 133660 3228
rect 133420 3176 133660 3198
rect 140298 3146 140302 3466
rect 140336 3146 140340 3466
<< error_s >>
rect 346562 620583 348166 620633
rect 348174 620583 348374 620633
rect 348463 620617 348663 620667
rect 368090 620625 368290 620675
rect 368379 620591 368579 620641
rect 368587 620591 370191 620641
rect 348829 620499 349153 620549
rect 349219 620517 349419 620567
rect 367334 620525 367534 620575
rect 367600 620507 367924 620557
rect 349039 620365 349153 620415
rect 349305 620383 349419 620433
rect 367334 620391 367448 620441
rect 367600 620373 367714 620423
rect 348783 620261 348897 620311
rect 367856 620269 367970 620319
rect 348783 620061 349139 620111
rect 349205 620061 349405 620111
rect 367348 620069 367548 620119
rect 367614 620069 367970 620119
rect 346562 619931 348166 619981
rect 348178 619931 348378 619981
rect 348463 619931 348663 619981
rect 368090 619939 368290 619989
rect 368375 619939 368575 619989
rect 368587 619939 370191 619989
rect 346154 619549 347474 619599
rect 347608 619549 349212 619599
rect 349220 619549 349420 619599
rect 367333 619557 367533 619607
rect 367541 619557 369145 619607
rect 369279 619557 370599 619607
rect 346154 618897 347446 618947
rect 347608 618897 349212 618947
rect 349224 618897 349424 618947
rect 367329 618905 367529 618955
rect 367541 618905 369145 618955
rect 369307 618905 370599 618955
<< mvpsubdiff >>
rect 345740 628255 345764 629032
rect 371078 628255 371102 629032
<< mvpsubdiffcont >>
rect 345764 628255 371078 629032
<< locali >>
rect 345748 628255 345764 629032
rect 371078 628255 371094 629032
<< viali >>
rect 357593 628300 359298 629000
<< metal1 >>
rect 357470 629399 359442 629457
rect 357470 628057 357538 629399
rect 359388 628057 359442 629399
rect 357470 627990 359442 628057
<< via1 >>
rect 357538 629000 359388 629399
rect 357538 628300 357593 629000
rect 357593 628300 359298 629000
rect 359298 628300 359388 629000
rect 357538 628057 359388 628300
<< metal2 >>
rect 357470 629399 359442 629457
rect 357470 628057 357538 629399
rect 359388 628057 359442 629399
rect 357470 627990 359442 628057
rect 524 -800 636 480
rect 1706 -800 1818 480
rect 2888 -800 3000 480
rect 4070 -800 4182 480
rect 5252 -800 5364 480
rect 6434 -800 6546 480
rect 7616 -800 7728 480
rect 8798 -800 8910 480
rect 9980 -800 10092 480
rect 11162 -800 11274 480
rect 12344 -800 12456 480
rect 13526 -800 13638 480
rect 14708 -800 14820 480
rect 15890 -800 16002 480
rect 17072 -800 17184 480
rect 18254 -800 18366 480
rect 19436 -800 19548 480
rect 20618 -800 20730 480
rect 21800 -800 21912 480
rect 22982 -800 23094 480
rect 24164 -800 24276 480
rect 25346 -800 25458 480
rect 26528 -800 26640 480
rect 27710 -800 27822 480
rect 28892 -800 29004 480
rect 30074 -800 30186 480
rect 31256 -800 31368 480
rect 32438 -800 32550 480
rect 33620 -800 33732 480
rect 34802 -800 34914 480
rect 35984 -800 36096 480
rect 37166 -800 37278 480
rect 38348 -800 38460 480
rect 39530 -800 39642 480
rect 40712 -800 40824 480
rect 41894 -800 42006 480
rect 43076 -800 43188 480
rect 44258 -800 44370 480
rect 45440 -800 45552 480
rect 46622 -800 46734 480
rect 47804 -800 47916 480
rect 48986 -800 49098 480
rect 50168 -800 50280 480
rect 51350 -800 51462 480
rect 52532 -800 52644 480
rect 53714 -800 53826 480
rect 54896 -800 55008 480
rect 56078 -800 56190 480
rect 57260 -800 57372 480
rect 58442 -800 58554 480
rect 59624 -800 59736 480
rect 60806 -800 60918 480
rect 61988 -800 62100 480
rect 63170 -800 63282 480
rect 64352 -800 64464 480
rect 65534 -800 65646 480
rect 66716 -800 66828 480
rect 67898 -800 68010 480
rect 69080 -800 69192 480
rect 70262 -800 70374 480
rect 71444 -800 71556 480
rect 72626 -800 72738 480
rect 73808 -800 73920 480
rect 74990 -800 75102 480
rect 76172 -800 76284 480
rect 77354 -800 77466 480
rect 78536 -800 78648 480
rect 79718 -800 79830 480
rect 80900 -800 81012 480
rect 82082 -800 82194 480
rect 83264 -800 83376 480
rect 84446 -800 84558 480
rect 85628 -800 85740 480
rect 86810 -800 86922 480
rect 87992 -800 88104 480
rect 89174 -800 89286 480
rect 90356 -800 90468 480
rect 91538 -800 91650 480
rect 92720 -800 92832 480
rect 93902 -800 94014 480
rect 95084 -800 95196 480
rect 96266 -800 96378 480
rect 97448 -800 97560 480
rect 98630 -800 98742 480
rect 99812 -800 99924 480
rect 100994 -800 101106 480
rect 102176 -800 102288 480
rect 103358 -800 103470 480
rect 104540 -800 104652 480
rect 105722 -800 105834 480
rect 106904 -800 107016 480
rect 108086 -800 108198 480
rect 109268 -800 109380 480
rect 110450 -800 110562 480
rect 111632 -800 111744 480
rect 112814 -800 112926 480
rect 113996 -800 114108 480
rect 115178 -800 115290 480
rect 116360 -800 116472 480
rect 117542 -800 117654 480
rect 118724 -800 118836 480
rect 119906 -800 120018 480
rect 121088 -800 121200 480
rect 122270 -800 122382 480
rect 123452 -800 123564 480
rect 124634 -800 124746 480
rect 125816 -800 125928 480
rect 126998 -800 127110 480
rect 128180 -800 128292 480
rect 129362 -800 129474 480
rect 130544 -800 130656 480
rect 131726 -800 131838 480
rect 132908 -800 133020 480
rect 134090 -800 134202 480
rect 135272 -800 135384 480
rect 136454 -800 136566 480
rect 137636 -800 137748 480
rect 138818 -800 138930 480
rect 140000 -800 140112 480
rect 141182 -800 141294 480
rect 142364 -800 142476 480
rect 143546 -800 143658 480
rect 144728 -800 144840 480
rect 145910 -800 146022 480
rect 147092 -800 147204 480
rect 148274 -800 148386 480
rect 149456 -800 149568 480
rect 150638 -800 150750 480
rect 151820 -800 151932 480
rect 153002 -800 153114 480
rect 154184 -800 154296 480
rect 155366 -800 155478 480
rect 156548 -800 156660 480
rect 157730 -800 157842 480
rect 158912 -800 159024 480
rect 160094 -800 160206 480
rect 161276 -800 161388 480
rect 162458 -800 162570 480
rect 163640 -800 163752 480
rect 164822 -800 164934 480
rect 166004 -800 166116 480
rect 167186 -800 167298 480
rect 168368 -800 168480 480
rect 169550 -800 169662 480
rect 170732 -800 170844 480
rect 171914 -800 172026 480
rect 173096 -800 173208 480
rect 174278 -800 174390 480
rect 175460 -800 175572 480
rect 176642 -800 176754 480
rect 177824 -800 177936 480
rect 179006 -800 179118 480
rect 180188 -800 180300 480
rect 181370 -800 181482 480
rect 182552 -800 182664 480
rect 183734 -800 183846 480
rect 184916 -800 185028 480
rect 186098 -800 186210 480
rect 187280 -800 187392 480
rect 188462 -800 188574 480
rect 189644 -800 189756 480
rect 190826 -800 190938 480
rect 192008 -800 192120 480
rect 193190 -800 193302 480
rect 194372 -800 194484 480
rect 195554 -800 195666 480
rect 196736 -800 196848 480
rect 197918 -800 198030 480
rect 199100 -800 199212 480
rect 200282 -800 200394 480
rect 201464 -800 201576 480
rect 202646 -800 202758 480
rect 203828 -800 203940 480
rect 205010 -800 205122 480
rect 206192 -800 206304 480
rect 207374 -800 207486 480
rect 208556 -800 208668 480
rect 209738 -800 209850 480
rect 210920 -800 211032 480
rect 212102 -800 212214 480
rect 213284 -800 213396 480
rect 214466 -800 214578 480
rect 215648 -800 215760 480
rect 216830 -800 216942 480
rect 218012 -800 218124 480
rect 219194 -800 219306 480
rect 220376 -800 220488 480
rect 221558 -800 221670 480
rect 222740 -800 222852 480
rect 223922 -800 224034 480
rect 225104 -800 225216 480
rect 226286 -800 226398 480
rect 227468 -800 227580 480
rect 228650 -800 228762 480
rect 229832 -800 229944 480
rect 231014 -800 231126 480
rect 232196 -800 232308 480
rect 233378 -800 233490 480
rect 234560 -800 234672 480
rect 235742 -800 235854 480
rect 236924 -800 237036 480
rect 238106 -800 238218 480
rect 239288 -800 239400 480
rect 240470 -800 240582 480
rect 241652 -800 241764 480
rect 242834 -800 242946 480
rect 244016 -800 244128 480
rect 245198 -800 245310 480
rect 246380 -800 246492 480
rect 247562 -800 247674 480
rect 248744 -800 248856 480
rect 249926 -800 250038 480
rect 251108 -800 251220 480
rect 252290 -800 252402 480
rect 253472 -800 253584 480
rect 254654 -800 254766 480
rect 255836 -800 255948 480
rect 257018 -800 257130 480
rect 258200 -800 258312 480
rect 259382 -800 259494 480
rect 260564 -800 260676 480
rect 261746 -800 261858 480
rect 262928 -800 263040 480
rect 264110 -800 264222 480
rect 265292 -800 265404 480
rect 266474 -800 266586 480
rect 267656 -800 267768 480
rect 268838 -800 268950 480
rect 270020 -800 270132 480
rect 271202 -800 271314 480
rect 272384 -800 272496 480
rect 273566 -800 273678 480
rect 274748 -800 274860 480
rect 275930 -800 276042 480
rect 277112 -800 277224 480
rect 278294 -800 278406 480
rect 279476 -800 279588 480
rect 280658 -800 280770 480
rect 281840 -800 281952 480
rect 283022 -800 283134 480
rect 284204 -800 284316 480
rect 285386 -800 285498 480
rect 286568 -800 286680 480
rect 287750 -800 287862 480
rect 288932 -800 289044 480
rect 290114 -800 290226 480
rect 291296 -800 291408 480
rect 292478 -800 292590 480
rect 293660 -800 293772 480
rect 294842 -800 294954 480
rect 296024 -800 296136 480
rect 297206 -800 297318 480
rect 298388 -800 298500 480
rect 299570 -800 299682 480
rect 300752 -800 300864 480
rect 301934 -800 302046 480
rect 303116 -800 303228 480
rect 304298 -800 304410 480
rect 305480 -800 305592 480
rect 306662 -800 306774 480
rect 307844 -800 307956 480
rect 309026 -800 309138 480
rect 310208 -800 310320 480
rect 311390 -800 311502 480
rect 312572 -800 312684 480
rect 313754 -800 313866 480
rect 314936 -800 315048 480
rect 316118 -800 316230 480
rect 317300 -800 317412 480
rect 318482 -800 318594 480
rect 319664 -800 319776 480
rect 320846 -800 320958 480
rect 322028 -800 322140 480
rect 323210 -800 323322 480
rect 324392 -800 324504 480
rect 325574 -800 325686 480
rect 326756 -800 326868 480
rect 327938 -800 328050 480
rect 329120 -800 329232 480
rect 330302 -800 330414 480
rect 331484 -800 331596 480
rect 332666 -800 332778 480
rect 333848 -800 333960 480
rect 335030 -800 335142 480
rect 336212 -800 336324 480
rect 337394 -800 337506 480
rect 338576 -800 338688 480
rect 339758 -800 339870 480
rect 340940 -800 341052 480
rect 342122 -800 342234 480
rect 343304 -800 343416 480
rect 344486 -800 344598 480
rect 345668 -800 345780 480
rect 346850 -800 346962 480
rect 348032 -800 348144 480
rect 349214 -800 349326 480
rect 350396 -800 350508 480
rect 351578 -800 351690 480
rect 352760 -800 352872 480
rect 353942 -800 354054 480
rect 355124 -800 355236 480
rect 356306 -800 356418 480
rect 357488 -800 357600 480
rect 358670 -800 358782 480
rect 359852 -800 359964 480
rect 361034 -800 361146 480
rect 362216 -800 362328 480
rect 363398 -800 363510 480
rect 364580 -800 364692 480
rect 365762 -800 365874 480
rect 366944 -800 367056 480
rect 368126 -800 368238 480
rect 369308 -800 369420 480
rect 370490 -800 370602 480
rect 371672 -800 371784 480
rect 372854 -800 372966 480
rect 374036 -800 374148 480
rect 375218 -800 375330 480
rect 376400 -800 376512 480
rect 377582 -800 377694 480
rect 378764 -800 378876 480
rect 379946 -800 380058 480
rect 381128 -800 381240 480
rect 382310 -800 382422 480
rect 383492 -800 383604 480
rect 384674 -800 384786 480
rect 385856 -800 385968 480
rect 387038 -800 387150 480
rect 388220 -800 388332 480
rect 389402 -800 389514 480
rect 390584 -800 390696 480
rect 391766 -800 391878 480
rect 392948 -800 393060 480
rect 394130 -800 394242 480
rect 395312 -800 395424 480
rect 396494 -800 396606 480
rect 397676 -800 397788 480
rect 398858 -800 398970 480
rect 400040 -800 400152 480
rect 401222 -800 401334 480
rect 402404 -800 402516 480
rect 403586 -800 403698 480
rect 404768 -800 404880 480
rect 405950 -800 406062 480
rect 407132 -800 407244 480
rect 408314 -800 408426 480
rect 409496 -800 409608 480
rect 410678 -800 410790 480
rect 411860 -800 411972 480
rect 413042 -800 413154 480
rect 414224 -800 414336 480
rect 415406 -800 415518 480
rect 416588 -800 416700 480
rect 417770 -800 417882 480
rect 418952 -800 419064 480
rect 420134 -800 420246 480
rect 421316 -800 421428 480
rect 422498 -800 422610 480
rect 423680 -800 423792 480
rect 424862 -800 424974 480
rect 426044 -800 426156 480
rect 427226 -800 427338 480
rect 428408 -800 428520 480
rect 429590 -800 429702 480
rect 430772 -800 430884 480
rect 431954 -800 432066 480
rect 433136 -800 433248 480
rect 434318 -800 434430 480
rect 435500 -800 435612 480
rect 436682 -800 436794 480
rect 437864 -800 437976 480
rect 439046 -800 439158 480
rect 440228 -800 440340 480
rect 441410 -800 441522 480
rect 442592 -800 442704 480
rect 443774 -800 443886 480
rect 444956 -800 445068 480
rect 446138 -800 446250 480
rect 447320 -800 447432 480
rect 448502 -800 448614 480
rect 449684 -800 449796 480
rect 450866 -800 450978 480
rect 452048 -800 452160 480
rect 453230 -800 453342 480
rect 454412 -800 454524 480
rect 455594 -800 455706 480
rect 456776 -800 456888 480
rect 457958 -800 458070 480
rect 459140 -800 459252 480
rect 460322 -800 460434 480
rect 461504 -800 461616 480
rect 462686 -800 462798 480
rect 463868 -800 463980 480
rect 465050 -800 465162 480
rect 466232 -800 466344 480
rect 467414 -800 467526 480
rect 468596 -800 468708 480
rect 469778 -800 469890 480
rect 470960 -800 471072 480
rect 472142 -800 472254 480
rect 473324 -800 473436 480
rect 474506 -800 474618 480
rect 475688 -800 475800 480
rect 476870 -800 476982 480
rect 478052 -800 478164 480
rect 479234 -800 479346 480
rect 480416 -800 480528 480
rect 481598 -800 481710 480
rect 482780 -800 482892 480
rect 483962 -800 484074 480
rect 485144 -800 485256 480
rect 486326 -800 486438 480
rect 487508 -800 487620 480
rect 488690 -800 488802 480
rect 489872 -800 489984 480
rect 491054 -800 491166 480
rect 492236 -800 492348 480
rect 493418 -800 493530 480
rect 494600 -800 494712 480
rect 495782 -800 495894 480
rect 496964 -800 497076 480
rect 498146 -800 498258 480
rect 499328 -800 499440 480
rect 500510 -800 500622 480
rect 501692 -800 501804 480
rect 502874 -800 502986 480
rect 504056 -800 504168 480
rect 505238 -800 505350 480
rect 506420 -800 506532 480
rect 507602 -800 507714 480
rect 508784 -800 508896 480
rect 509966 -800 510078 480
rect 511148 -800 511260 480
rect 512330 -800 512442 480
rect 513512 -800 513624 480
rect 514694 -800 514806 480
rect 515876 -800 515988 480
rect 517058 -800 517170 480
rect 518240 -800 518352 480
rect 519422 -800 519534 480
rect 520604 -800 520716 480
rect 521786 -800 521898 480
rect 522968 -800 523080 480
rect 524150 -800 524262 480
rect 525332 -800 525444 480
rect 526514 -800 526626 480
rect 527696 -800 527808 480
rect 528878 -800 528990 480
rect 530060 -800 530172 480
rect 531242 -800 531354 480
rect 532424 -800 532536 480
rect 533606 -800 533718 480
rect 534788 -800 534900 480
rect 535970 -800 536082 480
rect 537152 -800 537264 480
rect 538334 -800 538446 480
rect 539516 -800 539628 480
rect 540698 -800 540810 480
rect 541880 -800 541992 480
rect 543062 -800 543174 480
rect 544244 -800 544356 480
rect 545426 -800 545538 480
rect 546608 -800 546720 480
rect 547790 -800 547902 480
rect 548972 -800 549084 480
rect 550154 -800 550266 480
rect 551336 -800 551448 480
rect 552518 -800 552630 480
rect 553700 -800 553812 480
rect 554882 -800 554994 480
rect 556064 -800 556176 480
rect 557246 -800 557358 480
rect 558428 -800 558540 480
rect 559610 -800 559722 480
rect 560792 -800 560904 480
rect 561974 -800 562086 480
rect 563156 -800 563268 480
rect 564338 -800 564450 480
rect 565520 -800 565632 480
rect 566702 -800 566814 480
rect 567884 -800 567996 480
rect 569066 -800 569178 480
rect 570248 -800 570360 480
rect 571430 -800 571542 480
rect 572612 -800 572724 480
rect 573794 -800 573906 480
rect 574976 -800 575088 480
rect 576158 -800 576270 480
rect 577340 -800 577452 480
rect 578522 -800 578634 480
rect 579704 -800 579816 480
rect 580886 -800 580998 480
rect 582068 -800 582180 480
rect 583250 -800 583362 480
<< via2 >>
rect 357538 628057 359388 629399
<< metal3 >>
rect 16194 702300 21194 704800
rect 68194 702300 73194 704800
rect 120194 702300 125194 704800
rect 165594 702300 170594 704800
rect 170894 700788 173094 704800
rect 170894 690603 173094 700738
rect -800 680242 1700 685242
rect 170894 683764 173094 684327
rect 173394 700786 175594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 173394 690603 175594 700736
rect 173394 683764 175594 684327
rect 222594 700836 224794 704800
rect 222594 690636 224794 700786
rect 222594 683913 224794 684360
rect 225094 700846 227294 704800
rect 227594 702300 232594 704800
rect 225094 690636 227294 700796
rect 225094 683913 227294 684360
rect 318994 649497 323994 704800
rect 324294 701130 326494 704800
rect 324294 690618 326494 701080
rect 326794 701150 328994 704800
rect 326794 694292 328994 701100
rect 329294 694292 334294 704800
rect 413394 702300 418394 704800
rect 465394 702300 470394 704800
rect 326794 692092 334294 694292
rect 324294 684038 326494 684344
rect -800 643842 1660 648642
rect 318994 642983 323994 643740
rect 329294 649497 334294 692092
rect 329294 642983 334294 643740
rect 510594 690564 515394 704800
rect -800 633842 1660 638642
rect 510594 637598 515394 684332
rect 510594 631116 515394 631780
rect 520594 690564 525394 704800
rect 566594 702300 571594 704800
rect 520594 637598 525394 684332
rect 582300 677984 584800 682984
rect 560050 639784 560566 644584
rect 566742 639784 584800 644584
rect 520594 631116 525394 631780
rect 560050 629784 560566 634584
rect 566742 629784 584800 634584
rect 357470 629399 359442 629457
rect 357470 628057 357538 629399
rect 359388 628057 359442 629399
rect 357470 627990 359442 628057
rect 339960 620294 345660 620363
rect 371099 620302 533609 620371
rect -800 559442 1660 564242
rect -800 549442 1660 554242
rect 339960 511642 340072 620294
rect 341733 619574 341739 619684
rect 341849 619637 341855 619684
rect 533089 619645 533095 619647
rect 341849 619577 345660 619637
rect 371099 619585 533095 619645
rect 533089 619583 533095 619585
rect 533159 619583 533165 619647
rect 341849 619574 341855 619577
rect 533105 619280 533111 619282
rect -800 511530 340072 511642
rect 340967 619212 345660 619272
rect 371099 619220 533111 619280
rect 533105 619218 533111 619220
rect 533175 619218 533181 619282
rect -800 510348 480 510460
rect -800 509166 480 509278
rect -800 507984 480 508096
rect -800 506802 480 506914
rect -800 505620 480 505732
rect -800 468308 480 468420
rect -800 467126 480 467238
rect -800 465944 480 466056
rect -800 464762 480 464874
rect 340967 463692 341079 619212
rect -800 463580 341079 463692
rect 341738 618632 341850 618638
rect -800 462398 660 462510
rect 780 462398 13894 462510
rect 17564 462398 17711 462510
rect -800 425086 480 425198
rect -800 423904 480 424016
rect -800 422722 480 422834
rect -800 421540 480 421652
rect 341738 420470 341850 618520
rect -800 420358 341850 420470
rect -800 419176 676 419288
rect 738 419176 13887 419288
rect 17599 419176 17694 419288
rect 533497 405408 533609 620302
rect 533894 619647 533958 619653
rect 533958 619585 539606 619645
rect 533894 619577 533958 619583
rect 533904 619282 533968 619288
rect 533968 619220 537488 619280
rect 533904 619212 533968 619218
rect 537376 454558 537488 619220
rect 539494 498980 539606 619585
rect 583520 589472 584800 589584
rect 583520 588290 584800 588402
rect 583520 587108 584800 587220
rect 583520 585926 584800 586038
rect 583520 584744 584800 584856
rect 583520 583562 584800 583674
rect 555452 550562 556229 555362
rect 562346 550562 584800 555362
rect 555452 540562 556229 545362
rect 562346 540562 584800 545362
rect 573371 500050 573548 500162
rect 576743 500050 583220 500162
rect 583318 500050 584800 500162
rect 539494 498868 584800 498980
rect 583520 497686 584800 497798
rect 583520 496504 584800 496616
rect 583520 495322 584800 495434
rect 583520 494140 584800 494252
rect 573405 455628 573556 455740
rect 576731 455628 583180 455740
rect 583296 455628 584800 455740
rect 537376 454446 584800 454558
rect 583520 453264 584800 453376
rect 583520 452082 584800 452194
rect 583520 450900 584800 451012
rect 583520 449718 584800 449830
rect 583520 411206 584800 411318
rect 583520 410024 584800 410136
rect 583520 408842 584800 408954
rect 583520 407660 584800 407772
rect 583520 406478 584800 406590
rect 533497 405296 584800 405408
rect -800 381864 480 381976
rect -800 380682 480 380794
rect -800 379500 480 379612
rect -800 378318 480 378430
rect -800 377136 480 377248
rect -800 375954 480 376066
rect 583520 364784 584800 364896
rect 583520 363602 584800 363714
rect 583520 362420 584800 362532
rect 583520 361238 584800 361350
rect 583520 360056 584800 360168
rect 583520 358874 584800 358986
rect -800 338642 480 338754
rect -800 337460 480 337572
rect -800 336278 480 336390
rect -800 335096 480 335208
rect -800 333914 480 334026
rect -800 332732 480 332844
rect 583520 319562 584800 319674
rect 583520 318380 584800 318492
rect 583520 317198 584800 317310
rect 583520 316016 584800 316128
rect 583520 314834 584800 314946
rect 583520 313652 584800 313764
rect -800 295420 480 295532
rect -800 294238 480 294350
rect -800 293056 480 293168
rect -800 291874 480 291986
rect -800 290692 480 290804
rect -800 289510 480 289622
rect 583520 275140 584800 275252
rect 583520 273958 584800 274070
rect 583520 272776 584800 272888
rect 583520 271594 584800 271706
rect 583520 270412 584800 270524
rect 583520 269230 584800 269342
rect -800 252398 480 252510
rect -800 251216 480 251328
rect -800 250034 480 250146
rect -800 248852 480 248964
rect -800 247670 480 247782
rect -800 246488 480 246600
rect 582340 235230 584800 240030
rect 582340 225230 584800 230030
rect -800 214888 1660 219688
rect -800 204888 1660 209688
rect 13406 191430 13991 196230
rect 17427 191430 573605 196230
rect 576629 191430 584800 196230
rect 582340 181430 584800 186230
rect -800 172888 1660 177688
rect -800 162888 1660 167688
rect 582340 146830 584800 151630
rect 582340 136830 584800 141630
rect -800 124776 480 124888
rect -800 123594 480 123706
rect -800 122412 480 122524
rect -800 121230 480 121342
rect -800 120048 480 120160
rect -800 118866 480 118978
rect 583520 95118 584800 95230
rect 583520 93936 584800 94048
rect 583520 92754 584800 92866
rect 583520 91572 584800 91684
rect -800 81554 480 81666
rect -800 80372 480 80484
rect -800 79190 480 79302
rect -800 78008 480 78120
rect -800 76826 480 76938
rect -800 75644 480 75756
rect 583520 50460 584800 50572
rect 583520 49278 584800 49390
rect 583520 48096 584800 48208
rect 583520 46914 584800 47026
rect -800 38332 480 38444
rect -800 37150 480 37262
rect -800 35968 480 36080
rect -800 34786 480 34898
rect -800 33604 480 33716
rect -800 32422 480 32534
rect 583520 24002 584800 24114
rect 583520 22820 584800 22932
rect 583520 21638 584800 21750
rect 583520 20456 584800 20568
rect 583520 19274 584800 19386
rect 583520 18092 584800 18204
rect -800 16910 480 17022
rect 583520 16910 584800 17022
rect -800 15728 480 15840
rect 583520 15728 584800 15840
rect -800 14546 480 14658
rect 583520 14546 584800 14658
rect -800 13364 480 13476
rect 583520 13364 584800 13476
rect -800 12182 480 12294
rect 583520 12182 584800 12294
rect -800 11000 480 11112
rect 583520 11000 584800 11112
rect -800 9818 480 9930
rect 583520 9818 584800 9930
rect -800 8636 480 8748
rect 583520 8636 584800 8748
rect -800 7454 480 7566
rect 583520 7454 584800 7566
rect -800 6272 480 6384
rect 583520 6272 584800 6384
rect -800 5090 480 5202
rect 583520 5090 584800 5202
rect -800 3908 480 4020
rect 583520 3908 584800 4020
rect -800 2726 480 2838
rect 583520 2726 584800 2838
rect -800 1544 480 1656
rect 583520 1544 584800 1656
<< rmetal3 >>
rect 170894 700738 173094 700788
rect 173394 700736 175594 700786
rect 222594 700786 224794 700836
rect 225094 700796 227294 700846
rect 324294 701080 326494 701130
rect 326794 701100 328994 701150
rect 660 462398 780 462510
rect 676 419176 738 419288
rect 583220 500050 583318 500162
rect 583180 455628 583296 455740
<< via3 >>
rect 170894 684327 173094 690603
rect 173394 684327 175594 690603
rect 222594 684360 224794 690636
rect 225094 684360 227294 690636
rect 324294 684344 326494 690618
rect 318994 643740 323994 649497
rect 329294 643740 334294 649497
rect 510594 684332 515394 690564
rect 510594 631780 515394 637598
rect 520594 684332 525394 690564
rect 560566 639784 566742 644584
rect 520594 631780 525394 637598
rect 560566 629784 566742 634584
rect 357538 628057 359388 629399
rect 341739 619574 341849 619684
rect 533095 619583 533159 619647
rect 533111 619218 533175 619282
rect 341738 618520 341850 618632
rect 13894 462398 17564 462510
rect 13887 419176 17599 419288
rect 533894 619583 533958 619647
rect 533904 619218 533968 619282
rect 556229 550562 562346 555362
rect 556229 540562 562346 545362
rect 573548 500050 576743 500162
rect 573556 455628 576731 455740
rect 13991 191430 17427 196230
rect 573605 191430 576629 196230
<< metal4 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
rect 170628 690636 526162 690737
rect 170628 690603 222594 690636
rect 170628 684327 170894 690603
rect 173094 684327 173394 690603
rect 175594 684360 222594 690603
rect 224794 684360 225094 690636
rect 227294 690618 526162 690636
rect 227294 684360 324294 690618
rect 175594 684344 324294 684360
rect 326494 690564 526162 690618
rect 326494 684344 510594 690564
rect 175594 684332 510594 684344
rect 515394 684332 520594 690564
rect 525394 684332 526162 690564
rect 175594 684327 526162 684332
rect 170628 684183 526162 684327
rect 318330 649837 359973 649898
rect 318330 649497 357559 649837
rect 318330 643740 318994 649497
rect 323994 643740 329294 649497
rect 334294 643740 357559 649497
rect 318330 643394 357559 643740
rect 359314 643394 359973 649837
rect 318330 643344 359973 643394
rect 560425 644584 566979 644980
rect 560425 639784 560566 644584
rect 566742 639784 566979 644584
rect 356144 637598 525696 637898
rect 356144 631780 510594 637598
rect 515394 631780 520594 637598
rect 525394 631780 525696 637598
rect 356144 631344 525696 631780
rect 560425 634584 566979 639784
rect 357442 629399 359470 631344
rect 357442 628057 357538 629399
rect 359388 628057 359470 629399
rect 357442 619873 359470 628057
rect 560425 629784 560566 634584
rect 566742 629784 566979 634584
rect 341738 619684 341850 619685
rect 341738 619574 341739 619684
rect 341849 619574 341850 619684
rect 341738 618633 341850 619574
rect 356867 619473 359885 619873
rect 533094 619647 533160 619648
rect 533094 619583 533095 619647
rect 533159 619645 533160 619647
rect 533893 619647 533959 619648
rect 533893 619645 533894 619647
rect 533159 619585 533894 619645
rect 533159 619583 533160 619585
rect 533094 619582 533160 619583
rect 533893 619583 533894 619585
rect 533958 619583 533959 619647
rect 533893 619582 533959 619583
rect 533110 619282 533176 619283
rect 533110 619218 533111 619282
rect 533175 619280 533176 619282
rect 533903 619282 533969 619283
rect 533903 619280 533904 619282
rect 533175 619220 533904 619280
rect 533175 619218 533176 619220
rect 533110 619217 533176 619218
rect 533903 619218 533904 619220
rect 533968 619218 533969 619282
rect 533903 619217 533969 619218
rect 341737 618632 341851 618633
rect 341737 618520 341738 618632
rect 341850 618520 341851 618632
rect 341737 618519 341851 618520
rect 345773 613756 346828 618849
rect 351928 617829 353757 618856
rect 351928 615249 352028 617829
rect 353603 615249 353757 617829
rect 351928 615131 353757 615249
rect 363328 617835 365157 618884
rect 363328 615255 363412 617835
rect 364987 615255 365157 617835
rect 363328 615131 365157 615255
rect 369823 613756 370980 618859
rect 560425 613756 566979 629784
rect 345256 607202 566979 613756
rect 362658 601572 562613 601756
rect 362658 597231 363414 601572
rect 364992 597231 562613 601572
rect 362658 595202 562613 597231
rect 556059 555362 562613 595202
rect 556059 550562 556229 555362
rect 562346 550562 562613 555362
rect 556059 545362 562613 550562
rect 556059 540562 556229 545362
rect 562346 540562 562613 545362
rect 556059 540155 562613 540562
rect 573464 500162 576816 500473
rect 573464 500050 573548 500162
rect 576743 500050 576816 500162
rect 13814 462510 17684 462771
rect 13814 462398 13894 462510
rect 17564 462398 17684 462510
rect 13814 419288 17684 462398
rect 13814 419176 13887 419288
rect 17599 419176 17684 419288
rect 13814 227257 17684 419176
rect 573464 455740 576816 500050
rect 573464 455628 573556 455740
rect 576731 455628 576816 455740
rect 13811 196230 17688 227257
rect 13811 191430 13991 196230
rect 17427 191430 17688 196230
rect 13811 191098 17688 191430
rect 573464 196230 576816 455628
rect 573464 191430 573605 196230
rect 576629 191430 576816 196230
rect 573464 191191 576816 191430
<< via4 >>
rect 357559 643394 359314 649837
rect 352028 615249 353603 617829
rect 363412 615255 364987 617835
rect 363414 597231 364992 601572
<< metal5 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
rect 357521 649837 359350 649991
rect 357521 643394 357559 649837
rect 359314 643394 359350 649837
rect 351918 617829 353747 617929
rect 351918 615249 352028 617829
rect 353603 615249 353747 617829
rect 351918 614900 353747 615249
rect 357521 614900 359350 643394
rect 351918 613071 359350 614900
rect 363318 617835 365147 617929
rect 363318 615255 363412 617835
rect 364987 615255 365147 617835
rect 363318 601572 365147 615255
rect 363318 597231 363414 601572
rect 364992 597231 365147 601572
rect 363318 597052 365147 597231
<< comment >>
rect -100 704000 584100 704100
rect -100 0 0 704000
rect 584000 0 584100 704000
rect -100 -100 584100 0
use ColROs  ColROs_0
timestamp 1695461588
transform 1 0 47061 0 1 9739
box -33468 -9022 186662 48942
use sky130_fd_pr__res_generic_m3_DPAT6Q  R1
timestamp 0
transform 1 0 1100 0 1 687
box 0 0 1 1
use sky130_fd_pr__res_generic_m3_DPAT6Q  R2
timestamp 0
transform 1 0 3300 0 1 687
box 0 0 1 1
use sky130_fd_pr__res_generic_m3_DPAT6Q  R4
timestamp 0
transform 1 0 5500 0 1 687
box 0 0 1 1
use sky130_fd_pr__res_generic_m3_DPAT6Q  R5
timestamp 0
transform 1 0 7700 0 1 687
box 0 0 1 1
use sky130_fd_pr__res_generic_m3_DPAT6Q  R6
timestamp 0
transform 1 0 9900 0 1 687
box 0 0 1 1
use sky130_fd_pr__res_generic_m3_DPAT6Q  R7
timestamp 0
transform 1 0 12100 0 1 687
box 0 0 1 1
use sky130_fd_pr__res_generic_m3_2QNVX3  R8
timestamp 0
transform 1 0 13256 0 1 706
box 0 0 1 1
use sky130_fd_pr__res_generic_m3_SS5VKG  R9
timestamp 0
transform 1 0 13368 0 1 688
box 0 0 1 1
use sky130_fd_pr__res_generic_m3_HK2ST4  R11
timestamp 0
transform 1 0 13480 0 1 715
box 0 0 1 1
use sky130_fd_pr__res_generic_m3_BHQV68  R12
timestamp 0
transform 1 0 13592 0 1 717
box 0 0 1 1
use user_analog_proj_example  user_analog_proj_example_0 /run/media/thuat/build/cmos/MulColRO/mag
timestamp 1639841760
transform 1 0 345668 0 -1 627114
box -59 -22 25476 8324
use ColROs  x3
timestamp 1695461588
transform 1 0 41048 0 1 9622
box -33468 -9022 186662 48942
<< labels >>
flabel metal3 s 583520 269230 584800 269342 0 FreeSans 1120 0 0 0 gpio_analog[0]
port 0 nsew signal bidirectional
flabel metal3 s -800 381864 480 381976 0 FreeSans 1120 0 0 0 gpio_analog[10]
port 1 nsew signal bidirectional
flabel metal3 s -800 338642 480 338754 0 FreeSans 1120 0 0 0 gpio_analog[11]
port 2 nsew signal bidirectional
flabel metal3 s -800 295420 480 295532 0 FreeSans 1120 0 0 0 gpio_analog[12]
port 3 nsew signal bidirectional
flabel metal3 s -800 252398 480 252510 0 FreeSans 1120 0 0 0 gpio_analog[13]
port 4 nsew signal bidirectional
flabel metal3 s -800 124776 480 124888 0 FreeSans 1120 0 0 0 gpio_analog[14]
port 5 nsew signal bidirectional
flabel metal3 s -800 81554 480 81666 0 FreeSans 1120 0 0 0 gpio_analog[15]
port 6 nsew signal bidirectional
flabel metal3 s -800 38332 480 38444 0 FreeSans 1120 0 0 0 gpio_analog[16]
port 7 nsew signal bidirectional
flabel metal3 s -800 16910 480 17022 0 FreeSans 1120 0 0 0 gpio_analog[17]
port 8 nsew signal bidirectional
flabel metal3 s 583520 313652 584800 313764 0 FreeSans 1120 0 0 0 gpio_analog[1]
port 9 nsew signal bidirectional
flabel metal3 s 583520 358874 584800 358986 0 FreeSans 1120 0 0 0 gpio_analog[2]
port 10 nsew signal bidirectional
flabel metal3 s 583520 405296 584800 405408 0 FreeSans 1120 0 0 0 gpio_analog[3]
port 11 nsew signal bidirectional
flabel metal3 s 583520 449718 584800 449830 0 FreeSans 1120 0 0 0 gpio_analog[4]
port 12 nsew signal bidirectional
flabel metal3 s 583520 494140 584800 494252 0 FreeSans 1120 0 0 0 gpio_analog[5]
port 13 nsew signal bidirectional
flabel metal3 s 583520 583562 584800 583674 0 FreeSans 1120 0 0 0 gpio_analog[6]
port 14 nsew signal bidirectional
flabel metal3 s -800 511530 480 511642 0 FreeSans 1120 0 0 0 gpio_analog[7]
port 15 nsew signal bidirectional
flabel metal3 s -800 468308 480 468420 0 FreeSans 1120 0 0 0 gpio_analog[8]
port 16 nsew signal bidirectional
flabel metal3 s -800 425086 480 425198 0 FreeSans 1120 0 0 0 gpio_analog[9]
port 17 nsew signal bidirectional
flabel metal3 s 583520 270412 584800 270524 0 FreeSans 1120 0 0 0 gpio_noesd[0]
port 18 nsew signal bidirectional
flabel metal3 s -800 380682 480 380794 0 FreeSans 1120 0 0 0 gpio_noesd[10]
port 19 nsew signal bidirectional
flabel metal3 s -800 337460 480 337572 0 FreeSans 1120 0 0 0 gpio_noesd[11]
port 20 nsew signal bidirectional
flabel metal3 s -800 294238 480 294350 0 FreeSans 1120 0 0 0 gpio_noesd[12]
port 21 nsew signal bidirectional
flabel metal3 s -800 251216 480 251328 0 FreeSans 1120 0 0 0 gpio_noesd[13]
port 22 nsew signal bidirectional
flabel metal3 s -800 123594 480 123706 0 FreeSans 1120 0 0 0 gpio_noesd[14]
port 23 nsew signal bidirectional
flabel metal3 s -800 80372 480 80484 0 FreeSans 1120 0 0 0 gpio_noesd[15]
port 24 nsew signal bidirectional
flabel metal3 s -800 37150 480 37262 0 FreeSans 1120 0 0 0 gpio_noesd[16]
port 25 nsew signal bidirectional
flabel metal3 s -800 15728 480 15840 0 FreeSans 1120 0 0 0 gpio_noesd[17]
port 26 nsew signal bidirectional
flabel metal3 s 583520 314834 584800 314946 0 FreeSans 1120 0 0 0 gpio_noesd[1]
port 27 nsew signal bidirectional
flabel metal3 s 583520 360056 584800 360168 0 FreeSans 1120 0 0 0 gpio_noesd[2]
port 28 nsew signal bidirectional
flabel metal3 s 583520 406478 584800 406590 0 FreeSans 1120 0 0 0 gpio_noesd[3]
port 29 nsew signal bidirectional
flabel metal3 s 583520 450900 584800 451012 0 FreeSans 1120 0 0 0 gpio_noesd[4]
port 30 nsew signal bidirectional
flabel metal3 s 583520 495322 584800 495434 0 FreeSans 1120 0 0 0 gpio_noesd[5]
port 31 nsew signal bidirectional
flabel metal3 s 583520 584744 584800 584856 0 FreeSans 1120 0 0 0 gpio_noesd[6]
port 32 nsew signal bidirectional
flabel metal3 s -800 510348 480 510460 0 FreeSans 1120 0 0 0 gpio_noesd[7]
port 33 nsew signal bidirectional
flabel metal3 s -800 467126 480 467238 0 FreeSans 1120 0 0 0 gpio_noesd[8]
port 34 nsew signal bidirectional
flabel metal3 s -800 423904 480 424016 0 FreeSans 1120 0 0 0 gpio_noesd[9]
port 35 nsew signal bidirectional
flabel metal3 s 582300 677984 584800 682984 0 FreeSans 1120 0 0 0 io_analog[0]
port 36 nsew signal bidirectional
flabel metal3 s 0 680242 1700 685242 0 FreeSans 1120 0 0 0 io_analog[10]
port 37 nsew signal bidirectional
flabel metal3 s 566594 702300 571594 704800 0 FreeSans 1920 180 0 0 io_analog[1]
port 38 nsew signal bidirectional
flabel metal3 s 465394 702300 470394 704800 0 FreeSans 1920 180 0 0 io_analog[2]
port 39 nsew signal bidirectional
flabel metal3 s 413394 702300 418394 704800 0 FreeSans 1920 180 0 0 io_analog[3]
port 40 nsew signal bidirectional
flabel metal3 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal4 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal5 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal3 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal4 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal5 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal3 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal4 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal5 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal3 s 120194 702300 125194 704800 0 FreeSans 1920 180 0 0 io_analog[7]
port 44 nsew signal bidirectional
flabel metal3 s 68194 702300 73194 704800 0 FreeSans 1920 180 0 0 io_analog[8]
port 45 nsew signal bidirectional
flabel metal3 s 16194 702300 21194 704800 0 FreeSans 1920 180 0 0 io_analog[9]
port 46 nsew signal bidirectional
flabel metal3 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal4 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal5 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal3 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal4 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal5 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal3 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal4 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal5 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal3 s 326794 702300 328994 704800 0 FreeSans 1920 180 0 0 io_clamp_high[0]
port 50 nsew signal bidirectional
flabel metal3 s 225094 702300 227294 704800 0 FreeSans 1920 180 0 0 io_clamp_high[1]
port 51 nsew signal bidirectional
flabel metal3 s 173394 702300 175594 704800 0 FreeSans 1920 180 0 0 io_clamp_high[2]
port 52 nsew signal bidirectional
flabel metal3 s 324294 702300 326494 704800 0 FreeSans 1920 180 0 0 io_clamp_low[0]
port 53 nsew signal bidirectional
flabel metal3 s 222594 702300 224794 704800 0 FreeSans 1920 180 0 0 io_clamp_low[1]
port 54 nsew signal bidirectional
flabel metal3 s 170894 702300 173094 704800 0 FreeSans 1920 180 0 0 io_clamp_low[2]
port 55 nsew signal bidirectional
flabel metal3 s 583520 2726 584800 2838 0 FreeSans 1120 0 0 0 io_in[0]
port 56 nsew signal input
flabel metal3 s 583520 408842 584800 408954 0 FreeSans 1120 0 0 0 io_in[10]
port 57 nsew signal input
flabel metal3 s 583520 453264 584800 453376 0 FreeSans 1120 0 0 0 io_in[11]
port 58 nsew signal input
flabel metal3 s 583520 497686 584800 497798 0 FreeSans 1120 0 0 0 io_in[12]
port 59 nsew signal input
flabel metal3 s 583520 587108 584800 587220 0 FreeSans 1120 0 0 0 io_in[13]
port 60 nsew signal input
flabel metal3 s -800 507984 480 508096 0 FreeSans 1120 0 0 0 io_in[14]
port 61 nsew signal input
flabel metal3 s -800 464762 480 464874 0 FreeSans 1120 0 0 0 io_in[15]
port 62 nsew signal input
flabel metal3 s -800 421540 480 421652 0 FreeSans 1120 0 0 0 io_in[16]
port 63 nsew signal input
flabel metal3 s -800 378318 480 378430 0 FreeSans 1120 0 0 0 io_in[17]
port 64 nsew signal input
flabel metal3 s -800 335096 480 335208 0 FreeSans 1120 0 0 0 io_in[18]
port 65 nsew signal input
flabel metal3 s -800 291874 480 291986 0 FreeSans 1120 0 0 0 io_in[19]
port 66 nsew signal input
flabel metal3 s 583520 7454 584800 7566 0 FreeSans 1120 0 0 0 io_in[1]
port 67 nsew signal input
flabel metal3 s -800 248852 480 248964 0 FreeSans 1120 0 0 0 io_in[20]
port 68 nsew signal input
flabel metal3 s -800 121230 480 121342 0 FreeSans 1120 0 0 0 io_in[21]
port 69 nsew signal input
flabel metal3 s -800 78008 480 78120 0 FreeSans 1120 0 0 0 io_in[22]
port 70 nsew signal input
flabel metal3 s -800 34786 480 34898 0 FreeSans 1120 0 0 0 io_in[23]
port 71 nsew signal input
flabel metal3 s -800 13364 480 13476 0 FreeSans 1120 0 0 0 io_in[24]
port 72 nsew signal input
flabel metal3 s -800 8636 480 8748 0 FreeSans 1120 0 0 0 io_in[25]
port 73 nsew signal input
flabel metal3 s -800 3908 480 4020 0 FreeSans 1120 0 0 0 io_in[26]
port 74 nsew signal input
flabel metal3 s 583520 12182 584800 12294 0 FreeSans 1120 0 0 0 io_in[2]
port 75 nsew signal input
flabel metal3 s 583520 16910 584800 17022 0 FreeSans 1120 0 0 0 io_in[3]
port 76 nsew signal input
flabel metal3 s 583520 21638 584800 21750 0 FreeSans 1120 0 0 0 io_in[4]
port 77 nsew signal input
flabel metal3 s 583520 48096 584800 48208 0 FreeSans 1120 0 0 0 io_in[5]
port 78 nsew signal input
flabel metal3 s 583520 92754 584800 92866 0 FreeSans 1120 0 0 0 io_in[6]
port 79 nsew signal input
flabel metal3 s 583520 272776 584800 272888 0 FreeSans 1120 0 0 0 io_in[7]
port 80 nsew signal input
flabel metal3 s 583520 317198 584800 317310 0 FreeSans 1120 0 0 0 io_in[8]
port 81 nsew signal input
flabel metal3 s 583520 362420 584800 362532 0 FreeSans 1120 0 0 0 io_in[9]
port 82 nsew signal input
flabel metal3 s 583520 1544 584800 1656 0 FreeSans 1120 0 0 0 io_in_3v3[0]
port 83 nsew signal input
flabel metal3 s 583520 407660 584800 407772 0 FreeSans 1120 0 0 0 io_in_3v3[10]
port 84 nsew signal input
flabel metal3 s 583520 452082 584800 452194 0 FreeSans 1120 0 0 0 io_in_3v3[11]
port 85 nsew signal input
flabel metal3 s 583520 496504 584800 496616 0 FreeSans 1120 0 0 0 io_in_3v3[12]
port 86 nsew signal input
flabel metal3 s 583520 585926 584800 586038 0 FreeSans 1120 0 0 0 io_in_3v3[13]
port 87 nsew signal input
flabel metal3 s -800 509166 480 509278 0 FreeSans 1120 0 0 0 io_in_3v3[14]
port 88 nsew signal input
flabel metal3 s -800 465944 480 466056 0 FreeSans 1120 0 0 0 io_in_3v3[15]
port 89 nsew signal input
flabel metal3 s -800 422722 480 422834 0 FreeSans 1120 0 0 0 io_in_3v3[16]
port 90 nsew signal input
flabel metal3 s -800 379500 480 379612 0 FreeSans 1120 0 0 0 io_in_3v3[17]
port 91 nsew signal input
flabel metal3 s -800 336278 480 336390 0 FreeSans 1120 0 0 0 io_in_3v3[18]
port 92 nsew signal input
flabel metal3 s -800 293056 480 293168 0 FreeSans 1120 0 0 0 io_in_3v3[19]
port 93 nsew signal input
flabel metal3 s 583520 6272 584800 6384 0 FreeSans 1120 0 0 0 io_in_3v3[1]
port 94 nsew signal input
flabel metal3 s -800 250034 480 250146 0 FreeSans 1120 0 0 0 io_in_3v3[20]
port 95 nsew signal input
flabel metal3 s -800 122412 480 122524 0 FreeSans 1120 0 0 0 io_in_3v3[21]
port 96 nsew signal input
flabel metal3 s -800 79190 480 79302 0 FreeSans 1120 0 0 0 io_in_3v3[22]
port 97 nsew signal input
flabel metal3 s -800 35968 480 36080 0 FreeSans 1120 0 0 0 io_in_3v3[23]
port 98 nsew signal input
flabel metal3 s -800 14546 480 14658 0 FreeSans 1120 0 0 0 io_in_3v3[24]
port 99 nsew signal input
flabel metal3 s -800 9818 480 9930 0 FreeSans 1120 0 0 0 io_in_3v3[25]
port 100 nsew signal input
flabel metal3 s -800 5090 480 5202 0 FreeSans 1120 0 0 0 io_in_3v3[26]
port 101 nsew signal input
flabel metal3 s 583520 11000 584800 11112 0 FreeSans 1120 0 0 0 io_in_3v3[2]
port 102 nsew signal input
flabel metal3 s 583520 15728 584800 15840 0 FreeSans 1120 0 0 0 io_in_3v3[3]
port 103 nsew signal input
flabel metal3 s 583520 20456 584800 20568 0 FreeSans 1120 0 0 0 io_in_3v3[4]
port 104 nsew signal input
flabel metal3 s 583520 46914 584800 47026 0 FreeSans 1120 0 0 0 io_in_3v3[5]
port 105 nsew signal input
flabel metal3 s 583520 91572 584800 91684 0 FreeSans 1120 0 0 0 io_in_3v3[6]
port 106 nsew signal input
flabel metal3 s 583520 271594 584800 271706 0 FreeSans 1120 0 0 0 io_in_3v3[7]
port 107 nsew signal input
flabel metal3 s 583520 316016 584800 316128 0 FreeSans 1120 0 0 0 io_in_3v3[8]
port 108 nsew signal input
flabel metal3 s 583520 361238 584800 361350 0 FreeSans 1120 0 0 0 io_in_3v3[9]
port 109 nsew signal input
flabel metal3 s 583520 5090 584800 5202 0 FreeSans 1120 0 0 0 io_oeb[0]
port 110 nsew signal tristate
flabel metal3 s 583520 411206 584800 411318 0 FreeSans 1120 0 0 0 io_oeb[10]
port 111 nsew signal tristate
flabel metal3 s 583520 455628 584800 455740 0 FreeSans 1120 0 0 0 io_oeb[11]
port 112 nsew signal tristate
flabel metal3 s 583520 500050 584800 500162 0 FreeSans 1120 0 0 0 io_oeb[12]
port 113 nsew signal tristate
flabel metal3 s 583520 589472 584800 589584 0 FreeSans 1120 0 0 0 io_oeb[13]
port 114 nsew signal tristate
flabel metal3 s -800 505620 480 505732 0 FreeSans 1120 0 0 0 io_oeb[14]
port 115 nsew signal tristate
flabel metal3 s -800 462398 480 462510 0 FreeSans 1120 0 0 0 io_oeb[15]
port 116 nsew signal tristate
flabel metal3 s -800 419176 480 419288 0 FreeSans 1120 0 0 0 io_oeb[16]
port 117 nsew signal tristate
flabel metal3 s -800 375954 480 376066 0 FreeSans 1120 0 0 0 io_oeb[17]
port 118 nsew signal tristate
flabel metal3 s -800 332732 480 332844 0 FreeSans 1120 0 0 0 io_oeb[18]
port 119 nsew signal tristate
flabel metal3 s -800 289510 480 289622 0 FreeSans 1120 0 0 0 io_oeb[19]
port 120 nsew signal tristate
flabel metal3 s 583520 9818 584800 9930 0 FreeSans 1120 0 0 0 io_oeb[1]
port 121 nsew signal tristate
flabel metal3 s -800 246488 480 246600 0 FreeSans 1120 0 0 0 io_oeb[20]
port 122 nsew signal tristate
flabel metal3 s -800 118866 480 118978 0 FreeSans 1120 0 0 0 io_oeb[21]
port 123 nsew signal tristate
flabel metal3 s -800 75644 480 75756 0 FreeSans 1120 0 0 0 io_oeb[22]
port 124 nsew signal tristate
flabel metal3 s -800 32422 480 32534 0 FreeSans 1120 0 0 0 io_oeb[23]
port 125 nsew signal tristate
flabel metal3 s -800 11000 480 11112 0 FreeSans 1120 0 0 0 io_oeb[24]
port 126 nsew signal tristate
flabel metal3 s -800 6272 480 6384 0 FreeSans 1120 0 0 0 io_oeb[25]
port 127 nsew signal tristate
flabel metal3 s -800 1544 480 1656 0 FreeSans 1120 0 0 0 io_oeb[26]
port 128 nsew signal tristate
flabel metal3 s 583520 14546 584800 14658 0 FreeSans 1120 0 0 0 io_oeb[2]
port 129 nsew signal tristate
flabel metal3 s 583520 19274 584800 19386 0 FreeSans 1120 0 0 0 io_oeb[3]
port 130 nsew signal tristate
flabel metal3 s 583520 24002 584800 24114 0 FreeSans 1120 0 0 0 io_oeb[4]
port 131 nsew signal tristate
flabel metal3 s 583520 50460 584800 50572 0 FreeSans 1120 0 0 0 io_oeb[5]
port 132 nsew signal tristate
flabel metal3 s 583520 95118 584800 95230 0 FreeSans 1120 0 0 0 io_oeb[6]
port 133 nsew signal tristate
flabel metal3 s 583520 275140 584800 275252 0 FreeSans 1120 0 0 0 io_oeb[7]
port 134 nsew signal tristate
flabel metal3 s 583520 319562 584800 319674 0 FreeSans 1120 0 0 0 io_oeb[8]
port 135 nsew signal tristate
flabel metal3 s 583520 364784 584800 364896 0 FreeSans 1120 0 0 0 io_oeb[9]
port 136 nsew signal tristate
flabel metal3 s 583520 3908 584800 4020 0 FreeSans 1120 0 0 0 io_out[0]
port 137 nsew signal tristate
flabel metal3 s 583520 410024 584800 410136 0 FreeSans 1120 0 0 0 io_out[10]
port 138 nsew signal tristate
flabel metal3 s 583520 454446 584800 454558 0 FreeSans 1120 0 0 0 io_out[11]
port 139 nsew signal tristate
flabel metal3 s 583520 498868 584800 498980 0 FreeSans 1120 0 0 0 io_out[12]
port 140 nsew signal tristate
flabel metal3 s 583520 588290 584800 588402 0 FreeSans 1120 0 0 0 io_out[13]
port 141 nsew signal tristate
flabel metal3 s -800 506802 480 506914 0 FreeSans 1120 0 0 0 io_out[14]
port 142 nsew signal tristate
flabel metal3 s -800 463580 480 463692 0 FreeSans 1120 0 0 0 io_out[15]
port 143 nsew signal tristate
flabel metal3 s -800 420358 480 420470 0 FreeSans 1120 0 0 0 io_out[16]
port 144 nsew signal tristate
flabel metal3 s -800 377136 480 377248 0 FreeSans 1120 0 0 0 io_out[17]
port 145 nsew signal tristate
flabel metal3 s -800 333914 480 334026 0 FreeSans 1120 0 0 0 io_out[18]
port 146 nsew signal tristate
flabel metal3 s -800 290692 480 290804 0 FreeSans 1120 0 0 0 io_out[19]
port 147 nsew signal tristate
flabel metal3 s 583520 8636 584800 8748 0 FreeSans 1120 0 0 0 io_out[1]
port 148 nsew signal tristate
flabel metal3 s -800 247670 480 247782 0 FreeSans 1120 0 0 0 io_out[20]
port 149 nsew signal tristate
flabel metal3 s -800 120048 480 120160 0 FreeSans 1120 0 0 0 io_out[21]
port 150 nsew signal tristate
flabel metal3 s -800 76826 480 76938 0 FreeSans 1120 0 0 0 io_out[22]
port 151 nsew signal tristate
flabel metal3 s -800 33604 480 33716 0 FreeSans 1120 0 0 0 io_out[23]
port 152 nsew signal tristate
flabel metal3 s -800 12182 480 12294 0 FreeSans 1120 0 0 0 io_out[24]
port 153 nsew signal tristate
flabel metal3 s -800 7454 480 7566 0 FreeSans 1120 0 0 0 io_out[25]
port 154 nsew signal tristate
flabel metal3 s -800 2726 480 2838 0 FreeSans 1120 0 0 0 io_out[26]
port 155 nsew signal tristate
flabel metal3 s 583520 13364 584800 13476 0 FreeSans 1120 0 0 0 io_out[2]
port 156 nsew signal tristate
flabel metal3 s 583520 18092 584800 18204 0 FreeSans 1120 0 0 0 io_out[3]
port 157 nsew signal tristate
flabel metal3 s 583520 22820 584800 22932 0 FreeSans 1120 0 0 0 io_out[4]
port 158 nsew signal tristate
flabel metal3 s 583520 49278 584800 49390 0 FreeSans 1120 0 0 0 io_out[5]
port 159 nsew signal tristate
flabel metal3 s 583520 93936 584800 94048 0 FreeSans 1120 0 0 0 io_out[6]
port 160 nsew signal tristate
flabel metal3 s 583520 273958 584800 274070 0 FreeSans 1120 0 0 0 io_out[7]
port 161 nsew signal tristate
flabel metal3 s 583520 318380 584800 318492 0 FreeSans 1120 0 0 0 io_out[8]
port 162 nsew signal tristate
flabel metal3 s 583520 363602 584800 363714 0 FreeSans 1120 0 0 0 io_out[9]
port 163 nsew signal tristate
flabel metal2 s 125816 -800 125928 480 0 FreeSans 1120 90 0 0 la_data_in[0]
port 164 nsew signal input
flabel metal2 s 480416 -800 480528 480 0 FreeSans 1120 90 0 0 la_data_in[100]
port 165 nsew signal input
flabel metal2 s 483962 -800 484074 480 0 FreeSans 1120 90 0 0 la_data_in[101]
port 166 nsew signal input
flabel metal2 s 487508 -800 487620 480 0 FreeSans 1120 90 0 0 la_data_in[102]
port 167 nsew signal input
flabel metal2 s 491054 -800 491166 480 0 FreeSans 1120 90 0 0 la_data_in[103]
port 168 nsew signal input
flabel metal2 s 494600 -800 494712 480 0 FreeSans 1120 90 0 0 la_data_in[104]
port 169 nsew signal input
flabel metal2 s 498146 -800 498258 480 0 FreeSans 1120 90 0 0 la_data_in[105]
port 170 nsew signal input
flabel metal2 s 501692 -800 501804 480 0 FreeSans 1120 90 0 0 la_data_in[106]
port 171 nsew signal input
flabel metal2 s 505238 -800 505350 480 0 FreeSans 1120 90 0 0 la_data_in[107]
port 172 nsew signal input
flabel metal2 s 508784 -800 508896 480 0 FreeSans 1120 90 0 0 la_data_in[108]
port 173 nsew signal input
flabel metal2 s 512330 -800 512442 480 0 FreeSans 1120 90 0 0 la_data_in[109]
port 174 nsew signal input
flabel metal2 s 161276 -800 161388 480 0 FreeSans 1120 90 0 0 la_data_in[10]
port 175 nsew signal input
flabel metal2 s 515876 -800 515988 480 0 FreeSans 1120 90 0 0 la_data_in[110]
port 176 nsew signal input
flabel metal2 s 519422 -800 519534 480 0 FreeSans 1120 90 0 0 la_data_in[111]
port 177 nsew signal input
flabel metal2 s 522968 -800 523080 480 0 FreeSans 1120 90 0 0 la_data_in[112]
port 178 nsew signal input
flabel metal2 s 526514 -800 526626 480 0 FreeSans 1120 90 0 0 la_data_in[113]
port 179 nsew signal input
flabel metal2 s 530060 -800 530172 480 0 FreeSans 1120 90 0 0 la_data_in[114]
port 180 nsew signal input
flabel metal2 s 533606 -800 533718 480 0 FreeSans 1120 90 0 0 la_data_in[115]
port 181 nsew signal input
flabel metal2 s 537152 -800 537264 480 0 FreeSans 1120 90 0 0 la_data_in[116]
port 182 nsew signal input
flabel metal2 s 540698 -800 540810 480 0 FreeSans 1120 90 0 0 la_data_in[117]
port 183 nsew signal input
flabel metal2 s 544244 -800 544356 480 0 FreeSans 1120 90 0 0 la_data_in[118]
port 184 nsew signal input
flabel metal2 s 547790 -800 547902 480 0 FreeSans 1120 90 0 0 la_data_in[119]
port 185 nsew signal input
flabel metal2 s 164822 -800 164934 480 0 FreeSans 1120 90 0 0 la_data_in[11]
port 186 nsew signal input
flabel metal2 s 551336 -800 551448 480 0 FreeSans 1120 90 0 0 la_data_in[120]
port 187 nsew signal input
flabel metal2 s 554882 -800 554994 480 0 FreeSans 1120 90 0 0 la_data_in[121]
port 188 nsew signal input
flabel metal2 s 558428 -800 558540 480 0 FreeSans 1120 90 0 0 la_data_in[122]
port 189 nsew signal input
flabel metal2 s 561974 -800 562086 480 0 FreeSans 1120 90 0 0 la_data_in[123]
port 190 nsew signal input
flabel metal2 s 565520 -800 565632 480 0 FreeSans 1120 90 0 0 la_data_in[124]
port 191 nsew signal input
flabel metal2 s 569066 -800 569178 480 0 FreeSans 1120 90 0 0 la_data_in[125]
port 192 nsew signal input
flabel metal2 s 572612 -800 572724 480 0 FreeSans 1120 90 0 0 la_data_in[126]
port 193 nsew signal input
flabel metal2 s 576158 -800 576270 480 0 FreeSans 1120 90 0 0 la_data_in[127]
port 194 nsew signal input
flabel metal2 s 168368 -800 168480 480 0 FreeSans 1120 90 0 0 la_data_in[12]
port 195 nsew signal input
flabel metal2 s 171914 -800 172026 480 0 FreeSans 1120 90 0 0 la_data_in[13]
port 196 nsew signal input
flabel metal2 s 175460 -800 175572 480 0 FreeSans 1120 90 0 0 la_data_in[14]
port 197 nsew signal input
flabel metal2 s 179006 -800 179118 480 0 FreeSans 1120 90 0 0 la_data_in[15]
port 198 nsew signal input
flabel metal2 s 182552 -800 182664 480 0 FreeSans 1120 90 0 0 la_data_in[16]
port 199 nsew signal input
flabel metal2 s 186098 -800 186210 480 0 FreeSans 1120 90 0 0 la_data_in[17]
port 200 nsew signal input
flabel metal2 s 189644 -800 189756 480 0 FreeSans 1120 90 0 0 la_data_in[18]
port 201 nsew signal input
flabel metal2 s 193190 -800 193302 480 0 FreeSans 1120 90 0 0 la_data_in[19]
port 202 nsew signal input
flabel metal2 s 129362 -800 129474 480 0 FreeSans 1120 90 0 0 la_data_in[1]
port 203 nsew signal input
flabel metal2 s 196736 -800 196848 480 0 FreeSans 1120 90 0 0 la_data_in[20]
port 204 nsew signal input
flabel metal2 s 200282 -800 200394 480 0 FreeSans 1120 90 0 0 la_data_in[21]
port 205 nsew signal input
flabel metal2 s 203828 -800 203940 480 0 FreeSans 1120 90 0 0 la_data_in[22]
port 206 nsew signal input
flabel metal2 s 207374 -800 207486 480 0 FreeSans 1120 90 0 0 la_data_in[23]
port 207 nsew signal input
flabel metal2 s 210920 -800 211032 480 0 FreeSans 1120 90 0 0 la_data_in[24]
port 208 nsew signal input
flabel metal2 s 214466 -800 214578 480 0 FreeSans 1120 90 0 0 la_data_in[25]
port 209 nsew signal input
flabel metal2 s 218012 -800 218124 480 0 FreeSans 1120 90 0 0 la_data_in[26]
port 210 nsew signal input
flabel metal2 s 221558 -800 221670 480 0 FreeSans 1120 90 0 0 la_data_in[27]
port 211 nsew signal input
flabel metal2 s 225104 -800 225216 480 0 FreeSans 1120 90 0 0 la_data_in[28]
port 212 nsew signal input
flabel metal2 s 228650 -800 228762 480 0 FreeSans 1120 90 0 0 la_data_in[29]
port 213 nsew signal input
flabel metal2 s 132908 -800 133020 480 0 FreeSans 1120 90 0 0 la_data_in[2]
port 214 nsew signal input
flabel metal2 s 232196 -800 232308 480 0 FreeSans 1120 90 0 0 la_data_in[30]
port 215 nsew signal input
flabel metal2 s 235742 -800 235854 480 0 FreeSans 1120 90 0 0 la_data_in[31]
port 216 nsew signal input
flabel metal2 s 239288 -800 239400 480 0 FreeSans 1120 90 0 0 la_data_in[32]
port 217 nsew signal input
flabel metal2 s 242834 -800 242946 480 0 FreeSans 1120 90 0 0 la_data_in[33]
port 218 nsew signal input
flabel metal2 s 246380 -800 246492 480 0 FreeSans 1120 90 0 0 la_data_in[34]
port 219 nsew signal input
flabel metal2 s 249926 -800 250038 480 0 FreeSans 1120 90 0 0 la_data_in[35]
port 220 nsew signal input
flabel metal2 s 253472 -800 253584 480 0 FreeSans 1120 90 0 0 la_data_in[36]
port 221 nsew signal input
flabel metal2 s 257018 -800 257130 480 0 FreeSans 1120 90 0 0 la_data_in[37]
port 222 nsew signal input
flabel metal2 s 260564 -800 260676 480 0 FreeSans 1120 90 0 0 la_data_in[38]
port 223 nsew signal input
flabel metal2 s 264110 -800 264222 480 0 FreeSans 1120 90 0 0 la_data_in[39]
port 224 nsew signal input
flabel metal2 s 136454 -800 136566 480 0 FreeSans 1120 90 0 0 la_data_in[3]
port 225 nsew signal input
flabel metal2 s 267656 -800 267768 480 0 FreeSans 1120 90 0 0 la_data_in[40]
port 226 nsew signal input
flabel metal2 s 271202 -800 271314 480 0 FreeSans 1120 90 0 0 la_data_in[41]
port 227 nsew signal input
flabel metal2 s 274748 -800 274860 480 0 FreeSans 1120 90 0 0 la_data_in[42]
port 228 nsew signal input
flabel metal2 s 278294 -800 278406 480 0 FreeSans 1120 90 0 0 la_data_in[43]
port 229 nsew signal input
flabel metal2 s 281840 -800 281952 480 0 FreeSans 1120 90 0 0 la_data_in[44]
port 230 nsew signal input
flabel metal2 s 285386 -800 285498 480 0 FreeSans 1120 90 0 0 la_data_in[45]
port 231 nsew signal input
flabel metal2 s 288932 -800 289044 480 0 FreeSans 1120 90 0 0 la_data_in[46]
port 232 nsew signal input
flabel metal2 s 292478 -800 292590 480 0 FreeSans 1120 90 0 0 la_data_in[47]
port 233 nsew signal input
flabel metal2 s 296024 -800 296136 480 0 FreeSans 1120 90 0 0 la_data_in[48]
port 234 nsew signal input
flabel metal2 s 299570 -800 299682 480 0 FreeSans 1120 90 0 0 la_data_in[49]
port 235 nsew signal input
flabel metal2 s 140000 -800 140112 480 0 FreeSans 1120 90 0 0 la_data_in[4]
port 236 nsew signal input
flabel metal2 s 303116 -800 303228 480 0 FreeSans 1120 90 0 0 la_data_in[50]
port 237 nsew signal input
flabel metal2 s 306662 -800 306774 480 0 FreeSans 1120 90 0 0 la_data_in[51]
port 238 nsew signal input
flabel metal2 s 310208 -800 310320 480 0 FreeSans 1120 90 0 0 la_data_in[52]
port 239 nsew signal input
flabel metal2 s 313754 -800 313866 480 0 FreeSans 1120 90 0 0 la_data_in[53]
port 240 nsew signal input
flabel metal2 s 317300 -800 317412 480 0 FreeSans 1120 90 0 0 la_data_in[54]
port 241 nsew signal input
flabel metal2 s 320846 -800 320958 480 0 FreeSans 1120 90 0 0 la_data_in[55]
port 242 nsew signal input
flabel metal2 s 324392 -800 324504 480 0 FreeSans 1120 90 0 0 la_data_in[56]
port 243 nsew signal input
flabel metal2 s 327938 -800 328050 480 0 FreeSans 1120 90 0 0 la_data_in[57]
port 244 nsew signal input
flabel metal2 s 331484 -800 331596 480 0 FreeSans 1120 90 0 0 la_data_in[58]
port 245 nsew signal input
flabel metal2 s 335030 -800 335142 480 0 FreeSans 1120 90 0 0 la_data_in[59]
port 246 nsew signal input
flabel metal2 s 143546 -800 143658 480 0 FreeSans 1120 90 0 0 la_data_in[5]
port 247 nsew signal input
flabel metal2 s 338576 -800 338688 480 0 FreeSans 1120 90 0 0 la_data_in[60]
port 248 nsew signal input
flabel metal2 s 342122 -800 342234 480 0 FreeSans 1120 90 0 0 la_data_in[61]
port 249 nsew signal input
flabel metal2 s 345668 -800 345780 480 0 FreeSans 1120 90 0 0 la_data_in[62]
port 250 nsew signal input
flabel metal2 s 349214 -800 349326 480 0 FreeSans 1120 90 0 0 la_data_in[63]
port 251 nsew signal input
flabel metal2 s 352760 -800 352872 480 0 FreeSans 1120 90 0 0 la_data_in[64]
port 252 nsew signal input
flabel metal2 s 356306 -800 356418 480 0 FreeSans 1120 90 0 0 la_data_in[65]
port 253 nsew signal input
flabel metal2 s 359852 -800 359964 480 0 FreeSans 1120 90 0 0 la_data_in[66]
port 254 nsew signal input
flabel metal2 s 363398 -800 363510 480 0 FreeSans 1120 90 0 0 la_data_in[67]
port 255 nsew signal input
flabel metal2 s 366944 -800 367056 480 0 FreeSans 1120 90 0 0 la_data_in[68]
port 256 nsew signal input
flabel metal2 s 370490 -800 370602 480 0 FreeSans 1120 90 0 0 la_data_in[69]
port 257 nsew signal input
flabel metal2 s 147092 -800 147204 480 0 FreeSans 1120 90 0 0 la_data_in[6]
port 258 nsew signal input
flabel metal2 s 374036 -800 374148 480 0 FreeSans 1120 90 0 0 la_data_in[70]
port 259 nsew signal input
flabel metal2 s 377582 -800 377694 480 0 FreeSans 1120 90 0 0 la_data_in[71]
port 260 nsew signal input
flabel metal2 s 381128 -800 381240 480 0 FreeSans 1120 90 0 0 la_data_in[72]
port 261 nsew signal input
flabel metal2 s 384674 -800 384786 480 0 FreeSans 1120 90 0 0 la_data_in[73]
port 262 nsew signal input
flabel metal2 s 388220 -800 388332 480 0 FreeSans 1120 90 0 0 la_data_in[74]
port 263 nsew signal input
flabel metal2 s 391766 -800 391878 480 0 FreeSans 1120 90 0 0 la_data_in[75]
port 264 nsew signal input
flabel metal2 s 395312 -800 395424 480 0 FreeSans 1120 90 0 0 la_data_in[76]
port 265 nsew signal input
flabel metal2 s 398858 -800 398970 480 0 FreeSans 1120 90 0 0 la_data_in[77]
port 266 nsew signal input
flabel metal2 s 402404 -800 402516 480 0 FreeSans 1120 90 0 0 la_data_in[78]
port 267 nsew signal input
flabel metal2 s 405950 -800 406062 480 0 FreeSans 1120 90 0 0 la_data_in[79]
port 268 nsew signal input
flabel metal2 s 150638 -800 150750 480 0 FreeSans 1120 90 0 0 la_data_in[7]
port 269 nsew signal input
flabel metal2 s 409496 -800 409608 480 0 FreeSans 1120 90 0 0 la_data_in[80]
port 270 nsew signal input
flabel metal2 s 413042 -800 413154 480 0 FreeSans 1120 90 0 0 la_data_in[81]
port 271 nsew signal input
flabel metal2 s 416588 -800 416700 480 0 FreeSans 1120 90 0 0 la_data_in[82]
port 272 nsew signal input
flabel metal2 s 420134 -800 420246 480 0 FreeSans 1120 90 0 0 la_data_in[83]
port 273 nsew signal input
flabel metal2 s 423680 -800 423792 480 0 FreeSans 1120 90 0 0 la_data_in[84]
port 274 nsew signal input
flabel metal2 s 427226 -800 427338 480 0 FreeSans 1120 90 0 0 la_data_in[85]
port 275 nsew signal input
flabel metal2 s 430772 -800 430884 480 0 FreeSans 1120 90 0 0 la_data_in[86]
port 276 nsew signal input
flabel metal2 s 434318 -800 434430 480 0 FreeSans 1120 90 0 0 la_data_in[87]
port 277 nsew signal input
flabel metal2 s 437864 -800 437976 480 0 FreeSans 1120 90 0 0 la_data_in[88]
port 278 nsew signal input
flabel metal2 s 441410 -800 441522 480 0 FreeSans 1120 90 0 0 la_data_in[89]
port 279 nsew signal input
flabel metal2 s 154184 -800 154296 480 0 FreeSans 1120 90 0 0 la_data_in[8]
port 280 nsew signal input
flabel metal2 s 444956 -800 445068 480 0 FreeSans 1120 90 0 0 la_data_in[90]
port 281 nsew signal input
flabel metal2 s 448502 -800 448614 480 0 FreeSans 1120 90 0 0 la_data_in[91]
port 282 nsew signal input
flabel metal2 s 452048 -800 452160 480 0 FreeSans 1120 90 0 0 la_data_in[92]
port 283 nsew signal input
flabel metal2 s 455594 -800 455706 480 0 FreeSans 1120 90 0 0 la_data_in[93]
port 284 nsew signal input
flabel metal2 s 459140 -800 459252 480 0 FreeSans 1120 90 0 0 la_data_in[94]
port 285 nsew signal input
flabel metal2 s 462686 -800 462798 480 0 FreeSans 1120 90 0 0 la_data_in[95]
port 286 nsew signal input
flabel metal2 s 466232 -800 466344 480 0 FreeSans 1120 90 0 0 la_data_in[96]
port 287 nsew signal input
flabel metal2 s 469778 -800 469890 480 0 FreeSans 1120 90 0 0 la_data_in[97]
port 288 nsew signal input
flabel metal2 s 473324 -800 473436 480 0 FreeSans 1120 90 0 0 la_data_in[98]
port 289 nsew signal input
flabel metal2 s 476870 -800 476982 480 0 FreeSans 1120 90 0 0 la_data_in[99]
port 290 nsew signal input
flabel metal2 s 157730 -800 157842 480 0 FreeSans 1120 90 0 0 la_data_in[9]
port 291 nsew signal input
flabel metal2 s 126998 -800 127110 480 0 FreeSans 1120 90 0 0 la_data_out[0]
port 292 nsew signal tristate
flabel metal2 s 481598 -800 481710 480 0 FreeSans 1120 90 0 0 la_data_out[100]
port 293 nsew signal tristate
flabel metal2 s 485144 -800 485256 480 0 FreeSans 1120 90 0 0 la_data_out[101]
port 294 nsew signal tristate
flabel metal2 s 488690 -800 488802 480 0 FreeSans 1120 90 0 0 la_data_out[102]
port 295 nsew signal tristate
flabel metal2 s 492236 -800 492348 480 0 FreeSans 1120 90 0 0 la_data_out[103]
port 296 nsew signal tristate
flabel metal2 s 495782 -800 495894 480 0 FreeSans 1120 90 0 0 la_data_out[104]
port 297 nsew signal tristate
flabel metal2 s 499328 -800 499440 480 0 FreeSans 1120 90 0 0 la_data_out[105]
port 298 nsew signal tristate
flabel metal2 s 502874 -800 502986 480 0 FreeSans 1120 90 0 0 la_data_out[106]
port 299 nsew signal tristate
flabel metal2 s 506420 -800 506532 480 0 FreeSans 1120 90 0 0 la_data_out[107]
port 300 nsew signal tristate
flabel metal2 s 509966 -800 510078 480 0 FreeSans 1120 90 0 0 la_data_out[108]
port 301 nsew signal tristate
flabel metal2 s 513512 -800 513624 480 0 FreeSans 1120 90 0 0 la_data_out[109]
port 302 nsew signal tristate
flabel metal2 s 162458 -800 162570 480 0 FreeSans 1120 90 0 0 la_data_out[10]
port 303 nsew signal tristate
flabel metal2 s 517058 -800 517170 480 0 FreeSans 1120 90 0 0 la_data_out[110]
port 304 nsew signal tristate
flabel metal2 s 520604 -800 520716 480 0 FreeSans 1120 90 0 0 la_data_out[111]
port 305 nsew signal tristate
flabel metal2 s 524150 -800 524262 480 0 FreeSans 1120 90 0 0 la_data_out[112]
port 306 nsew signal tristate
flabel metal2 s 527696 -800 527808 480 0 FreeSans 1120 90 0 0 la_data_out[113]
port 307 nsew signal tristate
flabel metal2 s 531242 -800 531354 480 0 FreeSans 1120 90 0 0 la_data_out[114]
port 308 nsew signal tristate
flabel metal2 s 534788 -800 534900 480 0 FreeSans 1120 90 0 0 la_data_out[115]
port 309 nsew signal tristate
flabel metal2 s 538334 -800 538446 480 0 FreeSans 1120 90 0 0 la_data_out[116]
port 310 nsew signal tristate
flabel metal2 s 541880 -800 541992 480 0 FreeSans 1120 90 0 0 la_data_out[117]
port 311 nsew signal tristate
flabel metal2 s 545426 -800 545538 480 0 FreeSans 1120 90 0 0 la_data_out[118]
port 312 nsew signal tristate
flabel metal2 s 548972 -800 549084 480 0 FreeSans 1120 90 0 0 la_data_out[119]
port 313 nsew signal tristate
flabel metal2 s 166004 -800 166116 480 0 FreeSans 1120 90 0 0 la_data_out[11]
port 314 nsew signal tristate
flabel metal2 s 552518 -800 552630 480 0 FreeSans 1120 90 0 0 la_data_out[120]
port 315 nsew signal tristate
flabel metal2 s 556064 -800 556176 480 0 FreeSans 1120 90 0 0 la_data_out[121]
port 316 nsew signal tristate
flabel metal2 s 559610 -800 559722 480 0 FreeSans 1120 90 0 0 la_data_out[122]
port 317 nsew signal tristate
flabel metal2 s 563156 -800 563268 480 0 FreeSans 1120 90 0 0 la_data_out[123]
port 318 nsew signal tristate
flabel metal2 s 566702 -800 566814 480 0 FreeSans 1120 90 0 0 la_data_out[124]
port 319 nsew signal tristate
flabel metal2 s 570248 -800 570360 480 0 FreeSans 1120 90 0 0 la_data_out[125]
port 320 nsew signal tristate
flabel metal2 s 573794 -800 573906 480 0 FreeSans 1120 90 0 0 la_data_out[126]
port 321 nsew signal tristate
flabel metal2 s 577340 -800 577452 480 0 FreeSans 1120 90 0 0 la_data_out[127]
port 322 nsew signal tristate
flabel metal2 s 169550 -800 169662 480 0 FreeSans 1120 90 0 0 la_data_out[12]
port 323 nsew signal tristate
flabel metal2 s 173096 -800 173208 480 0 FreeSans 1120 90 0 0 la_data_out[13]
port 324 nsew signal tristate
flabel metal2 s 176642 -800 176754 480 0 FreeSans 1120 90 0 0 la_data_out[14]
port 325 nsew signal tristate
flabel metal2 s 180188 -800 180300 480 0 FreeSans 1120 90 0 0 la_data_out[15]
port 326 nsew signal tristate
flabel metal2 s 183734 -800 183846 480 0 FreeSans 1120 90 0 0 la_data_out[16]
port 327 nsew signal tristate
flabel metal2 s 187280 -800 187392 480 0 FreeSans 1120 90 0 0 la_data_out[17]
port 328 nsew signal tristate
flabel metal2 s 190826 -800 190938 480 0 FreeSans 1120 90 0 0 la_data_out[18]
port 329 nsew signal tristate
flabel metal2 s 194372 -800 194484 480 0 FreeSans 1120 90 0 0 la_data_out[19]
port 330 nsew signal tristate
flabel metal2 s 130544 -800 130656 480 0 FreeSans 1120 90 0 0 la_data_out[1]
port 331 nsew signal tristate
flabel metal2 s 197918 -800 198030 480 0 FreeSans 1120 90 0 0 la_data_out[20]
port 332 nsew signal tristate
flabel metal2 s 201464 -800 201576 480 0 FreeSans 1120 90 0 0 la_data_out[21]
port 333 nsew signal tristate
flabel metal2 s 205010 -800 205122 480 0 FreeSans 1120 90 0 0 la_data_out[22]
port 334 nsew signal tristate
flabel metal2 s 208556 -800 208668 480 0 FreeSans 1120 90 0 0 la_data_out[23]
port 335 nsew signal tristate
flabel metal2 s 212102 -800 212214 480 0 FreeSans 1120 90 0 0 la_data_out[24]
port 336 nsew signal tristate
flabel metal2 s 215648 -800 215760 480 0 FreeSans 1120 90 0 0 la_data_out[25]
port 337 nsew signal tristate
flabel metal2 s 219194 -800 219306 480 0 FreeSans 1120 90 0 0 la_data_out[26]
port 338 nsew signal tristate
flabel metal2 s 222740 -800 222852 480 0 FreeSans 1120 90 0 0 la_data_out[27]
port 339 nsew signal tristate
flabel metal2 s 226286 -800 226398 480 0 FreeSans 1120 90 0 0 la_data_out[28]
port 340 nsew signal tristate
flabel metal2 s 229832 -800 229944 480 0 FreeSans 1120 90 0 0 la_data_out[29]
port 341 nsew signal tristate
flabel metal2 s 134090 -800 134202 480 0 FreeSans 1120 90 0 0 la_data_out[2]
port 342 nsew signal tristate
flabel metal2 s 233378 -800 233490 480 0 FreeSans 1120 90 0 0 la_data_out[30]
port 343 nsew signal tristate
flabel metal2 s 236924 -800 237036 480 0 FreeSans 1120 90 0 0 la_data_out[31]
port 344 nsew signal tristate
flabel metal2 s 240470 -800 240582 480 0 FreeSans 1120 90 0 0 la_data_out[32]
port 345 nsew signal tristate
flabel metal2 s 244016 -800 244128 480 0 FreeSans 1120 90 0 0 la_data_out[33]
port 346 nsew signal tristate
flabel metal2 s 247562 -800 247674 480 0 FreeSans 1120 90 0 0 la_data_out[34]
port 347 nsew signal tristate
flabel metal2 s 251108 -800 251220 480 0 FreeSans 1120 90 0 0 la_data_out[35]
port 348 nsew signal tristate
flabel metal2 s 254654 -800 254766 480 0 FreeSans 1120 90 0 0 la_data_out[36]
port 349 nsew signal tristate
flabel metal2 s 258200 -800 258312 480 0 FreeSans 1120 90 0 0 la_data_out[37]
port 350 nsew signal tristate
flabel metal2 s 261746 -800 261858 480 0 FreeSans 1120 90 0 0 la_data_out[38]
port 351 nsew signal tristate
flabel metal2 s 265292 -800 265404 480 0 FreeSans 1120 90 0 0 la_data_out[39]
port 352 nsew signal tristate
flabel metal2 s 137636 -800 137748 480 0 FreeSans 1120 90 0 0 la_data_out[3]
port 353 nsew signal tristate
flabel metal2 s 268838 -800 268950 480 0 FreeSans 1120 90 0 0 la_data_out[40]
port 354 nsew signal tristate
flabel metal2 s 272384 -800 272496 480 0 FreeSans 1120 90 0 0 la_data_out[41]
port 355 nsew signal tristate
flabel metal2 s 275930 -800 276042 480 0 FreeSans 1120 90 0 0 la_data_out[42]
port 356 nsew signal tristate
flabel metal2 s 279476 -800 279588 480 0 FreeSans 1120 90 0 0 la_data_out[43]
port 357 nsew signal tristate
flabel metal2 s 283022 -800 283134 480 0 FreeSans 1120 90 0 0 la_data_out[44]
port 358 nsew signal tristate
flabel metal2 s 286568 -800 286680 480 0 FreeSans 1120 90 0 0 la_data_out[45]
port 359 nsew signal tristate
flabel metal2 s 290114 -800 290226 480 0 FreeSans 1120 90 0 0 la_data_out[46]
port 360 nsew signal tristate
flabel metal2 s 293660 -800 293772 480 0 FreeSans 1120 90 0 0 la_data_out[47]
port 361 nsew signal tristate
flabel metal2 s 297206 -800 297318 480 0 FreeSans 1120 90 0 0 la_data_out[48]
port 362 nsew signal tristate
flabel metal2 s 300752 -800 300864 480 0 FreeSans 1120 90 0 0 la_data_out[49]
port 363 nsew signal tristate
flabel metal2 s 141182 -800 141294 480 0 FreeSans 1120 90 0 0 la_data_out[4]
port 364 nsew signal tristate
flabel metal2 s 304298 -800 304410 480 0 FreeSans 1120 90 0 0 la_data_out[50]
port 365 nsew signal tristate
flabel metal2 s 307844 -800 307956 480 0 FreeSans 1120 90 0 0 la_data_out[51]
port 366 nsew signal tristate
flabel metal2 s 311390 -800 311502 480 0 FreeSans 1120 90 0 0 la_data_out[52]
port 367 nsew signal tristate
flabel metal2 s 314936 -800 315048 480 0 FreeSans 1120 90 0 0 la_data_out[53]
port 368 nsew signal tristate
flabel metal2 s 318482 -800 318594 480 0 FreeSans 1120 90 0 0 la_data_out[54]
port 369 nsew signal tristate
flabel metal2 s 322028 -800 322140 480 0 FreeSans 1120 90 0 0 la_data_out[55]
port 370 nsew signal tristate
flabel metal2 s 325574 -800 325686 480 0 FreeSans 1120 90 0 0 la_data_out[56]
port 371 nsew signal tristate
flabel metal2 s 329120 -800 329232 480 0 FreeSans 1120 90 0 0 la_data_out[57]
port 372 nsew signal tristate
flabel metal2 s 332666 -800 332778 480 0 FreeSans 1120 90 0 0 la_data_out[58]
port 373 nsew signal tristate
flabel metal2 s 336212 -800 336324 480 0 FreeSans 1120 90 0 0 la_data_out[59]
port 374 nsew signal tristate
flabel metal2 s 144728 -800 144840 480 0 FreeSans 1120 90 0 0 la_data_out[5]
port 375 nsew signal tristate
flabel metal2 s 339758 -800 339870 480 0 FreeSans 1120 90 0 0 la_data_out[60]
port 376 nsew signal tristate
flabel metal2 s 343304 -800 343416 480 0 FreeSans 1120 90 0 0 la_data_out[61]
port 377 nsew signal tristate
flabel metal2 s 346850 -800 346962 480 0 FreeSans 1120 90 0 0 la_data_out[62]
port 378 nsew signal tristate
flabel metal2 s 350396 -800 350508 480 0 FreeSans 1120 90 0 0 la_data_out[63]
port 379 nsew signal tristate
flabel metal2 s 353942 -800 354054 480 0 FreeSans 1120 90 0 0 la_data_out[64]
port 380 nsew signal tristate
flabel metal2 s 357488 -800 357600 480 0 FreeSans 1120 90 0 0 la_data_out[65]
port 381 nsew signal tristate
flabel metal2 s 361034 -800 361146 480 0 FreeSans 1120 90 0 0 la_data_out[66]
port 382 nsew signal tristate
flabel metal2 s 364580 -800 364692 480 0 FreeSans 1120 90 0 0 la_data_out[67]
port 383 nsew signal tristate
flabel metal2 s 368126 -800 368238 480 0 FreeSans 1120 90 0 0 la_data_out[68]
port 384 nsew signal tristate
flabel metal2 s 371672 -800 371784 480 0 FreeSans 1120 90 0 0 la_data_out[69]
port 385 nsew signal tristate
flabel metal2 s 148274 -800 148386 480 0 FreeSans 1120 90 0 0 la_data_out[6]
port 386 nsew signal tristate
flabel metal2 s 375218 -800 375330 480 0 FreeSans 1120 90 0 0 la_data_out[70]
port 387 nsew signal tristate
flabel metal2 s 378764 -800 378876 480 0 FreeSans 1120 90 0 0 la_data_out[71]
port 388 nsew signal tristate
flabel metal2 s 382310 -800 382422 480 0 FreeSans 1120 90 0 0 la_data_out[72]
port 389 nsew signal tristate
flabel metal2 s 385856 -800 385968 480 0 FreeSans 1120 90 0 0 la_data_out[73]
port 390 nsew signal tristate
flabel metal2 s 389402 -800 389514 480 0 FreeSans 1120 90 0 0 la_data_out[74]
port 391 nsew signal tristate
flabel metal2 s 392948 -800 393060 480 0 FreeSans 1120 90 0 0 la_data_out[75]
port 392 nsew signal tristate
flabel metal2 s 396494 -800 396606 480 0 FreeSans 1120 90 0 0 la_data_out[76]
port 393 nsew signal tristate
flabel metal2 s 400040 -800 400152 480 0 FreeSans 1120 90 0 0 la_data_out[77]
port 394 nsew signal tristate
flabel metal2 s 403586 -800 403698 480 0 FreeSans 1120 90 0 0 la_data_out[78]
port 395 nsew signal tristate
flabel metal2 s 407132 -800 407244 480 0 FreeSans 1120 90 0 0 la_data_out[79]
port 396 nsew signal tristate
flabel metal2 s 151820 -800 151932 480 0 FreeSans 1120 90 0 0 la_data_out[7]
port 397 nsew signal tristate
flabel metal2 s 410678 -800 410790 480 0 FreeSans 1120 90 0 0 la_data_out[80]
port 398 nsew signal tristate
flabel metal2 s 414224 -800 414336 480 0 FreeSans 1120 90 0 0 la_data_out[81]
port 399 nsew signal tristate
flabel metal2 s 417770 -800 417882 480 0 FreeSans 1120 90 0 0 la_data_out[82]
port 400 nsew signal tristate
flabel metal2 s 421316 -800 421428 480 0 FreeSans 1120 90 0 0 la_data_out[83]
port 401 nsew signal tristate
flabel metal2 s 424862 -800 424974 480 0 FreeSans 1120 90 0 0 la_data_out[84]
port 402 nsew signal tristate
flabel metal2 s 428408 -800 428520 480 0 FreeSans 1120 90 0 0 la_data_out[85]
port 403 nsew signal tristate
flabel metal2 s 431954 -800 432066 480 0 FreeSans 1120 90 0 0 la_data_out[86]
port 404 nsew signal tristate
flabel metal2 s 435500 -800 435612 480 0 FreeSans 1120 90 0 0 la_data_out[87]
port 405 nsew signal tristate
flabel metal2 s 439046 -800 439158 480 0 FreeSans 1120 90 0 0 la_data_out[88]
port 406 nsew signal tristate
flabel metal2 s 442592 -800 442704 480 0 FreeSans 1120 90 0 0 la_data_out[89]
port 407 nsew signal tristate
flabel metal2 s 155366 -800 155478 480 0 FreeSans 1120 90 0 0 la_data_out[8]
port 408 nsew signal tristate
flabel metal2 s 446138 -800 446250 480 0 FreeSans 1120 90 0 0 la_data_out[90]
port 409 nsew signal tristate
flabel metal2 s 449684 -800 449796 480 0 FreeSans 1120 90 0 0 la_data_out[91]
port 410 nsew signal tristate
flabel metal2 s 453230 -800 453342 480 0 FreeSans 1120 90 0 0 la_data_out[92]
port 411 nsew signal tristate
flabel metal2 s 456776 -800 456888 480 0 FreeSans 1120 90 0 0 la_data_out[93]
port 412 nsew signal tristate
flabel metal2 s 460322 -800 460434 480 0 FreeSans 1120 90 0 0 la_data_out[94]
port 413 nsew signal tristate
flabel metal2 s 463868 -800 463980 480 0 FreeSans 1120 90 0 0 la_data_out[95]
port 414 nsew signal tristate
flabel metal2 s 467414 -800 467526 480 0 FreeSans 1120 90 0 0 la_data_out[96]
port 415 nsew signal tristate
flabel metal2 s 470960 -800 471072 480 0 FreeSans 1120 90 0 0 la_data_out[97]
port 416 nsew signal tristate
flabel metal2 s 474506 -800 474618 480 0 FreeSans 1120 90 0 0 la_data_out[98]
port 417 nsew signal tristate
flabel metal2 s 478052 -800 478164 480 0 FreeSans 1120 90 0 0 la_data_out[99]
port 418 nsew signal tristate
flabel metal2 s 158912 -800 159024 480 0 FreeSans 1120 90 0 0 la_data_out[9]
port 419 nsew signal tristate
flabel metal2 s 128180 -800 128292 480 0 FreeSans 1120 90 0 0 la_oenb[0]
port 420 nsew signal input
flabel metal2 s 482780 -800 482892 480 0 FreeSans 1120 90 0 0 la_oenb[100]
port 421 nsew signal input
flabel metal2 s 486326 -800 486438 480 0 FreeSans 1120 90 0 0 la_oenb[101]
port 422 nsew signal input
flabel metal2 s 489872 -800 489984 480 0 FreeSans 1120 90 0 0 la_oenb[102]
port 423 nsew signal input
flabel metal2 s 493418 -800 493530 480 0 FreeSans 1120 90 0 0 la_oenb[103]
port 424 nsew signal input
flabel metal2 s 496964 -800 497076 480 0 FreeSans 1120 90 0 0 la_oenb[104]
port 425 nsew signal input
flabel metal2 s 500510 -800 500622 480 0 FreeSans 1120 90 0 0 la_oenb[105]
port 426 nsew signal input
flabel metal2 s 504056 -800 504168 480 0 FreeSans 1120 90 0 0 la_oenb[106]
port 427 nsew signal input
flabel metal2 s 507602 -800 507714 480 0 FreeSans 1120 90 0 0 la_oenb[107]
port 428 nsew signal input
flabel metal2 s 511148 -800 511260 480 0 FreeSans 1120 90 0 0 la_oenb[108]
port 429 nsew signal input
flabel metal2 s 514694 -800 514806 480 0 FreeSans 1120 90 0 0 la_oenb[109]
port 430 nsew signal input
flabel metal2 s 163640 -800 163752 480 0 FreeSans 1120 90 0 0 la_oenb[10]
port 431 nsew signal input
flabel metal2 s 518240 -800 518352 480 0 FreeSans 1120 90 0 0 la_oenb[110]
port 432 nsew signal input
flabel metal2 s 521786 -800 521898 480 0 FreeSans 1120 90 0 0 la_oenb[111]
port 433 nsew signal input
flabel metal2 s 525332 -800 525444 480 0 FreeSans 1120 90 0 0 la_oenb[112]
port 434 nsew signal input
flabel metal2 s 528878 -800 528990 480 0 FreeSans 1120 90 0 0 la_oenb[113]
port 435 nsew signal input
flabel metal2 s 532424 -800 532536 480 0 FreeSans 1120 90 0 0 la_oenb[114]
port 436 nsew signal input
flabel metal2 s 535970 -800 536082 480 0 FreeSans 1120 90 0 0 la_oenb[115]
port 437 nsew signal input
flabel metal2 s 539516 -800 539628 480 0 FreeSans 1120 90 0 0 la_oenb[116]
port 438 nsew signal input
flabel metal2 s 543062 -800 543174 480 0 FreeSans 1120 90 0 0 la_oenb[117]
port 439 nsew signal input
flabel metal2 s 546608 -800 546720 480 0 FreeSans 1120 90 0 0 la_oenb[118]
port 440 nsew signal input
flabel metal2 s 550154 -800 550266 480 0 FreeSans 1120 90 0 0 la_oenb[119]
port 441 nsew signal input
flabel metal2 s 167186 -800 167298 480 0 FreeSans 1120 90 0 0 la_oenb[11]
port 442 nsew signal input
flabel metal2 s 553700 -800 553812 480 0 FreeSans 1120 90 0 0 la_oenb[120]
port 443 nsew signal input
flabel metal2 s 557246 -800 557358 480 0 FreeSans 1120 90 0 0 la_oenb[121]
port 444 nsew signal input
flabel metal2 s 560792 -800 560904 480 0 FreeSans 1120 90 0 0 la_oenb[122]
port 445 nsew signal input
flabel metal2 s 564338 -800 564450 480 0 FreeSans 1120 90 0 0 la_oenb[123]
port 446 nsew signal input
flabel metal2 s 567884 -800 567996 480 0 FreeSans 1120 90 0 0 la_oenb[124]
port 447 nsew signal input
flabel metal2 s 571430 -800 571542 480 0 FreeSans 1120 90 0 0 la_oenb[125]
port 448 nsew signal input
flabel metal2 s 574976 -800 575088 480 0 FreeSans 1120 90 0 0 la_oenb[126]
port 449 nsew signal input
flabel metal2 s 578522 -800 578634 480 0 FreeSans 1120 90 0 0 la_oenb[127]
port 450 nsew signal input
flabel metal2 s 170732 -800 170844 480 0 FreeSans 1120 90 0 0 la_oenb[12]
port 451 nsew signal input
flabel metal2 s 174278 -800 174390 480 0 FreeSans 1120 90 0 0 la_oenb[13]
port 452 nsew signal input
flabel metal2 s 177824 -800 177936 480 0 FreeSans 1120 90 0 0 la_oenb[14]
port 453 nsew signal input
flabel metal2 s 181370 -800 181482 480 0 FreeSans 1120 90 0 0 la_oenb[15]
port 454 nsew signal input
flabel metal2 s 184916 -800 185028 480 0 FreeSans 1120 90 0 0 la_oenb[16]
port 455 nsew signal input
flabel metal2 s 188462 -800 188574 480 0 FreeSans 1120 90 0 0 la_oenb[17]
port 456 nsew signal input
flabel metal2 s 192008 -800 192120 480 0 FreeSans 1120 90 0 0 la_oenb[18]
port 457 nsew signal input
flabel metal2 s 195554 -800 195666 480 0 FreeSans 1120 90 0 0 la_oenb[19]
port 458 nsew signal input
flabel metal2 s 131726 -800 131838 480 0 FreeSans 1120 90 0 0 la_oenb[1]
port 459 nsew signal input
flabel metal2 s 199100 -800 199212 480 0 FreeSans 1120 90 0 0 la_oenb[20]
port 460 nsew signal input
flabel metal2 s 202646 -800 202758 480 0 FreeSans 1120 90 0 0 la_oenb[21]
port 461 nsew signal input
flabel metal2 s 206192 -800 206304 480 0 FreeSans 1120 90 0 0 la_oenb[22]
port 462 nsew signal input
flabel metal2 s 209738 -800 209850 480 0 FreeSans 1120 90 0 0 la_oenb[23]
port 463 nsew signal input
flabel metal2 s 213284 -800 213396 480 0 FreeSans 1120 90 0 0 la_oenb[24]
port 464 nsew signal input
flabel metal2 s 216830 -800 216942 480 0 FreeSans 1120 90 0 0 la_oenb[25]
port 465 nsew signal input
flabel metal2 s 220376 -800 220488 480 0 FreeSans 1120 90 0 0 la_oenb[26]
port 466 nsew signal input
flabel metal2 s 223922 -800 224034 480 0 FreeSans 1120 90 0 0 la_oenb[27]
port 467 nsew signal input
flabel metal2 s 227468 -800 227580 480 0 FreeSans 1120 90 0 0 la_oenb[28]
port 468 nsew signal input
flabel metal2 s 231014 -800 231126 480 0 FreeSans 1120 90 0 0 la_oenb[29]
port 469 nsew signal input
flabel metal2 s 135272 -800 135384 480 0 FreeSans 1120 90 0 0 la_oenb[2]
port 470 nsew signal input
flabel metal2 s 234560 -800 234672 480 0 FreeSans 1120 90 0 0 la_oenb[30]
port 471 nsew signal input
flabel metal2 s 238106 -800 238218 480 0 FreeSans 1120 90 0 0 la_oenb[31]
port 472 nsew signal input
flabel metal2 s 241652 -800 241764 480 0 FreeSans 1120 90 0 0 la_oenb[32]
port 473 nsew signal input
flabel metal2 s 245198 -800 245310 480 0 FreeSans 1120 90 0 0 la_oenb[33]
port 474 nsew signal input
flabel metal2 s 248744 -800 248856 480 0 FreeSans 1120 90 0 0 la_oenb[34]
port 475 nsew signal input
flabel metal2 s 252290 -800 252402 480 0 FreeSans 1120 90 0 0 la_oenb[35]
port 476 nsew signal input
flabel metal2 s 255836 -800 255948 480 0 FreeSans 1120 90 0 0 la_oenb[36]
port 477 nsew signal input
flabel metal2 s 259382 -800 259494 480 0 FreeSans 1120 90 0 0 la_oenb[37]
port 478 nsew signal input
flabel metal2 s 262928 -800 263040 480 0 FreeSans 1120 90 0 0 la_oenb[38]
port 479 nsew signal input
flabel metal2 s 266474 -800 266586 480 0 FreeSans 1120 90 0 0 la_oenb[39]
port 480 nsew signal input
flabel metal2 s 138818 -800 138930 480 0 FreeSans 1120 90 0 0 la_oenb[3]
port 481 nsew signal input
flabel metal2 s 270020 -800 270132 480 0 FreeSans 1120 90 0 0 la_oenb[40]
port 482 nsew signal input
flabel metal2 s 273566 -800 273678 480 0 FreeSans 1120 90 0 0 la_oenb[41]
port 483 nsew signal input
flabel metal2 s 277112 -800 277224 480 0 FreeSans 1120 90 0 0 la_oenb[42]
port 484 nsew signal input
flabel metal2 s 280658 -800 280770 480 0 FreeSans 1120 90 0 0 la_oenb[43]
port 485 nsew signal input
flabel metal2 s 284204 -800 284316 480 0 FreeSans 1120 90 0 0 la_oenb[44]
port 486 nsew signal input
flabel metal2 s 287750 -800 287862 480 0 FreeSans 1120 90 0 0 la_oenb[45]
port 487 nsew signal input
flabel metal2 s 291296 -800 291408 480 0 FreeSans 1120 90 0 0 la_oenb[46]
port 488 nsew signal input
flabel metal2 s 294842 -800 294954 480 0 FreeSans 1120 90 0 0 la_oenb[47]
port 489 nsew signal input
flabel metal2 s 298388 -800 298500 480 0 FreeSans 1120 90 0 0 la_oenb[48]
port 490 nsew signal input
flabel metal2 s 301934 -800 302046 480 0 FreeSans 1120 90 0 0 la_oenb[49]
port 491 nsew signal input
flabel metal2 s 142364 -800 142476 480 0 FreeSans 1120 90 0 0 la_oenb[4]
port 492 nsew signal input
flabel metal2 s 305480 -800 305592 480 0 FreeSans 1120 90 0 0 la_oenb[50]
port 493 nsew signal input
flabel metal2 s 309026 -800 309138 480 0 FreeSans 1120 90 0 0 la_oenb[51]
port 494 nsew signal input
flabel metal2 s 312572 -800 312684 480 0 FreeSans 1120 90 0 0 la_oenb[52]
port 495 nsew signal input
flabel metal2 s 316118 -800 316230 480 0 FreeSans 1120 90 0 0 la_oenb[53]
port 496 nsew signal input
flabel metal2 s 319664 -800 319776 480 0 FreeSans 1120 90 0 0 la_oenb[54]
port 497 nsew signal input
flabel metal2 s 323210 -800 323322 480 0 FreeSans 1120 90 0 0 la_oenb[55]
port 498 nsew signal input
flabel metal2 s 326756 -800 326868 480 0 FreeSans 1120 90 0 0 la_oenb[56]
port 499 nsew signal input
flabel metal2 s 330302 -800 330414 480 0 FreeSans 1120 90 0 0 la_oenb[57]
port 500 nsew signal input
flabel metal2 s 333848 -800 333960 480 0 FreeSans 1120 90 0 0 la_oenb[58]
port 501 nsew signal input
flabel metal2 s 337394 -800 337506 480 0 FreeSans 1120 90 0 0 la_oenb[59]
port 502 nsew signal input
flabel metal2 s 145910 -800 146022 480 0 FreeSans 1120 90 0 0 la_oenb[5]
port 503 nsew signal input
flabel metal2 s 340940 -800 341052 480 0 FreeSans 1120 90 0 0 la_oenb[60]
port 504 nsew signal input
flabel metal2 s 344486 -800 344598 480 0 FreeSans 1120 90 0 0 la_oenb[61]
port 505 nsew signal input
flabel metal2 s 348032 -800 348144 480 0 FreeSans 1120 90 0 0 la_oenb[62]
port 506 nsew signal input
flabel metal2 s 351578 -800 351690 480 0 FreeSans 1120 90 0 0 la_oenb[63]
port 507 nsew signal input
flabel metal2 s 355124 -800 355236 480 0 FreeSans 1120 90 0 0 la_oenb[64]
port 508 nsew signal input
flabel metal2 s 358670 -800 358782 480 0 FreeSans 1120 90 0 0 la_oenb[65]
port 509 nsew signal input
flabel metal2 s 362216 -800 362328 480 0 FreeSans 1120 90 0 0 la_oenb[66]
port 510 nsew signal input
flabel metal2 s 365762 -800 365874 480 0 FreeSans 1120 90 0 0 la_oenb[67]
port 511 nsew signal input
flabel metal2 s 369308 -800 369420 480 0 FreeSans 1120 90 0 0 la_oenb[68]
port 512 nsew signal input
flabel metal2 s 372854 -800 372966 480 0 FreeSans 1120 90 0 0 la_oenb[69]
port 513 nsew signal input
flabel metal2 s 149456 -800 149568 480 0 FreeSans 1120 90 0 0 la_oenb[6]
port 514 nsew signal input
flabel metal2 s 376400 -800 376512 480 0 FreeSans 1120 90 0 0 la_oenb[70]
port 515 nsew signal input
flabel metal2 s 379946 -800 380058 480 0 FreeSans 1120 90 0 0 la_oenb[71]
port 516 nsew signal input
flabel metal2 s 383492 -800 383604 480 0 FreeSans 1120 90 0 0 la_oenb[72]
port 517 nsew signal input
flabel metal2 s 387038 -800 387150 480 0 FreeSans 1120 90 0 0 la_oenb[73]
port 518 nsew signal input
flabel metal2 s 390584 -800 390696 480 0 FreeSans 1120 90 0 0 la_oenb[74]
port 519 nsew signal input
flabel metal2 s 394130 -800 394242 480 0 FreeSans 1120 90 0 0 la_oenb[75]
port 520 nsew signal input
flabel metal2 s 397676 -800 397788 480 0 FreeSans 1120 90 0 0 la_oenb[76]
port 521 nsew signal input
flabel metal2 s 401222 -800 401334 480 0 FreeSans 1120 90 0 0 la_oenb[77]
port 522 nsew signal input
flabel metal2 s 404768 -800 404880 480 0 FreeSans 1120 90 0 0 la_oenb[78]
port 523 nsew signal input
flabel metal2 s 408314 -800 408426 480 0 FreeSans 1120 90 0 0 la_oenb[79]
port 524 nsew signal input
flabel metal2 s 153002 -800 153114 480 0 FreeSans 1120 90 0 0 la_oenb[7]
port 525 nsew signal input
flabel metal2 s 411860 -800 411972 480 0 FreeSans 1120 90 0 0 la_oenb[80]
port 526 nsew signal input
flabel metal2 s 415406 -800 415518 480 0 FreeSans 1120 90 0 0 la_oenb[81]
port 527 nsew signal input
flabel metal2 s 418952 -800 419064 480 0 FreeSans 1120 90 0 0 la_oenb[82]
port 528 nsew signal input
flabel metal2 s 422498 -800 422610 480 0 FreeSans 1120 90 0 0 la_oenb[83]
port 529 nsew signal input
flabel metal2 s 426044 -800 426156 480 0 FreeSans 1120 90 0 0 la_oenb[84]
port 530 nsew signal input
flabel metal2 s 429590 -800 429702 480 0 FreeSans 1120 90 0 0 la_oenb[85]
port 531 nsew signal input
flabel metal2 s 433136 -800 433248 480 0 FreeSans 1120 90 0 0 la_oenb[86]
port 532 nsew signal input
flabel metal2 s 436682 -800 436794 480 0 FreeSans 1120 90 0 0 la_oenb[87]
port 533 nsew signal input
flabel metal2 s 440228 -800 440340 480 0 FreeSans 1120 90 0 0 la_oenb[88]
port 534 nsew signal input
flabel metal2 s 443774 -800 443886 480 0 FreeSans 1120 90 0 0 la_oenb[89]
port 535 nsew signal input
flabel metal2 s 156548 -800 156660 480 0 FreeSans 1120 90 0 0 la_oenb[8]
port 536 nsew signal input
flabel metal2 s 447320 -800 447432 480 0 FreeSans 1120 90 0 0 la_oenb[90]
port 537 nsew signal input
flabel metal2 s 450866 -800 450978 480 0 FreeSans 1120 90 0 0 la_oenb[91]
port 538 nsew signal input
flabel metal2 s 454412 -800 454524 480 0 FreeSans 1120 90 0 0 la_oenb[92]
port 539 nsew signal input
flabel metal2 s 457958 -800 458070 480 0 FreeSans 1120 90 0 0 la_oenb[93]
port 540 nsew signal input
flabel metal2 s 461504 -800 461616 480 0 FreeSans 1120 90 0 0 la_oenb[94]
port 541 nsew signal input
flabel metal2 s 465050 -800 465162 480 0 FreeSans 1120 90 0 0 la_oenb[95]
port 542 nsew signal input
flabel metal2 s 468596 -800 468708 480 0 FreeSans 1120 90 0 0 la_oenb[96]
port 543 nsew signal input
flabel metal2 s 472142 -800 472254 480 0 FreeSans 1120 90 0 0 la_oenb[97]
port 544 nsew signal input
flabel metal2 s 475688 -800 475800 480 0 FreeSans 1120 90 0 0 la_oenb[98]
port 545 nsew signal input
flabel metal2 s 479234 -800 479346 480 0 FreeSans 1120 90 0 0 la_oenb[99]
port 546 nsew signal input
flabel metal2 s 160094 -800 160206 480 0 FreeSans 1120 90 0 0 la_oenb[9]
port 547 nsew signal input
flabel metal2 s 579704 -800 579816 480 0 FreeSans 1120 90 0 0 user_clock2
port 548 nsew signal input
flabel metal2 s 580886 -800 580998 480 0 FreeSans 1120 90 0 0 user_irq[0]
port 549 nsew signal tristate
flabel metal2 s 582068 -800 582180 480 0 FreeSans 1120 90 0 0 user_irq[1]
port 550 nsew signal tristate
flabel metal2 s 583250 -800 583362 480 0 FreeSans 1120 90 0 0 user_irq[2]
port 551 nsew signal tristate
flabel metal3 s 582340 639784 584800 644584 0 FreeSans 1120 0 0 0 vccd1
port 552 nsew signal bidirectional
flabel metal3 s 582340 629784 584800 634584 0 FreeSans 1120 0 0 0 vccd1
port 553 nsew signal bidirectional
flabel metal3 s 0 643842 1660 648642 0 FreeSans 1120 0 0 0 vccd2
port 554 nsew signal bidirectional
flabel metal3 s 0 633842 1660 638642 0 FreeSans 1120 0 0 0 vccd2
port 555 nsew signal bidirectional
flabel metal3 s 582340 540562 584800 545362 0 FreeSans 1120 0 0 0 vdda1
port 556 nsew signal bidirectional
flabel metal3 s 582340 550562 584800 555362 0 FreeSans 1120 0 0 0 vdda1
port 557 nsew signal bidirectional
flabel metal3 s 582340 235230 584800 240030 0 FreeSans 1120 0 0 0 vdda1
port 558 nsew signal bidirectional
flabel metal3 s 582340 225230 584800 230030 0 FreeSans 1120 0 0 0 vdda1
port 559 nsew signal bidirectional
flabel metal3 s 0 204888 1660 209688 0 FreeSans 1120 0 0 0 vdda2
port 560 nsew signal bidirectional
flabel metal3 s 0 214888 1660 219688 0 FreeSans 1120 0 0 0 vdda2
port 561 nsew signal bidirectional
flabel metal3 s 520594 702340 525394 704800 0 FreeSans 1920 180 0 0 vssa1
port 562 nsew signal bidirectional
flabel metal3 s 510594 702340 515394 704800 0 FreeSans 1920 180 0 0 vssa1
port 563 nsew signal bidirectional
flabel metal3 s 582340 146830 584800 151630 0 FreeSans 1120 0 0 0 vssa1
port 564 nsew signal bidirectional
flabel metal3 s 582340 136830 584800 141630 0 FreeSans 1120 0 0 0 vssa1
port 565 nsew signal bidirectional
flabel metal3 s 0 559442 1660 564242 0 FreeSans 1120 0 0 0 vssa2
port 566 nsew signal bidirectional
flabel metal3 s 0 549442 1660 554242 0 FreeSans 1120 0 0 0 vssa2
port 567 nsew signal bidirectional
flabel metal3 s 582340 191430 584800 196230 0 FreeSans 1120 0 0 0 vssd1
port 568 nsew signal bidirectional
flabel metal3 s 582340 181430 584800 186230 0 FreeSans 1120 0 0 0 vssd1
port 569 nsew signal bidirectional
flabel metal3 s 0 172888 1660 177688 0 FreeSans 1120 0 0 0 vssd2
port 570 nsew signal bidirectional
flabel metal3 s 0 162888 1660 167688 0 FreeSans 1120 0 0 0 vssd2
port 571 nsew signal bidirectional
flabel metal2 s 524 -800 636 480 0 FreeSans 1120 90 0 0 wb_clk_i
port 572 nsew signal input
flabel metal2 s 1706 -800 1818 480 0 FreeSans 1120 90 0 0 wb_rst_i
port 573 nsew signal input
flabel metal2 s 2888 -800 3000 480 0 FreeSans 1120 90 0 0 wbs_ack_o
port 574 nsew signal tristate
flabel metal2 s 7616 -800 7728 480 0 FreeSans 1120 90 0 0 wbs_adr_i[0]
port 575 nsew signal input
flabel metal2 s 47804 -800 47916 480 0 FreeSans 1120 90 0 0 wbs_adr_i[10]
port 576 nsew signal input
flabel metal2 s 51350 -800 51462 480 0 FreeSans 1120 90 0 0 wbs_adr_i[11]
port 577 nsew signal input
flabel metal2 s 54896 -800 55008 480 0 FreeSans 1120 90 0 0 wbs_adr_i[12]
port 578 nsew signal input
flabel metal2 s 58442 -800 58554 480 0 FreeSans 1120 90 0 0 wbs_adr_i[13]
port 579 nsew signal input
flabel metal2 s 61988 -800 62100 480 0 FreeSans 1120 90 0 0 wbs_adr_i[14]
port 580 nsew signal input
flabel metal2 s 65534 -800 65646 480 0 FreeSans 1120 90 0 0 wbs_adr_i[15]
port 581 nsew signal input
flabel metal2 s 69080 -800 69192 480 0 FreeSans 1120 90 0 0 wbs_adr_i[16]
port 582 nsew signal input
flabel metal2 s 72626 -800 72738 480 0 FreeSans 1120 90 0 0 wbs_adr_i[17]
port 583 nsew signal input
flabel metal2 s 76172 -800 76284 480 0 FreeSans 1120 90 0 0 wbs_adr_i[18]
port 584 nsew signal input
flabel metal2 s 79718 -800 79830 480 0 FreeSans 1120 90 0 0 wbs_adr_i[19]
port 585 nsew signal input
flabel metal2 s 12344 -800 12456 480 0 FreeSans 1120 90 0 0 wbs_adr_i[1]
port 586 nsew signal input
flabel metal2 s 83264 -800 83376 480 0 FreeSans 1120 90 0 0 wbs_adr_i[20]
port 587 nsew signal input
flabel metal2 s 86810 -800 86922 480 0 FreeSans 1120 90 0 0 wbs_adr_i[21]
port 588 nsew signal input
flabel metal2 s 90356 -800 90468 480 0 FreeSans 1120 90 0 0 wbs_adr_i[22]
port 589 nsew signal input
flabel metal2 s 93902 -800 94014 480 0 FreeSans 1120 90 0 0 wbs_adr_i[23]
port 590 nsew signal input
flabel metal2 s 97448 -800 97560 480 0 FreeSans 1120 90 0 0 wbs_adr_i[24]
port 591 nsew signal input
flabel metal2 s 100994 -800 101106 480 0 FreeSans 1120 90 0 0 wbs_adr_i[25]
port 592 nsew signal input
flabel metal2 s 104540 -800 104652 480 0 FreeSans 1120 90 0 0 wbs_adr_i[26]
port 593 nsew signal input
flabel metal2 s 108086 -800 108198 480 0 FreeSans 1120 90 0 0 wbs_adr_i[27]
port 594 nsew signal input
flabel metal2 s 111632 -800 111744 480 0 FreeSans 1120 90 0 0 wbs_adr_i[28]
port 595 nsew signal input
flabel metal2 s 115178 -800 115290 480 0 FreeSans 1120 90 0 0 wbs_adr_i[29]
port 596 nsew signal input
flabel metal2 s 17072 -800 17184 480 0 FreeSans 1120 90 0 0 wbs_adr_i[2]
port 597 nsew signal input
flabel metal2 s 118724 -800 118836 480 0 FreeSans 1120 90 0 0 wbs_adr_i[30]
port 598 nsew signal input
flabel metal2 s 122270 -800 122382 480 0 FreeSans 1120 90 0 0 wbs_adr_i[31]
port 599 nsew signal input
flabel metal2 s 21800 -800 21912 480 0 FreeSans 1120 90 0 0 wbs_adr_i[3]
port 600 nsew signal input
flabel metal2 s 26528 -800 26640 480 0 FreeSans 1120 90 0 0 wbs_adr_i[4]
port 601 nsew signal input
flabel metal2 s 30074 -800 30186 480 0 FreeSans 1120 90 0 0 wbs_adr_i[5]
port 602 nsew signal input
flabel metal2 s 33620 -800 33732 480 0 FreeSans 1120 90 0 0 wbs_adr_i[6]
port 603 nsew signal input
flabel metal2 s 37166 -800 37278 480 0 FreeSans 1120 90 0 0 wbs_adr_i[7]
port 604 nsew signal input
flabel metal2 s 40712 -800 40824 480 0 FreeSans 1120 90 0 0 wbs_adr_i[8]
port 605 nsew signal input
flabel metal2 s 44258 -800 44370 480 0 FreeSans 1120 90 0 0 wbs_adr_i[9]
port 606 nsew signal input
flabel metal2 s 4070 -800 4182 480 0 FreeSans 1120 90 0 0 wbs_cyc_i
port 607 nsew signal input
flabel metal2 s 8798 -800 8910 480 0 FreeSans 1120 90 0 0 wbs_dat_i[0]
port 608 nsew signal input
flabel metal2 s 48986 -800 49098 480 0 FreeSans 1120 90 0 0 wbs_dat_i[10]
port 609 nsew signal input
flabel metal2 s 52532 -800 52644 480 0 FreeSans 1120 90 0 0 wbs_dat_i[11]
port 610 nsew signal input
flabel metal2 s 56078 -800 56190 480 0 FreeSans 1120 90 0 0 wbs_dat_i[12]
port 611 nsew signal input
flabel metal2 s 59624 -800 59736 480 0 FreeSans 1120 90 0 0 wbs_dat_i[13]
port 612 nsew signal input
flabel metal2 s 63170 -800 63282 480 0 FreeSans 1120 90 0 0 wbs_dat_i[14]
port 613 nsew signal input
flabel metal2 s 66716 -800 66828 480 0 FreeSans 1120 90 0 0 wbs_dat_i[15]
port 614 nsew signal input
flabel metal2 s 70262 -800 70374 480 0 FreeSans 1120 90 0 0 wbs_dat_i[16]
port 615 nsew signal input
flabel metal2 s 73808 -800 73920 480 0 FreeSans 1120 90 0 0 wbs_dat_i[17]
port 616 nsew signal input
flabel metal2 s 77354 -800 77466 480 0 FreeSans 1120 90 0 0 wbs_dat_i[18]
port 617 nsew signal input
flabel metal2 s 80900 -800 81012 480 0 FreeSans 1120 90 0 0 wbs_dat_i[19]
port 618 nsew signal input
flabel metal2 s 13526 -800 13638 480 0 FreeSans 1120 90 0 0 wbs_dat_i[1]
port 619 nsew signal input
flabel metal2 s 84446 -800 84558 480 0 FreeSans 1120 90 0 0 wbs_dat_i[20]
port 620 nsew signal input
flabel metal2 s 87992 -800 88104 480 0 FreeSans 1120 90 0 0 wbs_dat_i[21]
port 621 nsew signal input
flabel metal2 s 91538 -800 91650 480 0 FreeSans 1120 90 0 0 wbs_dat_i[22]
port 622 nsew signal input
flabel metal2 s 95084 -800 95196 480 0 FreeSans 1120 90 0 0 wbs_dat_i[23]
port 623 nsew signal input
flabel metal2 s 98630 -800 98742 480 0 FreeSans 1120 90 0 0 wbs_dat_i[24]
port 624 nsew signal input
flabel metal2 s 102176 -800 102288 480 0 FreeSans 1120 90 0 0 wbs_dat_i[25]
port 625 nsew signal input
flabel metal2 s 105722 -800 105834 480 0 FreeSans 1120 90 0 0 wbs_dat_i[26]
port 626 nsew signal input
flabel metal2 s 109268 -800 109380 480 0 FreeSans 1120 90 0 0 wbs_dat_i[27]
port 627 nsew signal input
flabel metal2 s 112814 -800 112926 480 0 FreeSans 1120 90 0 0 wbs_dat_i[28]
port 628 nsew signal input
flabel metal2 s 116360 -800 116472 480 0 FreeSans 1120 90 0 0 wbs_dat_i[29]
port 629 nsew signal input
flabel metal2 s 18254 -800 18366 480 0 FreeSans 1120 90 0 0 wbs_dat_i[2]
port 630 nsew signal input
flabel metal2 s 119906 -800 120018 480 0 FreeSans 1120 90 0 0 wbs_dat_i[30]
port 631 nsew signal input
flabel metal2 s 123452 -800 123564 480 0 FreeSans 1120 90 0 0 wbs_dat_i[31]
port 632 nsew signal input
flabel metal2 s 22982 -800 23094 480 0 FreeSans 1120 90 0 0 wbs_dat_i[3]
port 633 nsew signal input
flabel metal2 s 27710 -800 27822 480 0 FreeSans 1120 90 0 0 wbs_dat_i[4]
port 634 nsew signal input
flabel metal2 s 31256 -800 31368 480 0 FreeSans 1120 90 0 0 wbs_dat_i[5]
port 635 nsew signal input
flabel metal2 s 34802 -800 34914 480 0 FreeSans 1120 90 0 0 wbs_dat_i[6]
port 636 nsew signal input
flabel metal2 s 38348 -800 38460 480 0 FreeSans 1120 90 0 0 wbs_dat_i[7]
port 637 nsew signal input
flabel metal2 s 41894 -800 42006 480 0 FreeSans 1120 90 0 0 wbs_dat_i[8]
port 638 nsew signal input
flabel metal2 s 45440 -800 45552 480 0 FreeSans 1120 90 0 0 wbs_dat_i[9]
port 639 nsew signal input
flabel metal2 s 9980 -800 10092 480 0 FreeSans 1120 90 0 0 wbs_dat_o[0]
port 640 nsew signal tristate
flabel metal2 s 50168 -800 50280 480 0 FreeSans 1120 90 0 0 wbs_dat_o[10]
port 641 nsew signal tristate
flabel metal2 s 53714 -800 53826 480 0 FreeSans 1120 90 0 0 wbs_dat_o[11]
port 642 nsew signal tristate
flabel metal2 s 57260 -800 57372 480 0 FreeSans 1120 90 0 0 wbs_dat_o[12]
port 643 nsew signal tristate
flabel metal2 s 60806 -800 60918 480 0 FreeSans 1120 90 0 0 wbs_dat_o[13]
port 644 nsew signal tristate
flabel metal2 s 64352 -800 64464 480 0 FreeSans 1120 90 0 0 wbs_dat_o[14]
port 645 nsew signal tristate
flabel metal2 s 67898 -800 68010 480 0 FreeSans 1120 90 0 0 wbs_dat_o[15]
port 646 nsew signal tristate
flabel metal2 s 71444 -800 71556 480 0 FreeSans 1120 90 0 0 wbs_dat_o[16]
port 647 nsew signal tristate
flabel metal2 s 74990 -800 75102 480 0 FreeSans 1120 90 0 0 wbs_dat_o[17]
port 648 nsew signal tristate
flabel metal2 s 78536 -800 78648 480 0 FreeSans 1120 90 0 0 wbs_dat_o[18]
port 649 nsew signal tristate
flabel metal2 s 82082 -800 82194 480 0 FreeSans 1120 90 0 0 wbs_dat_o[19]
port 650 nsew signal tristate
flabel metal2 s 14708 -800 14820 480 0 FreeSans 1120 90 0 0 wbs_dat_o[1]
port 651 nsew signal tristate
flabel metal2 s 85628 -800 85740 480 0 FreeSans 1120 90 0 0 wbs_dat_o[20]
port 652 nsew signal tristate
flabel metal2 s 89174 -800 89286 480 0 FreeSans 1120 90 0 0 wbs_dat_o[21]
port 653 nsew signal tristate
flabel metal2 s 92720 -800 92832 480 0 FreeSans 1120 90 0 0 wbs_dat_o[22]
port 654 nsew signal tristate
flabel metal2 s 96266 -800 96378 480 0 FreeSans 1120 90 0 0 wbs_dat_o[23]
port 655 nsew signal tristate
flabel metal2 s 99812 -800 99924 480 0 FreeSans 1120 90 0 0 wbs_dat_o[24]
port 656 nsew signal tristate
flabel metal2 s 103358 -800 103470 480 0 FreeSans 1120 90 0 0 wbs_dat_o[25]
port 657 nsew signal tristate
flabel metal2 s 106904 -800 107016 480 0 FreeSans 1120 90 0 0 wbs_dat_o[26]
port 658 nsew signal tristate
flabel metal2 s 110450 -800 110562 480 0 FreeSans 1120 90 0 0 wbs_dat_o[27]
port 659 nsew signal tristate
flabel metal2 s 113996 -800 114108 480 0 FreeSans 1120 90 0 0 wbs_dat_o[28]
port 660 nsew signal tristate
flabel metal2 s 117542 -800 117654 480 0 FreeSans 1120 90 0 0 wbs_dat_o[29]
port 661 nsew signal tristate
flabel metal2 s 19436 -800 19548 480 0 FreeSans 1120 90 0 0 wbs_dat_o[2]
port 662 nsew signal tristate
flabel metal2 s 121088 -800 121200 480 0 FreeSans 1120 90 0 0 wbs_dat_o[30]
port 663 nsew signal tristate
flabel metal2 s 124634 -800 124746 480 0 FreeSans 1120 90 0 0 wbs_dat_o[31]
port 664 nsew signal tristate
flabel metal2 s 24164 -800 24276 480 0 FreeSans 1120 90 0 0 wbs_dat_o[3]
port 665 nsew signal tristate
flabel metal2 s 28892 -800 29004 480 0 FreeSans 1120 90 0 0 wbs_dat_o[4]
port 666 nsew signal tristate
flabel metal2 s 32438 -800 32550 480 0 FreeSans 1120 90 0 0 wbs_dat_o[5]
port 667 nsew signal tristate
flabel metal2 s 35984 -800 36096 480 0 FreeSans 1120 90 0 0 wbs_dat_o[6]
port 668 nsew signal tristate
flabel metal2 s 39530 -800 39642 480 0 FreeSans 1120 90 0 0 wbs_dat_o[7]
port 669 nsew signal tristate
flabel metal2 s 43076 -800 43188 480 0 FreeSans 1120 90 0 0 wbs_dat_o[8]
port 670 nsew signal tristate
flabel metal2 s 46622 -800 46734 480 0 FreeSans 1120 90 0 0 wbs_dat_o[9]
port 671 nsew signal tristate
flabel metal2 s 11162 -800 11274 480 0 FreeSans 1120 90 0 0 wbs_sel_i[0]
port 672 nsew signal input
flabel metal2 s 15890 -800 16002 480 0 FreeSans 1120 90 0 0 wbs_sel_i[1]
port 673 nsew signal input
flabel metal2 s 20618 -800 20730 480 0 FreeSans 1120 90 0 0 wbs_sel_i[2]
port 674 nsew signal input
flabel metal2 s 25346 -800 25458 480 0 FreeSans 1120 90 0 0 wbs_sel_i[3]
port 675 nsew signal input
flabel metal2 s 5252 -800 5364 480 0 FreeSans 1120 90 0 0 wbs_stb_i
port 676 nsew signal input
flabel metal2 s 6434 -800 6546 480 0 FreeSans 1120 90 0 0 wbs_we_i
port 677 nsew signal input
flabel metal3 572152 640142 580220 644150 0 FreeSans 16000 0 0 0 VCCD1
flabel metal3 567038 550960 577302 554546 0 FreeSans 16000 0 0 0 VDDA1
flabel metal3 511190 664896 514962 676272 0 FreeSans 16000 90 0 0 VSSA1
flabel metal3 561703 191929 571721 195859 0 FreeSans 16000 0 0 0 VSSD1
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
