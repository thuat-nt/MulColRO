magic
tech sky130A
magscale 1 2
timestamp 1696663834
<< locali >>
rect 15024 33870 16026 33956
rect 15024 32316 15094 33870
rect 15952 32316 16026 33870
rect 15024 12840 16026 32316
rect 20978 33782 21856 33892
rect 20978 32230 21072 33782
rect 21730 32230 21856 33782
rect 20978 7178 21856 32230
rect 35070 14078 36124 14218
rect 35070 13732 35278 14078
rect 35988 13732 36124 14078
rect 35070 13152 36124 13732
rect 35070 9588 36820 13152
rect 19378 -4796 20292 3040
rect 20858 -4796 21794 5776
rect 35070 4060 36124 9588
rect 47350 5426 50654 5440
rect 47350 5354 50706 5426
rect 47350 4580 47460 5354
rect 47976 4580 50706 5354
rect 47350 4492 50706 4580
rect 19376 -6136 21794 -4796
rect 35048 2518 36128 4060
rect 35048 1920 37074 2518
rect 35048 -1158 36128 1920
rect 35048 -1748 35172 -1158
rect 36030 -1748 36128 -1158
rect 35048 -5018 36128 -1748
rect 35028 -6136 36128 -5018
rect 49206 -5298 50706 4492
rect 19376 -6564 21750 -6136
rect 19376 -7296 19578 -6564
rect 21474 -7296 21750 -6564
rect 19376 -7420 21750 -7296
rect 35028 -6536 36104 -6136
rect 35028 -7242 35154 -6536
rect 35874 -7242 36104 -6536
rect 35028 -7448 36104 -7242
<< viali >>
rect 15094 32316 15952 33870
rect 21072 32230 21730 33782
rect 35278 13732 35988 14078
rect 47460 4580 47976 5354
rect 35172 -1748 36030 -1158
rect 19578 -7296 21474 -6564
rect 35154 -7242 35874 -6536
<< metal1 >>
rect 15054 33870 16000 33918
rect 15054 32316 15094 33870
rect 15952 32316 16000 33870
rect 15054 32232 16000 32316
rect 20852 33782 21926 33962
rect 20852 32230 21072 33782
rect 21730 32230 21926 33782
rect 20852 32198 21926 32230
rect 24116 33516 25278 33622
rect 24116 32264 24224 33516
rect 25188 32264 25278 33516
rect 24116 13726 25278 32264
rect 45892 33406 47008 33494
rect 45892 32264 45980 33406
rect 46904 32264 47008 33406
rect 34120 14078 36970 31590
rect 34120 13732 35278 14078
rect 35988 13732 36970 14078
rect 24116 13712 33790 13726
rect 24116 13504 33816 13712
rect 34120 13528 36970 13732
rect 33204 13126 33816 13504
rect 23816 4806 24178 5548
rect 22950 2730 24178 4806
rect 32920 -5816 34128 4972
rect 35888 4516 36952 13528
rect 45892 5554 47008 32264
rect 45892 5354 48080 5554
rect 45892 4580 47460 5354
rect 47976 4580 48080 5354
rect 45892 4506 48080 4580
rect 45910 4414 48080 4506
rect 35042 -1158 36108 -1020
rect 35042 -1748 35172 -1158
rect 36030 -1748 36108 -1158
rect 35042 -1886 36108 -1748
rect 19412 -6564 21708 -6412
rect 19412 -7296 19578 -6564
rect 21474 -7296 21708 -6564
rect 19412 -7420 21708 -7296
rect 34932 -6536 36094 -6398
rect 34932 -7242 35154 -6536
rect 35874 -7242 36094 -6536
rect 34932 -7448 36094 -7242
<< via1 >>
rect 15094 32316 15952 33870
rect 21072 32230 21730 33782
rect 24224 32264 25188 33516
rect 45980 32264 46904 33406
rect 22222 6310 22362 6456
rect 23548 -2018 23910 -962
rect 35172 -1748 36030 -1158
rect 19578 -7296 21474 -6564
rect 35154 -7242 35874 -6536
<< metal2 >>
rect 14628 33870 57258 36292
rect 14628 32316 15094 33870
rect 15952 33782 57258 33870
rect 15952 32316 21072 33782
rect 14628 32230 21072 32316
rect 21730 33516 57258 33782
rect 21730 32264 24224 33516
rect 25188 33406 57258 33516
rect 25188 32264 45980 33406
rect 46904 32264 57258 33406
rect 21730 32230 57258 32264
rect 14628 32156 57258 32230
rect 16718 9180 17114 9292
rect 16718 8572 16762 9180
rect 17070 8572 17114 9180
rect 16718 8460 17114 8572
rect 22200 6456 22376 6472
rect 22200 6310 22222 6456
rect 22362 6310 22376 6456
rect 22200 6290 22376 6310
rect 16844 2090 17410 2230
rect 16844 1868 16970 2090
rect 17302 1868 17410 2090
rect 16844 1720 17410 1868
rect 22858 -962 24172 2862
rect 25058 -200 26320 7816
rect 31452 3880 39416 31570
rect 43930 18196 56166 18372
rect 43930 17776 55314 18196
rect 56030 17776 56166 18196
rect 43930 17516 56166 17776
rect 22858 -2018 23548 -962
rect 23910 -2018 24172 -962
rect 35042 -1158 36108 -1020
rect 35042 -1748 35172 -1158
rect 36030 -1748 36108 -1158
rect 35042 -1886 36108 -1748
rect 22858 -4916 24172 -2018
rect 36202 -2642 36780 3880
rect 22856 -6136 24172 -4916
rect 14946 -6536 57118 -6394
rect 14946 -6564 35154 -6536
rect 14946 -7296 19578 -6564
rect 21474 -7242 35154 -6564
rect 35874 -7242 57118 -6536
rect 21474 -7296 57118 -7242
rect 14946 -10124 57118 -7296
<< via2 >>
rect 30942 27254 31096 27416
rect 26260 23556 27224 24248
rect 30930 18268 31106 18436
rect 26148 14606 27300 15542
rect 16762 8572 17070 9180
rect 25368 8598 25938 9180
rect 27202 8670 27364 8830
rect 21122 6370 21222 6454
rect 22236 6330 22348 6438
rect 16970 1868 17302 2090
rect 39996 27186 40162 27404
rect 44146 27008 44952 27430
rect 39952 17902 40124 18066
rect 55314 17776 56030 18196
rect 40068 8796 40228 8974
rect 44222 8624 45018 9066
rect 27102 -1626 27260 -1470
rect 31500 -1652 31890 -1280
rect 35172 -1748 36030 -1158
rect 41928 -2498 42036 -2434
rect 37518 -4376 37628 -4258
<< metal3 >>
rect 20978 30292 21706 30304
rect 20550 29986 22164 30292
rect 20550 28896 40436 29986
rect 20550 28632 22164 28896
rect 20978 28630 21706 28632
rect 20978 28072 21706 28078
rect 20572 27644 22186 28072
rect 20572 27416 31334 27644
rect 20572 27254 30942 27416
rect 31096 27254 31334 27416
rect 20572 26824 31334 27254
rect 39788 27404 40430 28896
rect 39788 27186 39996 27404
rect 40162 27186 40430 27404
rect 39788 27068 40430 27186
rect 44044 27430 45012 27488
rect 44044 27008 44146 27430
rect 44952 27008 45012 27430
rect 44044 26942 45012 27008
rect 20572 26412 22186 26824
rect 20978 26326 21706 26412
rect 26150 24248 27368 24346
rect 26150 23556 26260 24248
rect 27224 23556 27368 24248
rect 26150 23446 27368 23556
rect 20978 21304 21706 21354
rect 20594 20878 22208 21304
rect 20594 20000 40506 20878
rect 20594 19644 22208 20000
rect 20978 19632 21706 19644
rect 20978 19130 21706 19140
rect 20616 18664 22230 19130
rect 20616 18436 31258 18664
rect 20616 18268 30930 18436
rect 31106 18268 31258 18436
rect 20616 17856 31258 18268
rect 39654 18066 40490 20000
rect 39654 17902 39952 18066
rect 40124 17902 40490 18066
rect 20616 17470 22230 17856
rect 39654 17780 40490 17902
rect 55248 18196 56070 18248
rect 55248 17776 55314 18196
rect 56030 17776 56070 18196
rect 55248 17704 56070 17776
rect 20978 17454 21706 17470
rect 20932 17000 21984 17002
rect 20616 15340 22230 17000
rect 26094 15542 27478 15704
rect 20932 12410 21984 15340
rect 26094 14606 26148 15542
rect 27300 14606 27478 15542
rect 26094 14498 27478 14606
rect 20932 11616 40604 12410
rect 16744 9180 17092 9258
rect 16744 8572 16762 9180
rect 17070 8572 17092 9180
rect 16744 8506 17092 8572
rect 25252 9180 25996 9236
rect 25252 8598 25368 9180
rect 25938 8598 25996 9180
rect 39810 8974 40588 11616
rect 25252 8518 25996 8598
rect 27126 8830 27436 8888
rect 27126 8670 27202 8830
rect 27364 8670 27436 8830
rect 20890 6454 21304 6548
rect 27126 6498 27436 8670
rect 39810 8796 40068 8974
rect 40228 8796 40588 8974
rect 39810 8628 40588 8796
rect 44166 9066 45096 9160
rect 44166 8624 44222 9066
rect 45018 8624 45096 9066
rect 44166 8552 45096 8624
rect 20890 6370 21122 6454
rect 21222 6370 21304 6454
rect 16844 2090 17410 2230
rect 16844 1868 16970 2090
rect 17302 1868 17410 2090
rect 16844 1720 17410 1868
rect 20890 -902 21304 6370
rect 22180 6438 27460 6498
rect 22180 6330 22236 6438
rect 22348 6330 27460 6438
rect 22180 6258 27460 6330
rect 20636 -1196 21666 -902
rect 31352 -1108 32016 -1102
rect 20636 -1238 22676 -1196
rect 20636 -1250 22884 -1238
rect 24072 -1250 24426 -1238
rect 26880 -1250 27316 -1238
rect 20636 -1470 27318 -1250
rect 20636 -1626 27102 -1470
rect 27260 -1626 27318 -1470
rect 20636 -1924 27318 -1626
rect 31352 -1280 32018 -1108
rect 31352 -1652 31500 -1280
rect 31890 -1652 32018 -1280
rect 31352 -1894 32018 -1652
rect 35042 -1158 36108 -1020
rect 35042 -1748 35172 -1158
rect 36030 -1748 36108 -1158
rect 35042 -1886 36108 -1748
rect 31368 -1896 32018 -1894
rect 20636 -2074 21666 -1924
rect 22616 -1934 27318 -1924
rect 41868 -2234 42188 -2158
rect 41868 -2552 41898 -2234
rect 42136 -2552 42188 -2234
rect 41868 -2564 42188 -2552
rect 35964 -4114 37728 -4064
rect 35954 -4258 37728 -4114
rect 35954 -4376 37518 -4258
rect 37628 -4376 37728 -4258
rect 35954 -4586 37728 -4376
rect 35658 -4606 37728 -4586
rect 35658 -5760 36862 -4606
<< via3 >>
rect 44146 27008 44952 27430
rect 26260 23556 27224 24248
rect 55362 17824 55974 18154
rect 26148 14606 27300 15542
rect 16792 8698 17056 9048
rect 25490 8630 25844 9028
rect 44222 8624 45018 9066
rect 31512 -1646 31866 -1312
rect 35172 -1748 36030 -1158
rect 41898 -2434 42136 -2234
rect 41898 -2498 41928 -2434
rect 41928 -2498 42036 -2434
rect 42036 -2498 42136 -2434
rect 41898 -2552 42136 -2498
<< metal4 >>
rect 43928 27430 50272 27584
rect 43928 27008 44146 27430
rect 44952 27008 50272 27430
rect 43928 26774 50272 27008
rect 26058 24248 50282 24536
rect 26058 23556 26260 24248
rect 27224 23556 50282 24248
rect 26058 23260 50282 23556
rect 54812 18154 57228 31570
rect 54772 17824 55362 18154
rect 55974 17824 57228 18154
rect 16328 15236 18180 17016
rect 25976 15542 50196 15820
rect 16720 9332 17814 15236
rect 25976 14606 26148 15542
rect 27300 14606 50196 15542
rect 25976 14396 50196 14606
rect 16682 9048 26064 9332
rect 16682 8698 16792 9048
rect 17056 9028 26064 9048
rect 17056 8698 25490 9028
rect 16682 8630 25490 8698
rect 25844 8630 26064 9028
rect 16682 8386 26064 8630
rect 44038 9066 50258 9232
rect 44038 8624 44222 9066
rect 45018 8624 50258 9066
rect 44038 8436 50258 8624
rect 54812 6018 57228 17824
rect 54834 1498 57198 6018
rect 53568 1454 57198 1498
rect 46982 1092 57198 1454
rect 46982 1082 54970 1092
rect 53568 1048 54970 1082
rect 31368 -1158 42344 -1066
rect 31368 -1312 35172 -1158
rect 31368 -1646 31512 -1312
rect 31866 -1646 35172 -1312
rect 31368 -1748 35172 -1646
rect 36030 -1646 42344 -1158
rect 36030 -1748 42348 -1646
rect 31368 -1868 42348 -1748
rect 41794 -2234 42348 -1868
rect 41794 -2552 41898 -2234
rect 42136 -2552 42348 -2234
rect 41794 -2600 42348 -2552
use switch  x1
timestamp 1696663202
transform 0 1 36806 1 0 4546
box -53 -918 8642 10274
use switch  x2
timestamp 1696663202
transform 0 1 23934 -1 0 13086
box -53 -918 8642 10274
use curr_mir  x3
timestamp 1696147843
transform 0 -1 25426 1 0 1738
box 400 5130 11334 10390
use opamp  x4
timestamp 1696521366
transform 1 0 30358 0 -1 3752
box 6068 1244 19288 9014
use switch  x5
timestamp 1696663202
transform 0 1 36696 1 0 13644
box -53 -918 8642 10274
use switch  x6
timestamp 1696663202
transform 0 1 23834 -1 0 2788
box -53 -918 8642 10274
use not  x7
timestamp 1696661316
transform 1 0 20524 0 1 6226
box 472 -578 1868 1036
use switch  x8
timestamp 1696663202
transform 0 1 36738 1 0 22948
box -53 -918 8642 10274
use switch  x9
timestamp 1696663202
transform 0 -1 34358 1 0 14018
box -53 -918 8642 10274
use switch  x10
timestamp 1696663202
transform 0 -1 34358 1 0 22992
box -53 -918 8642 10274
use sky130_fd_pr__cap_mim_m3_1_3HBNLG  XC1
timestamp 1695395215
transform 1 0 51852 0 1 8768
box -3186 -3040 3186 3040
use sky130_fd_pr__cap_mim_m3_1_3HBNLG  XC2
timestamp 1695395215
transform 1 0 51818 0 1 15410
box -3186 -3040 3186 3040
use sky130_fd_pr__cap_mim_m3_1_3HBNLG  XC3
timestamp 1695395215
transform 1 0 51832 0 1 22082
box -3186 -3040 3186 3040
use sky130_fd_pr__cap_mim_m3_1_3HBNLG  XC4
timestamp 1695395215
transform 1 0 51864 0 1 28446
box -3186 -3040 3186 3040
<< labels >>
rlabel metal4 54834 1092 57198 17824 1 intout
port 7 nsew
rlabel metal3 35658 -5760 36862 -4586 1 opbias
port 13 nsew
rlabel metal3 20636 -2074 21666 -902 1 en
port 14 nsew
rlabel metal3 16844 1720 17410 2230 1 Vtune
port 15 nsew
rlabel metal4 16328 15236 18180 17016 1 intin
port 16 nsew
rlabel metal2 14946 -10124 57118 -6394 1 GROUND
port 18 nsew
rlabel metal2 14628 32156 57258 36292 1 VDD
port 17 nsew
rlabel metal3 20616 15340 22230 17000 1 sw1
port 12 nsew
rlabel metal3 20616 17470 22230 19130 1 sw2
port 11 nsew
rlabel metal3 20594 19644 22208 21304 1 rst
port 10 nsew
rlabel metal3 20572 26412 22186 28072 1 sw3
port 9 nsew
rlabel metal3 20550 28632 22164 30292 1 sw4
port 8 nsew
<< end >>
