magic
tech sky130A
magscale 1 2
timestamp 1698982829
<< metal3 >>
rect -386 412 386 440
rect -386 -412 302 412
rect 366 -412 386 412
rect -386 -440 386 -412
<< via3 >>
rect 302 -412 366 412
<< mimcap >>
rect -346 360 54 400
rect -346 -360 -306 360
rect 14 -360 54 360
rect -346 -400 54 -360
<< mimcapcontact >>
rect -306 -360 14 360
<< metal4 >>
rect 286 412 382 428
rect -307 360 15 361
rect -307 -360 -306 360
rect 14 -360 15 360
rect -307 -361 15 -360
rect 286 -412 302 412
rect 366 -412 382 412
rect 286 -428 382 -412
<< labels >>
rlabel mimcapcontact -306 -360 14 360 1 c0
port 1 nsew
rlabel via3 302 -412 366 412 1 c1
port 2 nsew
<< properties >>
string FIXED_BBOX -386 -440 94 440
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 2.0 l 4.0 val 18.28 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
