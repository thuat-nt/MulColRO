magic
tech sky130A
magscale 1 2
timestamp 1696148011
<< metal1 >>
rect 18616 30570 19744 30738
rect 5194 30338 5408 30390
rect 5194 30126 5242 30338
rect 5346 30126 5408 30338
rect 4402 16504 4670 16562
rect 4402 16386 4474 16504
rect 4596 16386 4670 16504
rect 4402 12478 4670 16386
rect 5194 12546 5408 30126
rect 18616 30216 18876 30570
rect 19496 30216 19744 30570
rect 6416 26036 6616 26060
rect 6416 25876 6428 26036
rect 6594 25876 6616 26036
rect 6416 25860 6616 25876
rect 5924 13738 6142 25550
rect 6464 16978 6664 16994
rect 6464 16806 6476 16978
rect 6648 16806 6664 16978
rect 6464 16794 6664 16806
rect 5914 12478 6108 12782
rect 4402 12464 6108 12478
rect 4402 12268 6114 12464
rect 5914 12264 6114 12268
rect 6544 11744 6754 12794
rect 6544 11532 6590 11744
rect 6694 11532 6754 11744
rect 6544 11480 6754 11532
rect 7414 11738 8536 22004
rect 18616 12220 19744 30216
rect 20522 20994 20722 21012
rect 20522 20832 20538 20994
rect 20706 20832 20722 20994
rect 20522 20812 20722 20832
rect 7414 11262 7642 11738
rect 8320 11262 8536 11738
rect 7414 11176 8536 11262
<< via1 >>
rect 5242 30126 5346 30338
rect 4474 16386 4596 16504
rect 18876 30216 19496 30570
rect 6428 25876 6594 26036
rect 6476 16806 6648 16978
rect 6590 11532 6694 11744
rect 20538 20832 20706 20994
rect 7642 11262 8320 11738
<< metal2 >>
rect 4240 30570 20872 33492
rect 4240 30338 18876 30570
rect 4240 30126 5242 30338
rect 5346 30216 18876 30338
rect 19496 30216 20872 30570
rect 5346 30126 20872 30216
rect 4240 30074 20872 30126
rect 6114 26036 10540 28732
rect 6114 25876 6428 26036
rect 6594 25876 10540 26036
rect 6114 25632 10540 25876
rect 5894 25484 6188 25538
rect 5894 25364 5976 25484
rect 6090 25364 6188 25484
rect 5894 25318 6188 25364
rect 11546 25516 11782 25550
rect 11546 25358 11580 25516
rect 11760 25358 11782 25516
rect 11546 25334 11782 25358
rect 15754 20994 20790 29664
rect 15754 20832 20538 20994
rect 20706 20832 20790 20994
rect 6130 16978 10556 19736
rect 6130 16806 6476 16978
rect 6648 16806 10556 16978
rect 6130 16636 10556 16806
rect 4384 16504 4702 16550
rect 4384 16386 4474 16504
rect 4596 16386 4702 16504
rect 4384 16330 4702 16386
rect 11578 16490 11778 16538
rect 11578 16358 11610 16490
rect 11752 16358 11778 16490
rect 11578 16288 11778 16358
rect 15754 12268 20790 20832
rect 4200 11744 20832 11840
rect 4200 11532 6590 11744
rect 6694 11738 20832 11744
rect 6694 11532 7642 11738
rect 4200 11262 7642 11532
rect 8320 11262 20832 11738
rect 4200 8422 20832 11262
<< via2 >>
rect 5976 25364 6090 25484
rect 11580 25358 11760 25516
rect 4474 16386 4596 16504
rect 11610 16358 11752 16490
<< metal3 >>
rect 5894 25516 11804 25562
rect 5894 25484 11580 25516
rect 5894 25364 5976 25484
rect 6090 25364 11580 25484
rect 5894 25358 11580 25364
rect 11760 25358 11804 25516
rect 5894 25312 11804 25358
rect 11550 16558 11810 16566
rect 4360 16504 11810 16558
rect 4360 16386 4474 16504
rect 4596 16490 11810 16504
rect 4596 16386 11610 16490
rect 4360 16358 11610 16386
rect 11752 16358 11810 16490
rect 4360 16308 11810 16358
rect 11550 16282 11810 16308
use not  x1
timestamp 1696147843
transform 0 -1 6186 1 0 12070
box 476 -578 1868 990
use switch  x5
timestamp 1696147897
transform 0 1 8322 -1 0 29778
box -53 -918 8642 11418
use switch  x6
timestamp 1696147897
transform 0 1 8340 -1 0 20784
box -53 -918 8642 11418
<< labels >>
flabel metal1 5914 12264 6114 12464 0 FreeSans 256 0 0 0 SEL0
port 0 nsew
flabel metal1 6416 25860 6616 26060 0 FreeSans 256 0 0 0 IN0
port 3 nsew
flabel metal1 6464 16794 6664 16994 0 FreeSans 256 0 0 0 IN1
port 1 nsew
flabel metal1 20522 20812 20722 21012 0 FreeSans 256 0 0 0 OUT
port 2 nsew
rlabel metal2 4200 8422 20832 11840 1 GROUND
port 4 nsew
rlabel metal2 4240 30074 20872 33492 1 VDD
port 5 nsew
rlabel metal2 10488 9224 13228 10790 1 GROUND
rlabel metal2 10988 30990 13728 32556 1 VDD
<< end >>
