magic
tech sky130A
magscale 1 2
timestamp 1695803350
<< locali >>
rect 28544 3482 30676 3802
rect 28544 1906 28840 3482
rect 30322 1906 30676 3482
rect 28544 -5660 30676 1906
rect 31294 -184 58150 1392
rect 31140 -5628 32068 -5622
rect 31140 -5640 41522 -5628
rect 41616 -5640 43872 -5626
rect 31140 -5660 43872 -5640
rect 28544 -6560 43872 -5660
rect 28544 -7800 32068 -6560
rect 28544 -8286 31344 -7800
rect 31754 -8286 32068 -7800
rect 28544 -12892 32068 -8286
rect 41440 -10236 43872 -6560
rect 54352 -9970 58052 -5034
rect 54352 -10146 57096 -9970
rect 41440 -10388 44696 -10236
rect 46574 -10388 50478 -10364
rect 41440 -10542 50478 -10388
rect 41428 -10876 50478 -10542
rect 41428 -10886 44696 -10876
rect 28544 -13518 31994 -12892
rect 28544 -18022 32100 -13518
rect 28544 -18552 31458 -18022
rect 31864 -18552 32100 -18022
rect 28544 -19844 32100 -18552
rect 41428 -15668 44134 -10886
rect 56708 -13184 57096 -10146
rect 56708 -13414 56844 -13184
rect 41428 -16182 50476 -15668
rect 41428 -19844 44134 -16182
rect 56708 -16460 57096 -13414
rect 28544 -20640 44134 -19844
rect 31174 -20776 44134 -20640
rect 41428 -20854 44134 -20776
rect 54374 -16476 57096 -16460
rect 54374 -21516 57924 -16476
rect 54386 -21540 57924 -21516
rect 31220 -27426 58000 -26394
rect 31244 -29004 58000 -27426
rect 31244 -30500 40896 -29004
rect 44220 -30500 58000 -29004
rect 31244 -30940 58000 -30500
<< viali >>
rect 28840 1906 30322 3482
rect 31344 -8286 31754 -7800
rect 31458 -18552 31864 -18022
rect 56844 -13414 57096 -13184
rect 40896 -30500 44220 -29004
<< metal1 >>
rect 28534 3482 30770 3764
rect 28534 1906 28840 3482
rect 30322 1906 30770 3482
rect 28534 1718 30770 1906
rect 28606 -2464 30536 -2376
rect 28606 -2788 30052 -2464
rect 30392 -2788 30536 -2464
rect 28606 -2878 30536 -2788
rect 31528 -2378 32032 -236
rect 32092 -1110 32216 -532
rect 32092 -1258 32094 -1110
rect 32214 -1258 32216 -1110
rect 32092 -1922 32216 -1258
rect 31528 -2886 31610 -2378
rect 31932 -2886 32032 -2378
rect 31336 -4018 31460 -3378
rect 31336 -4166 31338 -4018
rect 31458 -4166 31460 -4018
rect 31336 -4768 31460 -4166
rect 31528 -4960 32032 -2886
rect 32278 -2402 32782 -242
rect 32278 -2910 32348 -2402
rect 32670 -2910 32782 -2402
rect 32278 -4966 32782 -2910
rect 33048 -2384 33552 -248
rect 33612 -1062 33736 -552
rect 33612 -1210 33614 -1062
rect 33734 -1210 33736 -1062
rect 33612 -1942 33736 -1210
rect 33048 -2892 33122 -2384
rect 33444 -2892 33552 -2384
rect 32854 -3974 32978 -3368
rect 32854 -4122 32858 -3974
rect 32854 -4758 32978 -4122
rect 33048 -4972 33552 -2892
rect 33818 -2384 34322 -244
rect 33818 -2892 33912 -2384
rect 34234 -2892 34322 -2384
rect 33818 -4968 34322 -2892
rect 34558 -2372 35062 -244
rect 35120 -1102 35244 -552
rect 35120 -1250 35124 -1102
rect 35120 -1942 35244 -1250
rect 34558 -2880 34638 -2372
rect 34960 -2880 35062 -2372
rect 34372 -3958 34496 -3366
rect 34372 -4106 34376 -3958
rect 34372 -4756 34496 -4106
rect 34558 -4968 35062 -2880
rect 35312 -2350 35816 -248
rect 35312 -2858 35384 -2350
rect 35706 -2858 35816 -2350
rect 35312 -4972 35816 -2858
rect 36076 -2372 36580 -244
rect 36646 -1124 36770 -538
rect 36766 -1272 36770 -1124
rect 36646 -1928 36770 -1272
rect 36076 -2880 36146 -2372
rect 36468 -2880 36580 -2372
rect 35880 -3982 36004 -3372
rect 35880 -4130 35882 -3982
rect 36002 -4130 36004 -3982
rect 35880 -4762 36004 -4130
rect 36076 -4968 36580 -2880
rect 36852 -2344 37356 -248
rect 36852 -2852 36930 -2344
rect 37252 -2852 37356 -2344
rect 36852 -4972 37356 -2852
rect 37602 -2378 38106 -248
rect 38154 -1146 38278 -546
rect 38154 -1294 38158 -1146
rect 38154 -1936 38278 -1294
rect 37602 -2886 37708 -2378
rect 38030 -2886 38106 -2378
rect 37402 -4000 37526 -3352
rect 37402 -4148 37404 -4000
rect 37524 -4148 37526 -4000
rect 37402 -4742 37526 -4148
rect 37602 -4972 38106 -2886
rect 38350 -2362 38854 -248
rect 38350 -2870 38430 -2362
rect 38752 -2870 38854 -2362
rect 38350 -4972 38854 -2870
rect 39118 -2378 39622 -244
rect 39674 -1110 39798 -516
rect 39674 -1258 39678 -1110
rect 39674 -1906 39798 -1258
rect 39118 -2886 39186 -2378
rect 39508 -2886 39622 -2378
rect 38916 -3994 39040 -3362
rect 38916 -4142 38918 -3994
rect 39038 -4142 39040 -3994
rect 38916 -4752 39040 -4142
rect 39118 -4968 39622 -2886
rect 39862 -2378 40366 -248
rect 39862 -2886 39942 -2378
rect 40264 -2886 40366 -2378
rect 39862 -4972 40366 -2886
rect 40632 -2368 41136 -242
rect 41196 -1100 41320 -520
rect 41196 -1248 41200 -1100
rect 41196 -1910 41320 -1248
rect 40632 -2876 40710 -2368
rect 41032 -2876 41136 -2368
rect 40434 -4002 40558 -3394
rect 40434 -4150 40436 -4002
rect 40556 -4150 40558 -4002
rect 40434 -4784 40558 -4150
rect 40632 -4966 41136 -2876
rect 41380 -2362 41884 -252
rect 41380 -2870 41478 -2362
rect 41800 -2870 41884 -2362
rect 41380 -4976 41884 -2870
rect 42138 -2378 42642 -244
rect 42710 -1062 42834 -538
rect 42710 -1210 42712 -1062
rect 42832 -1210 42834 -1062
rect 42710 -1928 42834 -1210
rect 42138 -2886 42228 -2378
rect 42550 -2886 42642 -2378
rect 41952 -3996 42076 -3398
rect 41952 -4144 41956 -3996
rect 41952 -4788 42076 -4144
rect 42138 -4968 42642 -2886
rect 42908 -2368 43412 -248
rect 42908 -2876 43000 -2368
rect 43322 -2876 43412 -2368
rect 42908 -4972 43412 -2876
rect 43672 -2344 44176 -242
rect 44224 -1096 44348 -538
rect 44224 -1244 44228 -1096
rect 44224 -1928 44348 -1244
rect 43672 -2852 43768 -2344
rect 44090 -2852 44176 -2344
rect 43470 -3976 43594 -3388
rect 43470 -4124 43474 -3976
rect 43470 -4778 43594 -4124
rect 43672 -4966 44176 -2852
rect 44420 -2338 44924 -248
rect 44420 -2846 44496 -2338
rect 44818 -2846 44924 -2338
rect 44420 -4972 44924 -2846
rect 45174 -2362 45678 -244
rect 45738 -1082 45862 -546
rect 45738 -1230 45740 -1082
rect 45860 -1230 45862 -1082
rect 45738 -1936 45862 -1230
rect 45174 -2870 45262 -2362
rect 45584 -2870 45678 -2362
rect 44986 -3974 45110 -3358
rect 44986 -4122 44988 -3974
rect 45108 -4122 45110 -3974
rect 44986 -4748 45110 -4122
rect 45174 -4968 45678 -2870
rect 45936 -2368 46440 -242
rect 45936 -2876 46014 -2368
rect 46336 -2876 46440 -2368
rect 45936 -4966 46440 -2876
rect 46686 -2368 47190 -242
rect 47256 -1102 47380 -546
rect 47256 -1250 47258 -1102
rect 47378 -1250 47380 -1102
rect 47256 -1936 47380 -1250
rect 46686 -2876 46780 -2368
rect 47102 -2876 47190 -2368
rect 46494 -3966 46618 -3352
rect 46494 -4114 46496 -3966
rect 46616 -4114 46618 -3966
rect 46494 -4742 46618 -4114
rect 46686 -4966 47190 -2876
rect 47454 -2408 47958 -244
rect 47454 -2916 47526 -2408
rect 47848 -2916 47958 -2408
rect 47454 -4968 47958 -2916
rect 48214 -2418 48718 -242
rect 48770 -1104 48894 -538
rect 48770 -1252 48772 -1104
rect 48892 -1252 48894 -1104
rect 48770 -1928 48894 -1252
rect 48214 -2926 48298 -2418
rect 48620 -2926 48718 -2418
rect 48024 -3962 48148 -3378
rect 48144 -4110 48148 -3962
rect 48024 -4768 48148 -4110
rect 48214 -4966 48718 -2926
rect 48972 -2362 49476 -242
rect 48972 -2870 49072 -2362
rect 49394 -2870 49476 -2362
rect 48972 -4966 49476 -2870
rect 49722 -2368 50226 -248
rect 50284 -1102 50408 -526
rect 50404 -1250 50408 -1102
rect 50284 -1916 50408 -1250
rect 49722 -2876 49804 -2368
rect 50126 -2876 50226 -2368
rect 49532 -3974 49656 -3384
rect 49532 -4122 49534 -3974
rect 49654 -4122 49656 -3974
rect 49532 -4774 49656 -4122
rect 49722 -4972 50226 -2876
rect 50486 -2344 50990 -244
rect 50486 -2852 50578 -2344
rect 50900 -2852 50990 -2344
rect 50486 -4968 50990 -2852
rect 51232 -2332 51736 -238
rect 51804 -1112 51928 -546
rect 51804 -1260 51806 -1112
rect 51926 -1260 51928 -1112
rect 51804 -1936 51928 -1260
rect 51232 -2840 51328 -2332
rect 51650 -2840 51736 -2332
rect 51050 -3964 51174 -3390
rect 51050 -4112 51052 -3964
rect 51172 -4112 51174 -3964
rect 51050 -4780 51174 -4112
rect 51232 -4962 51736 -2840
rect 52008 -2364 52512 -244
rect 52008 -2872 52092 -2364
rect 52414 -2872 52512 -2364
rect 52008 -4968 52512 -2872
rect 52744 -2352 53248 -242
rect 53308 -1116 53432 -548
rect 53308 -1264 53310 -1116
rect 53430 -1264 53432 -1116
rect 53308 -1938 53432 -1264
rect 52744 -2860 52848 -2352
rect 53170 -2860 53248 -2352
rect 52564 -3982 52688 -3378
rect 52684 -4130 52688 -3982
rect 52564 -4768 52688 -4130
rect 52744 -4966 53248 -2860
rect 53510 -2366 54014 -244
rect 53510 -2874 53598 -2366
rect 53920 -2874 54014 -2366
rect 53510 -4968 54014 -2874
rect 54280 -2332 54784 -238
rect 54838 -1104 54962 -558
rect 54838 -1252 54842 -1104
rect 54838 -1948 54962 -1252
rect 54280 -2384 54806 -2332
rect 54280 -2892 54378 -2384
rect 54700 -2538 54806 -2384
rect 55032 -2382 55536 -238
rect 54700 -2892 54802 -2538
rect 54280 -2914 54802 -2892
rect 55032 -2890 55126 -2382
rect 55448 -2890 55536 -2382
rect 54084 -3960 54208 -3378
rect 54084 -4108 54088 -3960
rect 54084 -4768 54208 -4108
rect 54280 -4962 54784 -2914
rect 55032 -4962 55536 -2890
rect 55778 -2392 56282 -246
rect 56342 -1080 56466 -546
rect 56462 -1228 56466 -1080
rect 56342 -1936 56466 -1228
rect 55778 -2900 55882 -2392
rect 56204 -2900 56282 -2392
rect 55598 -3966 55722 -3388
rect 55598 -4114 55600 -3966
rect 55720 -4114 55722 -3966
rect 55598 -4778 55722 -4114
rect 55778 -4970 56282 -2900
rect 56546 -2382 57050 -242
rect 56546 -2890 56626 -2382
rect 56948 -2890 57050 -2382
rect 56546 -4966 57050 -2890
rect 57292 -2372 57796 -246
rect 57860 -1070 57984 -532
rect 57860 -1218 57864 -1070
rect 57860 -1922 57984 -1218
rect 57292 -2880 57376 -2372
rect 57698 -2880 57796 -2372
rect 57110 -3960 57234 -3394
rect 57110 -4108 57112 -3960
rect 57232 -4108 57234 -3960
rect 57110 -4784 57234 -4108
rect 57292 -4970 57796 -2880
rect 31242 -7784 31870 -7354
rect 31242 -8314 31344 -7784
rect 31750 -7800 31870 -7784
rect 31754 -8286 31870 -7800
rect 31750 -8314 31870 -8286
rect 31242 -8658 31870 -8314
rect 32438 -9412 34858 -6624
rect 35040 -7892 35336 -7160
rect 35040 -8280 35088 -7892
rect 35296 -8280 35336 -7892
rect 35040 -8930 35336 -8280
rect 32438 -9962 33246 -9412
rect 34070 -9962 34858 -9412
rect 32020 -11122 32308 -10538
rect 32020 -11566 32060 -11122
rect 32302 -11566 32308 -11122
rect 32020 -12120 32308 -11566
rect 32438 -12794 34858 -9962
rect 35488 -9424 37908 -6624
rect 35488 -9974 36258 -9424
rect 37082 -9974 37908 -9424
rect 35488 -12794 37908 -9974
rect 38590 -9434 41010 -6624
rect 41212 -7836 41436 -7172
rect 41212 -8334 41238 -7836
rect 41400 -8334 41436 -7836
rect 41212 -8896 41436 -8334
rect 46892 -8158 47344 -6882
rect 46892 -8412 47014 -8158
rect 47254 -8412 47344 -8158
rect 46892 -8472 47344 -8412
rect 38590 -9984 39420 -9434
rect 40244 -9984 41010 -9434
rect 38100 -11266 38436 -10706
rect 38100 -11682 38104 -11266
rect 38434 -11682 38436 -11266
rect 38100 -12224 38436 -11682
rect 38590 -12794 41010 -9984
rect 54606 -10192 55362 -10126
rect 54606 -10352 54748 -10192
rect 55104 -10352 55362 -10192
rect 54606 -10400 55362 -10352
rect 45196 -10786 45736 -10734
rect 48370 -10940 49098 -10922
rect 48370 -11000 48708 -10940
rect 48778 -11000 49098 -10940
rect 48370 -11018 49098 -11000
rect 44214 -11168 50376 -11056
rect 44214 -11410 46884 -11168
rect 47330 -11410 50376 -11168
rect 44214 -11562 50376 -11410
rect 45218 -11598 45852 -11596
rect 45218 -11658 45482 -11598
rect 45552 -11658 45852 -11598
rect 45218 -11662 45852 -11658
rect 44208 -11826 50370 -11716
rect 44208 -12068 46894 -11826
rect 47340 -12068 50370 -11826
rect 44208 -12222 50370 -12068
rect 48278 -12258 49406 -12250
rect 48278 -12318 48738 -12258
rect 48808 -12318 49406 -12258
rect 48278 -12330 49406 -12318
rect 44202 -12520 50364 -12376
rect 44202 -12762 46894 -12520
rect 47340 -12762 50364 -12520
rect 44202 -12882 50364 -12762
rect 45140 -12916 45774 -12912
rect 45140 -12976 45430 -12916
rect 45500 -12976 45774 -12916
rect 45140 -12978 45774 -12976
rect 54494 -13108 54690 -10478
rect 55230 -11588 56640 -10478
rect 55230 -11874 55462 -11588
rect 55670 -11874 56640 -11588
rect 55230 -13108 56640 -11874
rect 56006 -13266 56334 -13176
rect 56006 -13370 56122 -13266
rect 56248 -13370 56334 -13266
rect 56006 -13470 56334 -13370
rect 56792 -13184 57154 -13120
rect 56792 -13414 56844 -13184
rect 57096 -13414 57154 -13184
rect 56792 -13518 57154 -13414
rect 48444 -13572 49172 -13552
rect 32516 -16430 34936 -13614
rect 35582 -13618 36458 -13614
rect 37194 -13618 38002 -13614
rect 35096 -14802 35432 -14226
rect 35096 -15190 35120 -14802
rect 35396 -15190 35432 -14802
rect 35096 -15744 35432 -15190
rect 32516 -16980 33348 -16430
rect 34172 -16980 34936 -16430
rect 31358 -18022 31944 -17792
rect 31358 -18552 31458 -18022
rect 31864 -18552 31944 -18022
rect 31358 -18884 31944 -18552
rect 32026 -18044 32424 -17526
rect 32026 -18724 32084 -18044
rect 32366 -18724 32424 -18044
rect 32026 -19166 32424 -18724
rect 32516 -19784 34936 -16980
rect 35582 -16436 38002 -13618
rect 35582 -16986 36396 -16436
rect 37220 -16986 38002 -16436
rect 35582 -19784 38002 -16986
rect 38650 -16430 41070 -13610
rect 48444 -13632 48744 -13572
rect 48814 -13632 49172 -13572
rect 48444 -13648 49172 -13632
rect 54496 -13640 54690 -13556
rect 55230 -13640 56642 -13556
rect 44208 -13808 50370 -13676
rect 44208 -14050 46866 -13808
rect 47312 -14050 50370 -13808
rect 44208 -14182 50370 -14050
rect 41192 -14750 41528 -14202
rect 45116 -14232 45750 -14228
rect 45116 -14292 45418 -14232
rect 45488 -14292 45750 -14232
rect 45116 -14294 45750 -14292
rect 41192 -15138 41228 -14750
rect 41504 -15138 41528 -14750
rect 44208 -14466 50370 -14340
rect 44208 -14708 46888 -14466
rect 47334 -14708 50370 -14466
rect 44208 -14846 50370 -14708
rect 54496 -14708 56642 -13640
rect 48456 -14886 49172 -14878
rect 48456 -14946 48742 -14886
rect 48812 -14946 49172 -14886
rect 48456 -14958 49172 -14946
rect 41192 -15720 41528 -15138
rect 44214 -15120 50376 -14988
rect 44214 -15362 46894 -15120
rect 47340 -15362 50376 -15120
rect 44214 -15494 50376 -15362
rect 54496 -14994 55456 -14708
rect 55664 -14994 56642 -14708
rect 45094 -15544 45728 -15542
rect 45094 -15604 45384 -15544
rect 45454 -15604 45728 -15544
rect 45094 -15608 45728 -15604
rect 54496 -16024 56642 -14994
rect 54496 -16186 55034 -16024
rect 55194 -16186 56642 -16024
rect 38650 -16980 39402 -16430
rect 40226 -16980 41070 -16430
rect 54642 -16320 55034 -16306
rect 54642 -16424 54878 -16320
rect 55004 -16424 55034 -16320
rect 54642 -16438 55034 -16424
rect 38148 -18058 38490 -17532
rect 38148 -18478 38190 -18058
rect 38446 -18478 38490 -18058
rect 38148 -19212 38490 -18478
rect 38650 -19780 41070 -16980
rect 55420 -17236 55736 -17190
rect 55420 -17458 55462 -17236
rect 55682 -17458 55736 -17236
rect 55420 -18096 55736 -17458
rect 29038 -23756 30344 -23640
rect 29038 -24126 29836 -23756
rect 30200 -24126 30344 -23756
rect 29038 -24224 30344 -24126
rect 31476 -23676 31980 -21598
rect 32048 -22512 32172 -21798
rect 32048 -22660 32050 -22512
rect 32170 -22660 32172 -22512
rect 32048 -23188 32172 -22660
rect 31476 -24184 31568 -23676
rect 31890 -24184 31980 -23676
rect 31296 -25332 31420 -24658
rect 31416 -25480 31420 -25332
rect 31296 -26048 31420 -25480
rect 31476 -26328 31980 -24184
rect 32234 -23676 32738 -21598
rect 32234 -24184 32322 -23676
rect 32644 -24184 32738 -23676
rect 32234 -26328 32738 -24184
rect 33002 -23652 33506 -21596
rect 33564 -22506 33688 -21798
rect 33564 -22654 33566 -22506
rect 33686 -22654 33688 -22506
rect 33564 -23188 33688 -22654
rect 33002 -24160 33070 -23652
rect 33392 -24160 33506 -23652
rect 32808 -25340 32932 -24640
rect 32928 -25488 32932 -25340
rect 32808 -26030 32932 -25488
rect 33002 -26326 33506 -24160
rect 33746 -23686 34250 -21596
rect 33746 -24194 33842 -23686
rect 34164 -24194 34250 -23686
rect 33746 -26326 34250 -24194
rect 34500 -23672 35004 -21598
rect 35072 -22466 35196 -21798
rect 35072 -22614 35074 -22466
rect 35194 -22614 35196 -22466
rect 35072 -23188 35196 -22614
rect 34500 -24180 34580 -23672
rect 34902 -24180 35004 -23672
rect 34322 -25372 34446 -24642
rect 34442 -25520 34446 -25372
rect 34322 -26032 34446 -25520
rect 34500 -26328 35004 -24180
rect 35264 -23676 35768 -21596
rect 35264 -24184 35352 -23676
rect 35674 -24184 35768 -23676
rect 35264 -26326 35768 -24184
rect 36030 -23652 36534 -21602
rect 36596 -22488 36720 -21814
rect 36596 -22636 36600 -22488
rect 36596 -23204 36720 -22636
rect 36030 -24160 36112 -23652
rect 36434 -24160 36534 -23652
rect 35838 -25372 35962 -24666
rect 35838 -25520 35840 -25372
rect 35960 -25520 35962 -25372
rect 35838 -26056 35962 -25520
rect 36030 -26332 36534 -24160
rect 36760 -23652 37264 -21602
rect 36760 -24160 36880 -23652
rect 37202 -24160 37264 -23652
rect 36760 -26332 37264 -24160
rect 37542 -23664 38046 -21598
rect 38100 -22484 38224 -21840
rect 38220 -22632 38224 -22484
rect 38100 -23230 38224 -22632
rect 37542 -24172 37620 -23664
rect 37942 -24172 38046 -23664
rect 37354 -25374 37478 -24658
rect 37474 -25522 37478 -25374
rect 37354 -26048 37478 -25522
rect 37542 -26328 38046 -24172
rect 38282 -23672 38786 -21600
rect 38282 -24180 38374 -23672
rect 38696 -24180 38786 -23672
rect 38282 -26330 38786 -24180
rect 39058 -23666 39562 -21596
rect 39628 -22462 39752 -21798
rect 39628 -22610 39630 -22462
rect 39750 -22610 39752 -22462
rect 39628 -23188 39752 -22610
rect 39058 -24174 39152 -23666
rect 39474 -24174 39562 -23666
rect 38876 -25358 39000 -24656
rect 38996 -25506 39000 -25358
rect 38876 -26046 39000 -25506
rect 39058 -26326 39562 -24174
rect 39818 -23660 40322 -21596
rect 39818 -24168 39898 -23660
rect 40220 -24168 40322 -23660
rect 39818 -26326 40322 -24168
rect 40570 -23638 41074 -21600
rect 41148 -22466 41272 -21798
rect 41268 -22614 41272 -22466
rect 41148 -23188 41272 -22614
rect 40570 -24146 40676 -23638
rect 40998 -24146 41074 -23638
rect 40390 -25388 40514 -24640
rect 40390 -25536 40392 -25388
rect 40512 -25536 40514 -25388
rect 40390 -26030 40514 -25536
rect 40570 -26330 41074 -24146
rect 41324 -23658 41828 -21600
rect 41324 -24166 41402 -23658
rect 41724 -24166 41828 -23658
rect 41324 -26330 41828 -24166
rect 42080 -23656 42584 -21596
rect 42658 -22474 42782 -21804
rect 42778 -22622 42782 -22474
rect 42658 -23194 42782 -22622
rect 42080 -24164 42186 -23656
rect 42508 -24164 42584 -23656
rect 41896 -25390 42020 -24652
rect 41896 -25538 41898 -25390
rect 42018 -25538 42020 -25390
rect 41896 -26042 42020 -25538
rect 42080 -26326 42584 -24164
rect 42842 -23664 43346 -21596
rect 42842 -24172 42938 -23664
rect 43260 -24172 43346 -23664
rect 42842 -26326 43346 -24172
rect 43606 -23672 44110 -21598
rect 44172 -22478 44296 -21808
rect 44172 -22626 44176 -22478
rect 44172 -23198 44296 -22626
rect 43606 -24180 43682 -23672
rect 44004 -24180 44110 -23672
rect 43420 -25312 43544 -24646
rect 43420 -25460 43424 -25312
rect 43420 -26036 43544 -25460
rect 43606 -26328 44110 -24180
rect 44352 -23690 44856 -21598
rect 44352 -24198 44422 -23690
rect 44744 -24198 44856 -23690
rect 44352 -26328 44856 -24198
rect 45120 -23684 45624 -21598
rect 45690 -22466 45814 -21798
rect 45690 -22614 45692 -22466
rect 45812 -22614 45814 -22466
rect 45690 -23188 45814 -22614
rect 45120 -24192 45216 -23684
rect 45538 -24192 45624 -23684
rect 44930 -25336 45054 -24634
rect 44930 -25484 44932 -25336
rect 45052 -25484 45054 -25336
rect 44930 -26024 45054 -25484
rect 45120 -26328 45624 -24192
rect 45874 -23696 46378 -21600
rect 45874 -24204 45978 -23696
rect 46300 -24204 46378 -23696
rect 45874 -26330 46378 -24204
rect 46634 -23710 47138 -21600
rect 47198 -22482 47322 -21814
rect 47318 -22630 47322 -22482
rect 47198 -23204 47322 -22630
rect 46634 -24218 46722 -23710
rect 47044 -24218 47138 -23710
rect 46450 -25372 46574 -24642
rect 46570 -25520 46574 -25372
rect 46450 -26032 46574 -25520
rect 46634 -26330 47138 -24218
rect 47388 -23712 47892 -21598
rect 47388 -24220 47496 -23712
rect 47818 -24220 47892 -23712
rect 47388 -26328 47892 -24220
rect 48154 -23676 48658 -21598
rect 48716 -22462 48840 -21794
rect 48716 -22610 48720 -22462
rect 48716 -23184 48840 -22610
rect 48154 -24184 48232 -23676
rect 48554 -24184 48658 -23676
rect 47964 -25368 48088 -24652
rect 47964 -25516 47966 -25368
rect 48086 -25516 48088 -25368
rect 47964 -26042 48088 -25516
rect 48154 -26328 48658 -24184
rect 48924 -23678 49428 -21602
rect 48924 -24186 49026 -23678
rect 49348 -24186 49428 -23678
rect 48924 -26326 49428 -24186
rect 49670 -23674 50174 -21606
rect 50242 -22470 50366 -21804
rect 50242 -22618 50246 -22470
rect 50242 -23194 50366 -22618
rect 49670 -24182 49754 -23674
rect 50076 -24182 50174 -23674
rect 49476 -25350 49600 -24658
rect 49476 -25498 49480 -25350
rect 49476 -26048 49600 -25498
rect 49670 -26330 50174 -24182
rect 50424 -23666 50928 -21610
rect 50424 -24174 50502 -23666
rect 50824 -24174 50928 -23666
rect 50424 -26334 50928 -24174
rect 51182 -23658 51686 -21610
rect 51756 -22478 51880 -21808
rect 51756 -22626 51758 -22478
rect 51878 -22626 51880 -22478
rect 51756 -23198 51880 -22626
rect 51182 -24166 51268 -23658
rect 51590 -24166 51686 -23658
rect 51002 -25338 51126 -24650
rect 51002 -25486 51004 -25338
rect 51124 -25486 51126 -25338
rect 51002 -26040 51126 -25486
rect 51182 -26334 51686 -24166
rect 51942 -23660 52446 -21604
rect 51942 -24168 52038 -23660
rect 52360 -24168 52446 -23660
rect 51942 -26328 52446 -24168
rect 52692 -23640 53196 -21604
rect 53276 -22496 53400 -21810
rect 53276 -22644 53278 -22496
rect 53398 -22644 53400 -22496
rect 53276 -23200 53400 -22644
rect 52692 -24148 52776 -23640
rect 53098 -24148 53196 -23640
rect 52510 -25336 52634 -24662
rect 52510 -25484 52512 -25336
rect 52632 -25484 52634 -25336
rect 52510 -26052 52634 -25484
rect 52692 -26328 53196 -24148
rect 53458 -23660 53962 -21606
rect 53458 -24168 53536 -23660
rect 53858 -24168 53962 -23660
rect 53458 -26330 53962 -24168
rect 54234 -23686 54738 -21608
rect 54784 -22510 54908 -21788
rect 54784 -22658 54786 -22510
rect 54906 -22658 54908 -22510
rect 54784 -23178 54908 -22658
rect 54234 -24194 54324 -23686
rect 54646 -24194 54738 -23686
rect 54030 -25348 54154 -24646
rect 54030 -25496 54034 -25348
rect 54030 -26036 54154 -25496
rect 54234 -26332 54738 -24194
rect 54970 -23674 55474 -21604
rect 54970 -24182 55060 -23674
rect 55382 -24182 55474 -23674
rect 54970 -26328 55474 -24182
rect 55722 -23660 56226 -21602
rect 56302 -22488 56426 -21816
rect 56302 -22636 56304 -22488
rect 56424 -22636 56426 -22488
rect 56302 -23206 56426 -22636
rect 55722 -24168 55816 -23660
rect 56138 -24168 56226 -23660
rect 55548 -25350 55672 -24650
rect 55668 -25498 55672 -25350
rect 55548 -26040 55672 -25498
rect 55722 -26326 56226 -24168
rect 56482 -23682 56986 -21604
rect 56482 -24190 56564 -23682
rect 56886 -24190 56986 -23682
rect 56482 -26328 56986 -24190
rect 57238 -23704 57742 -21604
rect 57812 -22502 57936 -21824
rect 57932 -22650 57936 -22502
rect 57812 -23214 57936 -22650
rect 57238 -24212 57316 -23704
rect 57638 -24212 57742 -23704
rect 57062 -25366 57186 -24640
rect 57062 -25514 57066 -25366
rect 57062 -26030 57186 -25514
rect 57238 -26328 57742 -24212
rect 39994 -29004 44888 -28524
rect 39994 -30500 40896 -29004
rect 44220 -30500 44888 -29004
rect 39994 -31036 44888 -30500
<< via1 >>
rect 28840 1906 30322 3482
rect 30052 -2788 30392 -2464
rect 32094 -1258 32214 -1110
rect 31610 -2886 31932 -2378
rect 31338 -4166 31458 -4018
rect 32348 -2910 32670 -2402
rect 33614 -1210 33734 -1062
rect 33122 -2892 33444 -2384
rect 32858 -4122 32978 -3974
rect 33912 -2892 34234 -2384
rect 35124 -1250 35244 -1102
rect 34638 -2880 34960 -2372
rect 34376 -4106 34496 -3958
rect 35384 -2858 35706 -2350
rect 36646 -1272 36766 -1124
rect 36146 -2880 36468 -2372
rect 35882 -4130 36002 -3982
rect 36930 -2852 37252 -2344
rect 38158 -1294 38278 -1146
rect 37708 -2886 38030 -2378
rect 37404 -4148 37524 -4000
rect 38430 -2870 38752 -2362
rect 39678 -1258 39798 -1110
rect 39186 -2886 39508 -2378
rect 38918 -4142 39038 -3994
rect 39942 -2886 40264 -2378
rect 41200 -1248 41320 -1100
rect 40710 -2876 41032 -2368
rect 40436 -4150 40556 -4002
rect 41478 -2870 41800 -2362
rect 42712 -1210 42832 -1062
rect 42228 -2886 42550 -2378
rect 41956 -4144 42076 -3996
rect 43000 -2876 43322 -2368
rect 44228 -1244 44348 -1096
rect 43768 -2852 44090 -2344
rect 43474 -4124 43594 -3976
rect 44496 -2846 44818 -2338
rect 45740 -1230 45860 -1082
rect 45262 -2870 45584 -2362
rect 44988 -4122 45108 -3974
rect 46014 -2876 46336 -2368
rect 47258 -1250 47378 -1102
rect 46780 -2876 47102 -2368
rect 46496 -4114 46616 -3966
rect 47526 -2916 47848 -2408
rect 48772 -1252 48892 -1104
rect 48298 -2926 48620 -2418
rect 48024 -4110 48144 -3962
rect 49072 -2870 49394 -2362
rect 50284 -1250 50404 -1102
rect 49804 -2876 50126 -2368
rect 49534 -4122 49654 -3974
rect 50578 -2852 50900 -2344
rect 51806 -1260 51926 -1112
rect 51328 -2840 51650 -2332
rect 51052 -4112 51172 -3964
rect 52092 -2872 52414 -2364
rect 53310 -1264 53430 -1116
rect 52848 -2860 53170 -2352
rect 52564 -4130 52684 -3982
rect 53598 -2874 53920 -2366
rect 54842 -1252 54962 -1104
rect 54378 -2892 54700 -2384
rect 55126 -2890 55448 -2382
rect 54088 -4108 54208 -3960
rect 56342 -1228 56462 -1080
rect 55882 -2900 56204 -2392
rect 55600 -4114 55720 -3966
rect 56626 -2890 56948 -2382
rect 57864 -1218 57984 -1070
rect 57376 -2880 57698 -2372
rect 57112 -4108 57232 -3960
rect 31344 -7800 31750 -7784
rect 31344 -8286 31750 -7800
rect 31344 -8314 31750 -8286
rect 35088 -8280 35296 -7892
rect 33246 -9962 34070 -9412
rect 32060 -11566 32302 -11122
rect 36258 -9974 37082 -9424
rect 41238 -8334 41400 -7836
rect 47014 -8412 47254 -8158
rect 39420 -9984 40244 -9434
rect 38104 -11682 38434 -11266
rect 54748 -10352 55104 -10192
rect 48708 -11000 48778 -10940
rect 46884 -11410 47330 -11168
rect 45482 -11658 45552 -11598
rect 46894 -12068 47340 -11826
rect 48738 -12318 48808 -12258
rect 46894 -12762 47340 -12520
rect 45430 -12976 45500 -12916
rect 55462 -11874 55670 -11588
rect 56122 -13370 56248 -13266
rect 56844 -13414 57096 -13184
rect 35120 -15190 35396 -14802
rect 33348 -16980 34172 -16430
rect 31458 -18552 31864 -18022
rect 32084 -18724 32366 -18044
rect 36396 -16986 37220 -16436
rect 48744 -13632 48814 -13572
rect 46866 -14050 47312 -13808
rect 45418 -14292 45488 -14232
rect 41228 -15138 41504 -14750
rect 46888 -14708 47334 -14466
rect 48742 -14946 48812 -14886
rect 46894 -15362 47340 -15120
rect 55456 -14994 55664 -14708
rect 45384 -15604 45454 -15544
rect 39402 -16980 40226 -16430
rect 54878 -16424 55004 -16320
rect 38190 -18478 38446 -18058
rect 55462 -17458 55682 -17236
rect 29836 -24126 30200 -23756
rect 32050 -22660 32170 -22512
rect 31568 -24184 31890 -23676
rect 31296 -25480 31416 -25332
rect 32322 -24184 32644 -23676
rect 33566 -22654 33686 -22506
rect 33070 -24160 33392 -23652
rect 32808 -25488 32928 -25340
rect 33842 -24194 34164 -23686
rect 35074 -22614 35194 -22466
rect 34580 -24180 34902 -23672
rect 34322 -25520 34442 -25372
rect 35352 -24184 35674 -23676
rect 36600 -22636 36720 -22488
rect 36112 -24160 36434 -23652
rect 35840 -25520 35960 -25372
rect 36880 -24160 37202 -23652
rect 38100 -22632 38220 -22484
rect 37620 -24172 37942 -23664
rect 37354 -25522 37474 -25374
rect 38374 -24180 38696 -23672
rect 39630 -22610 39750 -22462
rect 39152 -24174 39474 -23666
rect 38876 -25506 38996 -25358
rect 39898 -24168 40220 -23660
rect 41148 -22614 41268 -22466
rect 40676 -24146 40998 -23638
rect 40392 -25536 40512 -25388
rect 41402 -24166 41724 -23658
rect 42658 -22622 42778 -22474
rect 42186 -24164 42508 -23656
rect 41898 -25538 42018 -25390
rect 42938 -24172 43260 -23664
rect 44176 -22626 44296 -22478
rect 43682 -24180 44004 -23672
rect 43424 -25460 43544 -25312
rect 44422 -24198 44744 -23690
rect 45692 -22614 45812 -22466
rect 45216 -24192 45538 -23684
rect 44932 -25484 45052 -25336
rect 45978 -24204 46300 -23696
rect 47198 -22630 47318 -22482
rect 46722 -24218 47044 -23710
rect 46450 -25520 46570 -25372
rect 47496 -24220 47818 -23712
rect 48720 -22610 48840 -22462
rect 48232 -24184 48554 -23676
rect 47966 -25516 48086 -25368
rect 49026 -24186 49348 -23678
rect 50246 -22618 50366 -22470
rect 49754 -24182 50076 -23674
rect 49480 -25498 49600 -25350
rect 50502 -24174 50824 -23666
rect 51758 -22626 51878 -22478
rect 51268 -24166 51590 -23658
rect 51004 -25486 51124 -25338
rect 52038 -24168 52360 -23660
rect 53278 -22644 53398 -22496
rect 52776 -24148 53098 -23640
rect 52512 -25484 52632 -25336
rect 53536 -24168 53858 -23660
rect 54786 -22658 54906 -22510
rect 54324 -24194 54646 -23686
rect 54034 -25496 54154 -25348
rect 55060 -24182 55382 -23674
rect 56304 -22636 56424 -22488
rect 55816 -24168 56138 -23660
rect 55548 -25498 55668 -25350
rect 56564 -24190 56886 -23682
rect 57812 -22650 57932 -22502
rect 57316 -24212 57638 -23704
rect 57066 -25514 57186 -25366
rect 40896 -30500 44220 -29004
<< metal2 >>
rect 28544 3482 58134 4684
rect 28544 1906 28840 3482
rect 30322 1906 58134 3482
rect 28544 1668 58134 1906
rect 42868 -462 44424 -444
rect 31220 -474 57948 -462
rect 31220 -908 58180 -474
rect 31220 -1062 54600 -908
rect 31220 -1110 33614 -1062
rect 31220 -1258 32094 -1110
rect 32214 -1210 33614 -1110
rect 33734 -1100 42712 -1062
rect 33734 -1102 41200 -1100
rect 33734 -1210 35124 -1102
rect 32214 -1250 35124 -1210
rect 35244 -1110 41200 -1102
rect 35244 -1124 39678 -1110
rect 35244 -1250 36646 -1124
rect 32214 -1258 36646 -1250
rect 31220 -1272 36646 -1258
rect 36766 -1146 39678 -1124
rect 36766 -1272 38158 -1146
rect 31220 -1294 38158 -1272
rect 38278 -1258 39678 -1146
rect 39798 -1248 41200 -1110
rect 41320 -1210 42712 -1100
rect 42832 -1082 54600 -1062
rect 42832 -1096 45740 -1082
rect 42832 -1210 44228 -1096
rect 41320 -1244 44228 -1210
rect 44348 -1230 45740 -1096
rect 45860 -1102 54600 -1082
rect 45860 -1230 47258 -1102
rect 44348 -1244 47258 -1230
rect 41320 -1248 47258 -1244
rect 39798 -1250 47258 -1248
rect 47378 -1104 50284 -1102
rect 47378 -1250 48772 -1104
rect 39798 -1252 48772 -1250
rect 48892 -1250 50284 -1104
rect 50404 -1112 54600 -1102
rect 55168 -1070 58180 -908
rect 55168 -1080 57864 -1070
rect 50404 -1250 51806 -1112
rect 48892 -1252 51806 -1250
rect 39798 -1258 51806 -1252
rect 38278 -1260 51806 -1258
rect 51926 -1116 54600 -1112
rect 51926 -1260 53310 -1116
rect 38278 -1264 53310 -1260
rect 53430 -1264 54600 -1116
rect 55168 -1228 56342 -1080
rect 56462 -1218 57864 -1080
rect 57984 -1218 58180 -1070
rect 56462 -1228 58180 -1218
rect 55168 -1236 58180 -1228
rect 38278 -1294 54600 -1264
rect 31220 -1742 54600 -1294
rect 55168 -1742 58150 -1236
rect 31220 -1962 54646 -1742
rect 31220 -1974 42898 -1962
rect 43902 -1974 54646 -1962
rect 54774 -1974 58150 -1742
rect 28240 -2210 30222 -2060
rect 30674 -2210 31272 -2176
rect 28240 -2222 31272 -2210
rect 54536 -2222 54960 -2210
rect 28240 -2266 58104 -2222
rect 28240 -3024 28412 -2266
rect 29010 -2332 58104 -2266
rect 29010 -2338 51328 -2332
rect 29010 -2344 44496 -2338
rect 29010 -2350 36930 -2344
rect 29010 -2372 35384 -2350
rect 29010 -2378 34638 -2372
rect 29010 -2464 31610 -2378
rect 29010 -2788 30052 -2464
rect 30392 -2788 31610 -2464
rect 29010 -2886 31610 -2788
rect 31932 -2384 34638 -2378
rect 31932 -2402 33122 -2384
rect 31932 -2886 32348 -2402
rect 29010 -2910 32348 -2886
rect 32670 -2892 33122 -2402
rect 33444 -2892 33912 -2384
rect 34234 -2880 34638 -2384
rect 34960 -2858 35384 -2372
rect 35706 -2372 36930 -2350
rect 35706 -2858 36146 -2372
rect 34960 -2880 36146 -2858
rect 36468 -2852 36930 -2372
rect 37252 -2362 43768 -2344
rect 37252 -2378 38430 -2362
rect 37252 -2852 37708 -2378
rect 36468 -2880 37708 -2852
rect 34234 -2886 37708 -2880
rect 38030 -2870 38430 -2378
rect 38752 -2368 41478 -2362
rect 38752 -2378 40710 -2368
rect 38752 -2870 39186 -2378
rect 38030 -2886 39186 -2870
rect 39508 -2886 39942 -2378
rect 40264 -2876 40710 -2378
rect 41032 -2870 41478 -2368
rect 41800 -2368 43768 -2362
rect 41800 -2378 43000 -2368
rect 41800 -2870 42228 -2378
rect 41032 -2876 42228 -2870
rect 40264 -2886 42228 -2876
rect 42550 -2876 43000 -2378
rect 43322 -2852 43768 -2368
rect 44090 -2846 44496 -2344
rect 44818 -2344 51328 -2338
rect 44818 -2362 50578 -2344
rect 44818 -2846 45262 -2362
rect 44090 -2852 45262 -2846
rect 43322 -2870 45262 -2852
rect 45584 -2368 49072 -2362
rect 45584 -2870 46014 -2368
rect 43322 -2876 46014 -2870
rect 46336 -2876 46780 -2368
rect 47102 -2408 49072 -2368
rect 47102 -2876 47526 -2408
rect 42550 -2886 47526 -2876
rect 34234 -2892 47526 -2886
rect 32670 -2910 47526 -2892
rect 29010 -2916 47526 -2910
rect 47848 -2418 49072 -2408
rect 47848 -2916 48298 -2418
rect 29010 -2926 48298 -2916
rect 48620 -2870 49072 -2418
rect 49394 -2368 50578 -2362
rect 49394 -2870 49804 -2368
rect 48620 -2876 49804 -2870
rect 50126 -2852 50578 -2368
rect 50900 -2840 51328 -2344
rect 51650 -2352 58104 -2332
rect 51650 -2364 52848 -2352
rect 51650 -2840 52092 -2364
rect 50900 -2852 52092 -2840
rect 50126 -2872 52092 -2852
rect 52414 -2860 52848 -2364
rect 53170 -2366 58104 -2352
rect 53170 -2860 53598 -2366
rect 52414 -2872 53598 -2860
rect 50126 -2874 53598 -2872
rect 53920 -2372 58104 -2366
rect 53920 -2382 57376 -2372
rect 53920 -2384 55126 -2382
rect 53920 -2874 54378 -2384
rect 50126 -2876 54378 -2874
rect 48620 -2892 54378 -2876
rect 54700 -2890 55126 -2384
rect 55448 -2392 56626 -2382
rect 55448 -2890 55882 -2392
rect 54700 -2892 55882 -2890
rect 48620 -2900 55882 -2892
rect 56204 -2890 56626 -2392
rect 56948 -2880 57376 -2382
rect 57698 -2880 58104 -2372
rect 56948 -2890 58104 -2880
rect 56204 -2900 58104 -2890
rect 48620 -2926 58104 -2900
rect 29010 -3024 58104 -2926
rect 28240 -3062 58104 -3024
rect 28240 -3072 30840 -3062
rect 28240 -3296 30222 -3072
rect 31182 -3078 58104 -3062
rect 31182 -3084 54646 -3078
rect 54774 -3084 58104 -3078
rect 54476 -3304 54960 -3288
rect 31128 -3958 58102 -3304
rect 31128 -3974 34376 -3958
rect 31128 -4018 32858 -3974
rect 31128 -4166 31338 -4018
rect 31458 -4122 32858 -4018
rect 32978 -4106 34376 -3974
rect 34496 -3960 58102 -3958
rect 34496 -3962 54088 -3960
rect 34496 -3966 48024 -3962
rect 34496 -3974 46496 -3966
rect 34496 -3976 44988 -3974
rect 34496 -3982 43474 -3976
rect 34496 -4106 35882 -3982
rect 32978 -4122 35882 -4106
rect 31458 -4130 35882 -4122
rect 36002 -3994 43474 -3982
rect 36002 -4000 38918 -3994
rect 36002 -4130 37404 -4000
rect 31458 -4148 37404 -4130
rect 37524 -4142 38918 -4000
rect 39038 -3996 43474 -3994
rect 39038 -4002 41956 -3996
rect 39038 -4142 40436 -4002
rect 37524 -4148 40436 -4142
rect 31458 -4150 40436 -4148
rect 40556 -4144 41956 -4002
rect 42076 -4124 43474 -3996
rect 43594 -4122 44988 -3976
rect 45108 -4114 46496 -3974
rect 46616 -4110 48024 -3966
rect 48144 -3964 54088 -3962
rect 48144 -3974 51052 -3964
rect 48144 -4110 49534 -3974
rect 46616 -4114 49534 -4110
rect 45108 -4122 49534 -4114
rect 49654 -4112 51052 -3974
rect 51172 -3982 54088 -3964
rect 51172 -4112 52564 -3982
rect 49654 -4122 52564 -4112
rect 43594 -4124 52564 -4122
rect 42076 -4130 52564 -4124
rect 52684 -4108 54088 -3982
rect 54208 -3966 57112 -3960
rect 54208 -4108 55600 -3966
rect 52684 -4114 55600 -4108
rect 55720 -4108 57112 -3966
rect 57232 -4108 58102 -3960
rect 55720 -4114 58102 -4108
rect 52684 -4130 58102 -4114
rect 42076 -4144 58102 -4130
rect 40556 -4150 58102 -4144
rect 31458 -4166 58102 -4150
rect 31128 -4812 58102 -4166
rect 31128 -4816 54646 -4812
rect 54774 -4816 56268 -4812
rect 57400 -4816 58102 -4812
rect 35344 -4822 36080 -4816
rect 47820 -5552 49596 -4816
rect 47820 -6218 60428 -5552
rect 46752 -6920 47448 -6848
rect 31094 -7784 41522 -7158
rect 31094 -8314 31344 -7784
rect 31750 -7836 41522 -7784
rect 31750 -7892 41238 -7836
rect 31750 -8280 35088 -7892
rect 35296 -8280 41238 -7892
rect 31750 -8314 41238 -8280
rect 31094 -8334 41238 -8314
rect 41400 -8334 41522 -7836
rect 46752 -7310 46932 -6920
rect 47314 -7310 47448 -6920
rect 46752 -8120 47448 -7310
rect 31094 -8938 41522 -8334
rect 46740 -8158 47448 -8120
rect 46740 -8412 47014 -8158
rect 47254 -8412 47448 -8158
rect 46740 -8636 47448 -8412
rect 41318 -9344 42274 -9318
rect 31960 -9412 42274 -9344
rect 31960 -9962 33246 -9412
rect 34070 -9424 42274 -9412
rect 34070 -9962 36258 -9424
rect 31960 -9974 36258 -9962
rect 37082 -9434 42274 -9424
rect 37082 -9974 39420 -9434
rect 31960 -9984 39420 -9974
rect 40244 -9496 42274 -9434
rect 40244 -9844 41676 -9496
rect 42114 -9844 42274 -9496
rect 40244 -9984 42274 -9844
rect 31960 -10036 42274 -9984
rect 31960 -10040 41522 -10036
rect 46752 -10164 47448 -8636
rect 46738 -10440 47448 -10164
rect 47820 -7908 58362 -6218
rect 59962 -7908 60428 -6218
rect 47820 -8666 60428 -7908
rect 31960 -10472 39908 -10454
rect 40964 -10472 41510 -10454
rect 31960 -10734 44486 -10472
rect 31960 -11122 46414 -10734
rect 31960 -11566 32060 -11122
rect 32302 -11266 46414 -11122
rect 32302 -11566 38104 -11266
rect 31960 -11682 38104 -11566
rect 38434 -11598 46414 -11266
rect 38434 -11658 45482 -11598
rect 45552 -11658 46414 -11598
rect 38434 -11682 46414 -11658
rect 31960 -12234 46414 -11682
rect 39782 -12268 46414 -12234
rect 44018 -12460 46414 -12268
rect 44634 -12916 46414 -12460
rect 44634 -12976 45430 -12916
rect 45500 -12976 46414 -12916
rect 44634 -13118 46414 -12976
rect 46738 -11168 47434 -10440
rect 47820 -10766 49596 -8666
rect 54690 -9954 55230 -9774
rect 54580 -10192 55310 -9954
rect 55426 -10074 55712 -9842
rect 54580 -10352 54748 -10192
rect 55104 -10352 55310 -10192
rect 47820 -10940 49606 -10766
rect 47820 -11000 48708 -10940
rect 48778 -11000 49606 -10940
rect 47820 -11072 49606 -11000
rect 46738 -11410 46884 -11168
rect 47330 -11410 47434 -11168
rect 46738 -11826 47434 -11410
rect 46738 -12068 46894 -11826
rect 47340 -12068 47434 -11826
rect 46738 -12520 47434 -12068
rect 46738 -12762 46894 -12520
rect 47340 -12762 47434 -12520
rect 44634 -14146 46414 -13428
rect 31938 -14184 39760 -14170
rect 40816 -14184 41550 -14170
rect 44018 -14184 46414 -14146
rect 31938 -14232 46414 -14184
rect 31938 -14292 45418 -14232
rect 45488 -14292 46414 -14232
rect 31938 -14750 46414 -14292
rect 31938 -14802 41228 -14750
rect 31938 -15190 35120 -14802
rect 35396 -15138 41228 -14802
rect 41504 -15138 46414 -14750
rect 35396 -15190 46414 -15138
rect 31938 -15544 46414 -15190
rect 31938 -15604 45384 -15544
rect 45454 -15604 46414 -15544
rect 31938 -15780 46414 -15604
rect 46738 -13808 47434 -12762
rect 47826 -11248 49606 -11072
rect 47826 -12258 49610 -11248
rect 47826 -12318 48738 -12258
rect 48808 -12318 49610 -12258
rect 47826 -12570 49610 -12318
rect 47826 -13116 49606 -12570
rect 54580 -12812 55310 -10352
rect 55430 -11588 55700 -10074
rect 55430 -11874 55462 -11588
rect 55670 -11874 55700 -11588
rect 54562 -12880 55328 -12812
rect 46738 -14050 46866 -13808
rect 47312 -14050 47434 -13808
rect 46738 -14466 47434 -14050
rect 46738 -14708 46888 -14466
rect 47334 -14708 47434 -14466
rect 46738 -15120 47434 -14708
rect 46738 -15362 46894 -15120
rect 47340 -15362 47434 -15120
rect 46738 -15748 47434 -15362
rect 47826 -13572 49606 -13426
rect 47826 -13632 48744 -13572
rect 48814 -13632 49606 -13572
rect 47826 -14010 49606 -13632
rect 54562 -13714 54646 -12880
rect 55214 -13714 55328 -12880
rect 47826 -14886 49610 -14010
rect 54562 -14092 55328 -13714
rect 47826 -14946 48742 -14886
rect 48812 -14946 49610 -14886
rect 47826 -15332 49610 -14946
rect 47826 -15682 49606 -15332
rect 47826 -15754 49608 -15682
rect 31938 -15932 44574 -15780
rect 31938 -15950 39760 -15932
rect 40816 -15950 41550 -15932
rect 35850 -16364 37590 -16328
rect 41438 -16364 42394 -16324
rect 32018 -16378 42394 -16364
rect 47832 -16378 49608 -15754
rect 32018 -16430 49608 -16378
rect 32018 -16980 33348 -16430
rect 34172 -16436 39402 -16430
rect 34172 -16980 36396 -16436
rect 32018 -16986 36396 -16980
rect 37220 -16980 39402 -16436
rect 40226 -16506 49608 -16430
rect 40226 -16854 41718 -16506
rect 42156 -16854 49608 -16506
rect 54580 -16320 55310 -14092
rect 54580 -16424 54878 -16320
rect 55004 -16424 55310 -16320
rect 54580 -16674 55310 -16424
rect 54580 -16688 55006 -16674
rect 55232 -16688 55310 -16674
rect 55430 -14708 55700 -11874
rect 55430 -14994 55456 -14708
rect 55664 -14994 55700 -14708
rect 55430 -16472 55700 -14994
rect 55832 -13006 56562 -9954
rect 55832 -13184 57222 -13006
rect 55832 -13266 56844 -13184
rect 55832 -13370 56122 -13266
rect 56248 -13370 56844 -13266
rect 55832 -13414 56844 -13370
rect 57096 -13414 57222 -13184
rect 55832 -13650 57222 -13414
rect 55430 -16688 55702 -16472
rect 55832 -16688 56562 -13650
rect 40226 -16980 49608 -16854
rect 37220 -16982 49608 -16980
rect 37220 -16986 42394 -16982
rect 32018 -17042 42394 -16986
rect 32018 -17060 41558 -17042
rect 35850 -17066 37600 -17060
rect 31154 -18022 41558 -17466
rect 31154 -18552 31458 -18022
rect 31864 -18044 41558 -18022
rect 31864 -18552 32084 -18044
rect 31154 -18724 32084 -18552
rect 32366 -18058 41558 -18044
rect 32366 -18478 38190 -18058
rect 38446 -18478 41558 -18058
rect 32366 -18724 41558 -18478
rect 31154 -19246 41558 -18724
rect 47832 -21762 49608 -16982
rect 55444 -17022 55702 -16688
rect 55432 -17236 55718 -17022
rect 55432 -17458 55462 -17236
rect 55682 -17458 55718 -17236
rect 55432 -17494 55718 -17458
rect 55444 -17710 55708 -17494
rect 51268 -17758 55756 -17710
rect 51268 -18068 51318 -17758
rect 51674 -18068 55756 -17758
rect 51268 -18118 55756 -18068
rect 31164 -21784 35322 -21762
rect 36050 -21784 58054 -21762
rect 31164 -22052 58054 -21784
rect 31090 -22462 58054 -22052
rect 31090 -22466 39630 -22462
rect 31090 -22506 35074 -22466
rect 31090 -22512 33566 -22506
rect 31090 -22580 32050 -22512
rect 31164 -22660 32050 -22580
rect 32170 -22654 33566 -22512
rect 33686 -22614 35074 -22506
rect 35194 -22484 39630 -22466
rect 35194 -22488 38100 -22484
rect 35194 -22614 36600 -22488
rect 33686 -22636 36600 -22614
rect 36720 -22632 38100 -22488
rect 38220 -22610 39630 -22484
rect 39750 -22466 48720 -22462
rect 39750 -22610 41148 -22466
rect 38220 -22614 41148 -22610
rect 41268 -22474 45692 -22466
rect 41268 -22614 42658 -22474
rect 38220 -22622 42658 -22614
rect 42778 -22478 45692 -22474
rect 42778 -22622 44176 -22478
rect 38220 -22626 44176 -22622
rect 44296 -22614 45692 -22478
rect 45812 -22482 48720 -22466
rect 45812 -22614 47198 -22482
rect 44296 -22626 47198 -22614
rect 38220 -22630 47198 -22626
rect 47318 -22610 48720 -22482
rect 48840 -22470 58054 -22462
rect 48840 -22610 50246 -22470
rect 47318 -22618 50246 -22610
rect 50366 -22478 58054 -22470
rect 50366 -22618 51758 -22478
rect 47318 -22626 51758 -22618
rect 51878 -22488 58054 -22478
rect 51878 -22496 56304 -22488
rect 51878 -22626 53278 -22496
rect 47318 -22630 53278 -22626
rect 38220 -22632 53278 -22630
rect 36720 -22636 53278 -22632
rect 33686 -22644 53278 -22636
rect 53398 -22510 56304 -22496
rect 53398 -22644 54786 -22510
rect 33686 -22654 54786 -22644
rect 32170 -22658 54786 -22654
rect 54906 -22636 56304 -22510
rect 56424 -22502 58054 -22488
rect 56424 -22636 57812 -22502
rect 54906 -22650 57812 -22636
rect 57932 -22650 58054 -22502
rect 54906 -22658 58054 -22650
rect 32170 -22660 58054 -22658
rect 27716 -23376 30216 -23220
rect 31164 -23254 58054 -22660
rect 31164 -23274 35322 -23254
rect 36050 -23274 58054 -23254
rect 27716 -24392 27972 -23376
rect 28674 -23486 30216 -23376
rect 30668 -23486 31110 -23476
rect 28674 -23494 31110 -23486
rect 28674 -23638 58052 -23494
rect 28674 -23652 40676 -23638
rect 28674 -23676 33070 -23652
rect 28674 -23756 31568 -23676
rect 28674 -24126 29836 -23756
rect 30200 -24126 31568 -23756
rect 28674 -24184 31568 -24126
rect 31890 -24184 32322 -23676
rect 32644 -24160 33070 -23676
rect 33392 -23672 36112 -23652
rect 33392 -23686 34580 -23672
rect 33392 -24160 33842 -23686
rect 32644 -24184 33842 -24160
rect 28674 -24194 33842 -24184
rect 34164 -24180 34580 -23686
rect 34902 -23676 36112 -23672
rect 34902 -24180 35352 -23676
rect 34164 -24184 35352 -24180
rect 35674 -24160 36112 -23676
rect 36434 -24160 36880 -23652
rect 37202 -23660 40676 -23652
rect 37202 -23664 39898 -23660
rect 37202 -24160 37620 -23664
rect 35674 -24172 37620 -24160
rect 37942 -23666 39898 -23664
rect 37942 -23672 39152 -23666
rect 37942 -24172 38374 -23672
rect 35674 -24180 38374 -24172
rect 38696 -24174 39152 -23672
rect 39474 -24168 39898 -23666
rect 40220 -24146 40676 -23660
rect 40998 -23640 58052 -23638
rect 40998 -23656 52776 -23640
rect 40998 -23658 42186 -23656
rect 40998 -24146 41402 -23658
rect 40220 -24166 41402 -24146
rect 41724 -24164 42186 -23658
rect 42508 -23658 52776 -23656
rect 42508 -23664 51268 -23658
rect 42508 -24164 42938 -23664
rect 41724 -24166 42938 -24164
rect 40220 -24168 42938 -24166
rect 39474 -24172 42938 -24168
rect 43260 -23666 51268 -23664
rect 43260 -23672 50502 -23666
rect 43260 -24172 43682 -23672
rect 39474 -24174 43682 -24172
rect 38696 -24180 43682 -24174
rect 44004 -23674 50502 -23672
rect 44004 -23676 49754 -23674
rect 44004 -23684 48232 -23676
rect 44004 -23690 45216 -23684
rect 44004 -24180 44422 -23690
rect 35674 -24184 44422 -24180
rect 34164 -24194 44422 -24184
rect 28674 -24198 44422 -24194
rect 44744 -24192 45216 -23690
rect 45538 -23696 48232 -23684
rect 45538 -24192 45978 -23696
rect 44744 -24198 45978 -24192
rect 28674 -24204 45978 -24198
rect 46300 -23710 48232 -23696
rect 46300 -24204 46722 -23710
rect 28674 -24218 46722 -24204
rect 47044 -23712 48232 -23710
rect 47044 -24218 47496 -23712
rect 28674 -24220 47496 -24218
rect 47818 -24184 48232 -23712
rect 48554 -23678 49754 -23676
rect 48554 -24184 49026 -23678
rect 47818 -24186 49026 -24184
rect 49348 -24182 49754 -23678
rect 50076 -24174 50502 -23674
rect 50824 -24166 51268 -23666
rect 51590 -23660 52776 -23658
rect 51590 -24166 52038 -23660
rect 50824 -24168 52038 -24166
rect 52360 -24148 52776 -23660
rect 53098 -23660 58052 -23640
rect 53098 -24148 53536 -23660
rect 52360 -24168 53536 -24148
rect 53858 -23674 55816 -23660
rect 53858 -23686 55060 -23674
rect 53858 -24168 54324 -23686
rect 50824 -24174 54324 -24168
rect 50076 -24182 54324 -24174
rect 49348 -24186 54324 -24182
rect 47818 -24194 54324 -24186
rect 54646 -24182 55060 -23686
rect 55382 -24168 55816 -23674
rect 56138 -23682 58052 -23660
rect 56138 -24168 56564 -23682
rect 55382 -24182 56564 -24168
rect 54646 -24190 56564 -24182
rect 56886 -23704 58052 -23682
rect 56886 -24190 57316 -23704
rect 54646 -24194 57316 -24190
rect 47818 -24212 57316 -24194
rect 57638 -24212 58052 -23704
rect 47818 -24220 58052 -24212
rect 28674 -24346 58052 -24220
rect 28674 -24348 30760 -24346
rect 28674 -24392 30216 -24348
rect 31098 -24356 58052 -24346
rect 27716 -24588 30216 -24392
rect 31172 -24608 43064 -24604
rect 43350 -24608 44064 -24604
rect 44418 -24608 58192 -24604
rect 31172 -24932 58192 -24608
rect 31172 -25312 54610 -24932
rect 31172 -25332 43424 -25312
rect 31172 -25480 31296 -25332
rect 31416 -25340 43424 -25332
rect 31416 -25480 32808 -25340
rect 31172 -25488 32808 -25480
rect 32928 -25358 43424 -25340
rect 32928 -25372 38876 -25358
rect 32928 -25488 34322 -25372
rect 31172 -25520 34322 -25488
rect 34442 -25520 35840 -25372
rect 35960 -25374 38876 -25372
rect 35960 -25520 37354 -25374
rect 31172 -25522 37354 -25520
rect 37474 -25506 38876 -25374
rect 38996 -25388 43424 -25358
rect 38996 -25506 40392 -25388
rect 37474 -25522 40392 -25506
rect 31172 -25536 40392 -25522
rect 40512 -25390 43424 -25388
rect 40512 -25536 41898 -25390
rect 31172 -25538 41898 -25536
rect 42018 -25460 43424 -25390
rect 43544 -25336 54610 -25312
rect 43544 -25460 44932 -25336
rect 42018 -25484 44932 -25460
rect 45052 -25338 52512 -25336
rect 45052 -25350 51004 -25338
rect 45052 -25368 49480 -25350
rect 45052 -25372 47966 -25368
rect 45052 -25484 46450 -25372
rect 42018 -25520 46450 -25484
rect 46570 -25516 47966 -25372
rect 48086 -25498 49480 -25368
rect 49600 -25486 51004 -25350
rect 51124 -25484 52512 -25338
rect 52632 -25348 54610 -25336
rect 52632 -25484 54034 -25348
rect 51124 -25486 54034 -25484
rect 49600 -25496 54034 -25486
rect 54154 -25496 54610 -25348
rect 49600 -25498 54610 -25496
rect 48086 -25516 54610 -25498
rect 46570 -25520 54610 -25516
rect 42018 -25538 54610 -25520
rect 31172 -25766 54610 -25538
rect 55178 -25350 58192 -24932
rect 55178 -25498 55548 -25350
rect 55668 -25366 58192 -25350
rect 55668 -25498 57066 -25366
rect 55178 -25514 57066 -25498
rect 57186 -25514 58192 -25366
rect 55178 -25766 58192 -25514
rect 31172 -26094 58192 -25766
rect 31172 -26112 57598 -26094
rect 31172 -26116 43064 -26112
rect 43346 -26128 44068 -26112
rect 44418 -26116 57598 -26112
rect 31210 -29004 60790 -28128
rect 31210 -30500 40896 -29004
rect 44220 -30500 60790 -29004
rect 31210 -31714 60790 -30500
<< via2 >>
rect 54600 -1104 55168 -908
rect 54600 -1252 54842 -1104
rect 54842 -1252 54962 -1104
rect 54962 -1252 55168 -1104
rect 54600 -1742 55168 -1252
rect 28412 -3024 29010 -2266
rect 46932 -7310 47314 -6920
rect 41676 -9844 42114 -9496
rect 58362 -7908 59962 -6218
rect 54646 -13714 55214 -12880
rect 41718 -16854 42156 -16506
rect 51318 -18068 51674 -17758
rect 27972 -24392 28674 -23376
rect 54610 -25766 55178 -24932
<< metal3 >>
rect 54468 -700 55254 -692
rect 54468 -908 55282 -700
rect 27778 -2266 29666 -1200
rect 27778 -3024 28412 -2266
rect 29010 -3024 29666 -2266
rect 27778 -4180 29666 -3024
rect 54468 -1742 54600 -908
rect 55168 -1742 55282 -908
rect 27804 -6920 47430 -6830
rect 27804 -7310 46932 -6920
rect 47314 -7310 47430 -6920
rect 27804 -7544 47430 -7310
rect 41574 -9496 42288 -9328
rect 41574 -9844 41676 -9496
rect 42114 -9844 42288 -9496
rect 41574 -16506 42288 -9844
rect 41574 -16854 41718 -16506
rect 42156 -16854 42288 -16506
rect 41574 -17040 42288 -16854
rect 54468 -12880 55254 -1742
rect 58186 -6218 61184 -4710
rect 58186 -7908 58362 -6218
rect 59962 -7908 61184 -6218
rect 58186 -9752 61184 -7908
rect 54468 -13714 54646 -12880
rect 55214 -13714 55282 -12880
rect 51236 -17636 51758 -17582
rect 27580 -17758 51758 -17636
rect 27580 -18068 51318 -17758
rect 51674 -18068 51758 -17758
rect 27580 -18188 51758 -18068
rect 27580 -18220 51730 -18188
rect 27400 -23376 29382 -22430
rect 27400 -24392 27972 -23376
rect 28674 -24392 29382 -23376
rect 27400 -25548 29382 -24392
rect 54468 -24932 55282 -13714
rect 54468 -25766 54610 -24932
rect 55178 -25766 55282 -24932
rect 54468 -25986 55282 -25766
use sky130_fd_pr__nfet_01v8_lvt_RM3WAQ  sky130_fd_pr__nfet_01v8_lvt_RM3WAQ_0
timestamp 1695195202
transform 1 0 44658 0 1 -2620
box -13432 -2496 13432 2496
use sky130_fd_pr__pfet_01v8_lvt_79GNHJ  XM1
timestamp 1695195202
transform 1 0 36748 0 1 -9709
box -4754 -3219 4754 3219
use sky130_fd_pr__pfet_01v8_lvt_79GNHJ  XM2
timestamp 1695195202
transform -1 0 36784 0 -1 -16695
box -4754 -3219 4754 3219
use sky130_fd_pr__nfet_01v8_lvt_9U978C  XM3
timestamp 1695195202
transform 0 1 55568 1 0 -13321
box -3225 -1210 3225 1210
use sky130_fd_pr__pfet_01v8_lvt_RM6ABE  XM4
timestamp 1695195202
transform 0 -1 47287 -1 0 -11958
box -1154 -3219 1154 3219
use sky130_fd_pr__pfet_01v8_lvt_RM6ABE  XM5
timestamp 1695195202
transform 0 1 47287 1 0 -14588
box -1154 -3219 1154 3219
use sky130_fd_pr__nfet_01v8_lvt_RM3WAQ  XM6
timestamp 1695195202
transform 1 0 44616 0 -1 -23968
box -13432 -2496 13432 2496
<< labels >>
flabel metal1 47012 -7176 47212 -6976 0 FreeSans 256 90 0 0 PCAS
port 0 nsew
flabel metal1 29132 -24022 29332 -23822 0 FreeSans 256 180 0 0 REF
port 2 nsew
flabel metal1 28706 -2732 28906 -2532 0 FreeSans 256 0 0 0 PIX
port 3 nsew
flabel metal1 55484 -18020 55684 -17820 0 FreeSans 256 270 0 0 GM_BIAS
port 4 nsew
rlabel metal3 27804 -7544 46932 -6830 1 PCAS
rlabel metal3 27778 -4180 28412 -1200 1 PIX
rlabel metal3 27400 -25548 27972 -22430 1 REF
rlabel metal3 27580 -18220 51318 -17636 1 GM_BIAS
rlabel metal3 59962 -9752 61184 -4710 1 OUT
port 7 nsew
rlabel metal2 28544 1668 58134 4684 1 VDD
port 5 nsew
rlabel metal2 31210 -31714 60790 -28128 1 GROUND
port 6 nsew
<< end >>
