magic
tech sky130A
timestamp 1698058409
<< locali >>
rect 7512 16935 8013 16978
rect 7512 16158 7547 16935
rect 7976 16158 8013 16935
rect 7512 6420 8013 16158
rect 10489 16891 10928 16946
rect 10489 16115 10536 16891
rect 10865 16115 10928 16891
rect 10489 3589 10928 16115
rect 17535 7039 18062 7109
rect 17535 6866 17639 7039
rect 17994 6866 18062 7039
rect 17535 6576 18062 6866
rect 17535 4794 18410 6576
rect 9689 -2398 10146 1520
rect 10429 -2398 10897 2888
rect 17535 2030 18062 4794
rect 23675 2713 25327 2720
rect 23675 2677 25353 2713
rect 23675 2290 23730 2677
rect 23988 2290 25353 2677
rect 23675 2246 25353 2290
rect 9688 -3068 10897 -2398
rect 17524 1259 18064 2030
rect 17524 960 18537 1259
rect 17524 -579 18064 960
rect 17524 -874 17586 -579
rect 18015 -874 18064 -579
rect 17524 -2509 18064 -874
rect 17514 -3068 18064 -2509
rect 24603 -2649 25353 2246
rect 9688 -3282 10875 -3068
rect 9688 -3648 9789 -3282
rect 10737 -3648 10875 -3282
rect 9688 -3710 10875 -3648
rect 17514 -3268 18052 -3068
rect 17514 -3621 17577 -3268
rect 17937 -3621 18052 -3268
rect 17514 -3724 18052 -3621
<< viali >>
rect 7547 16158 7976 16935
rect 10536 16115 10865 16891
rect 17639 6866 17994 7039
rect 23730 2290 23988 2677
rect 17586 -874 18015 -579
rect 9789 -3648 10737 -3282
rect 17577 -3621 17937 -3268
<< metal1 >>
rect 7527 16935 8000 16959
rect 7527 16158 7547 16935
rect 7976 16158 8000 16935
rect 7527 16116 8000 16158
rect 10426 16891 10963 16981
rect 10426 16115 10536 16891
rect 10865 16115 10963 16891
rect 10426 16099 10963 16115
rect 12058 16758 12639 16811
rect 12058 16132 12112 16758
rect 12594 16132 12639 16758
rect 12058 6863 12639 16132
rect 22946 16703 23504 16747
rect 22946 16132 22990 16703
rect 23452 16132 23504 16703
rect 17060 7039 18485 15795
rect 17060 6866 17639 7039
rect 17994 6866 18485 7039
rect 12058 6856 16895 6863
rect 12058 6752 16908 6856
rect 17060 6764 18485 6866
rect 16602 6563 16908 6752
rect 11908 2403 12089 2774
rect 11475 1365 12089 2403
rect 16460 -2908 17064 2486
rect 17944 2258 18476 6764
rect 22946 2777 23504 16132
rect 22946 2677 24040 2777
rect 22946 2290 23730 2677
rect 23988 2290 24040 2677
rect 22946 2253 24040 2290
rect 22955 2207 24040 2253
rect 17521 -579 18054 -510
rect 17521 -874 17586 -579
rect 18015 -874 18054 -579
rect 17521 -943 18054 -874
rect 9706 -3282 10854 -3206
rect 9706 -3648 9789 -3282
rect 10737 -3648 10854 -3282
rect 9706 -3710 10854 -3648
rect 17466 -3268 18047 -3199
rect 17466 -3621 17577 -3268
rect 17937 -3621 18047 -3268
rect 17466 -3724 18047 -3621
<< via1 >>
rect 7547 16158 7976 16935
rect 10536 16115 10865 16891
rect 12112 16132 12594 16758
rect 22990 16132 23452 16703
rect 11111 3155 11181 3228
rect 11774 -1009 11955 -481
rect 17586 -874 18015 -579
rect 9789 -3648 10737 -3282
rect 17577 -3621 17937 -3268
<< metal2 >>
rect 7314 16935 28629 18146
rect 7314 16158 7547 16935
rect 7976 16891 28629 16935
rect 7976 16158 10536 16891
rect 7314 16115 10536 16158
rect 10865 16758 28629 16891
rect 10865 16132 12112 16758
rect 12594 16703 28629 16758
rect 12594 16132 22990 16703
rect 23452 16132 28629 16703
rect 10865 16115 28629 16132
rect 7314 16078 28629 16115
rect 13069 12208 13442 13807
rect 13069 11703 13109 12208
rect 13371 11703 13442 12208
rect 13069 11658 13442 11703
rect 13047 7855 13480 9217
rect 13047 7343 13095 7855
rect 13412 7343 13480 7855
rect 13047 7303 13480 7343
rect 8327 4590 8706 4712
rect 8327 4286 8381 4590
rect 8535 4286 8706 4590
rect 8327 3155 8706 4286
rect 12606 4590 13047 4698
rect 12606 4299 12684 4590
rect 12969 4299 13047 4590
rect 12606 3908 13047 4299
rect 11100 3228 11188 3236
rect 11100 3155 11111 3228
rect 11181 3155 11188 3228
rect 11100 3145 11188 3155
rect 8422 1045 8705 1115
rect 8422 934 8485 1045
rect 8651 934 8705 1045
rect 8422 860 8705 934
rect 11429 -481 12086 1431
rect 12529 -100 13160 3908
rect 15726 1940 19708 15785
rect 21965 9098 28083 9186
rect 21965 8888 27657 9098
rect 28015 8888 28083 9098
rect 21965 8758 28083 8888
rect 11429 -1009 11774 -481
rect 11955 -1009 12086 -481
rect 11429 -2458 12086 -1009
rect 12606 -1012 13047 -100
rect 17521 -579 18054 -510
rect 17521 -874 17586 -579
rect 18015 -874 18054 -579
rect 17521 -943 18054 -874
rect 18101 -1321 18390 1940
rect 11428 -2484 12086 -2458
rect 11428 -3068 12130 -2484
rect 11463 -3197 12130 -3068
rect 7473 -3268 28559 -3197
rect 7473 -3282 17577 -3268
rect 7473 -3648 9789 -3282
rect 10737 -3621 17577 -3282
rect 17937 -3621 28559 -3268
rect 10737 -3648 28559 -3621
rect 7473 -5062 28559 -3648
<< via2 >>
rect 15471 13627 15548 13708
rect 13109 11703 13371 12208
rect 15465 9134 15553 9218
rect 13095 7343 13412 7855
rect 8381 4286 8535 4590
rect 12684 4299 12969 4590
rect 13601 4335 13682 4415
rect 10561 3185 10611 3227
rect 11118 3165 11174 3219
rect 8485 934 8651 1045
rect 19998 13593 20081 13702
rect 22073 13504 22476 13715
rect 19976 8951 20062 9033
rect 27657 8888 28015 9098
rect 20034 4398 20114 4487
rect 22111 4312 22509 4533
rect 13551 -813 13630 -735
rect 15750 -826 15945 -640
rect 17586 -874 18015 -579
rect 20964 -1249 21018 -1217
rect 18759 -2188 18814 -2129
<< metal3 >>
rect 10489 15146 10853 15152
rect 10275 14993 11082 15146
rect 10275 14448 20218 14993
rect 10275 14316 11082 14448
rect 10489 14315 10853 14316
rect 10489 14036 10853 14039
rect 10286 13822 11093 14036
rect 10286 13708 15667 13822
rect 10286 13627 15471 13708
rect 15548 13627 15667 13708
rect 10286 13412 15667 13627
rect 19894 13702 20215 14448
rect 19894 13593 19998 13702
rect 20081 13593 20215 13702
rect 19894 13534 20215 13593
rect 22022 13715 22506 13744
rect 22022 13504 22073 13715
rect 22476 13504 22506 13715
rect 22022 13471 22506 13504
rect 10286 13206 11093 13412
rect 10489 13163 10853 13206
rect 13079 12208 13435 12270
rect 13079 11703 13109 12208
rect 13371 11703 13435 12208
rect 13079 11658 13435 11703
rect 10489 10652 10853 10677
rect 10297 10439 11104 10652
rect 10297 10000 20253 10439
rect 10297 9822 11104 10000
rect 10489 9816 10853 9822
rect 10489 9565 10853 9570
rect 10308 9332 11115 9565
rect 10308 9218 15629 9332
rect 10308 9134 15465 9218
rect 15553 9134 15629 9218
rect 10308 8928 15629 9134
rect 19827 9033 20245 10000
rect 19827 8951 19976 9033
rect 20062 8951 20245 9033
rect 10308 8735 11115 8928
rect 19827 8890 20245 8951
rect 27624 9098 28035 9124
rect 27624 8888 27657 9098
rect 28015 8888 28035 9098
rect 27624 8852 28035 8888
rect 10489 8727 10853 8735
rect 10466 8500 10992 8501
rect 10308 7670 11115 8500
rect 13052 7855 13484 7909
rect 10466 6205 10992 7670
rect 13052 7343 13095 7855
rect 13412 7343 13484 7855
rect 13052 7310 13484 7343
rect 10466 5808 20302 6205
rect 8372 4590 8546 4629
rect 8372 4286 8381 4590
rect 8535 4286 8546 4590
rect 8372 4253 8546 4286
rect 12626 4590 12998 4618
rect 12626 4299 12684 4590
rect 12969 4299 12998 4590
rect 19905 4487 20294 5808
rect 12626 4259 12998 4299
rect 13563 4415 13718 4444
rect 13563 4335 13601 4415
rect 13682 4335 13718 4415
rect 10445 3227 10652 3274
rect 13563 3249 13718 4335
rect 19905 4398 20034 4487
rect 20114 4398 20294 4487
rect 19905 4314 20294 4398
rect 22083 4533 22548 4580
rect 22083 4312 22111 4533
rect 22509 4312 22548 4533
rect 22083 4276 22548 4312
rect 10445 3185 10561 3227
rect 10611 3185 10652 3227
rect 8422 1045 8705 1115
rect 8422 934 8485 1045
rect 8651 934 8705 1045
rect 8422 860 8705 934
rect 10445 -451 10652 3185
rect 11090 3219 13730 3249
rect 11090 3165 11118 3219
rect 11174 3165 13730 3219
rect 11090 3129 13730 3165
rect 10318 -598 10833 -451
rect 15676 -554 16008 -551
rect 10318 -619 11338 -598
rect 10318 -625 11442 -619
rect 12036 -625 12213 -619
rect 13440 -625 13658 -619
rect 10318 -735 13659 -625
rect 10318 -813 13551 -735
rect 13630 -813 13659 -735
rect 10318 -962 13659 -813
rect 15676 -640 16009 -554
rect 15676 -826 15750 -640
rect 15945 -826 16009 -640
rect 15676 -947 16009 -826
rect 17521 -579 18054 -510
rect 17521 -874 17586 -579
rect 18015 -874 18054 -579
rect 17521 -943 18054 -874
rect 15684 -948 16009 -947
rect 10318 -1037 10833 -962
rect 11308 -967 13659 -962
rect 20934 -1117 21094 -1079
rect 20934 -1276 20949 -1117
rect 21068 -1276 21094 -1117
rect 20934 -1282 21094 -1276
rect 17982 -2057 18864 -2032
rect 17977 -2129 18864 -2057
rect 17977 -2188 18759 -2129
rect 18814 -2188 18864 -2129
rect 17977 -2293 18864 -2188
rect 17829 -2303 18864 -2293
rect 17829 -2880 18431 -2303
<< via3 >>
rect 22073 13504 22476 13715
rect 13109 11703 13371 12208
rect 27681 8912 27987 9077
rect 13095 7343 13412 7855
rect 8396 4349 8528 4524
rect 12745 4315 12922 4514
rect 22111 4312 22509 4533
rect 15756 -823 15933 -656
rect 17586 -874 18015 -579
rect 20949 -1217 21068 -1117
rect 20949 -1249 20964 -1217
rect 20964 -1249 21018 -1217
rect 21018 -1249 21068 -1217
rect 20949 -1276 21068 -1249
<< metal4 >>
rect 21964 13715 25136 13792
rect 21964 13504 22073 13715
rect 22476 13504 25136 13715
rect 21964 13387 25136 13504
rect 13029 12208 25141 12268
rect 13029 11703 13109 12208
rect 13371 11703 25141 12208
rect 13029 11630 25141 11703
rect 27406 9077 28614 15785
rect 27386 8912 27681 9077
rect 27987 8912 28614 9077
rect 8164 7618 9090 8508
rect 12988 7855 25098 7910
rect 8360 4666 8907 7618
rect 12988 7343 13095 7855
rect 13412 7343 25098 7855
rect 12988 7198 25098 7343
rect 8341 4524 13032 4666
rect 8341 4349 8396 4524
rect 8528 4514 13032 4524
rect 8528 4349 12745 4514
rect 8341 4315 12745 4349
rect 12922 4315 13032 4514
rect 8341 4193 13032 4315
rect 22019 4533 25129 4616
rect 22019 4312 22111 4533
rect 22509 4312 25129 4533
rect 22019 4218 25129 4312
rect 27406 3009 28614 8912
rect 27417 749 28599 3009
rect 26784 727 28599 749
rect 23491 546 28599 727
rect 23491 541 27485 546
rect 26784 524 27485 541
rect 15684 -579 21172 -533
rect 15684 -656 17586 -579
rect 15684 -823 15756 -656
rect 15933 -823 17586 -656
rect 15684 -874 17586 -823
rect 18015 -823 21172 -579
rect 18015 -874 21174 -823
rect 15684 -934 21174 -874
rect 20897 -1117 21174 -934
rect 20897 -1276 20949 -1117
rect 21068 -1276 21174 -1117
rect 20897 -1300 21174 -1276
use switch  x1
timestamp 1698058409
transform 0 1 18403 1 0 2273
box -20 -459 4321 5137
use switch  x2
timestamp 1698058409
transform 0 1 11967 -1 0 6543
box -20 -459 4321 5137
use curr_mir  x3
timestamp 1698058334
transform 0 -1 12713 1 0 869
box 200 2565 6922 5195
use opamp  x4
timestamp 1696521366
transform 1 0 15179 0 -1 1876
box 3034 622 9644 4507
use switch  x5
timestamp 1698058409
transform 0 1 18348 1 0 6822
box -20 -459 4321 5137
use switch  x6
timestamp 1698058409
transform 0 1 11917 -1 0 1394
box -20 -459 4321 5137
use not  x7
timestamp 1696661316
transform 1 0 10262 0 1 3113
box 236 -289 934 518
use switch  x8
timestamp 1698058409
transform 0 1 18369 1 0 11474
box -20 -459 4321 5137
use switch  x9
timestamp 1698058409
transform 0 -1 17179 1 0 7009
box -20 -459 4321 5137
use switch  x10
timestamp 1698058409
transform 0 -1 17179 1 0 11496
box -20 -459 4321 5137
use sky130_fd_pr__cap_mim_m3_1_3HBNLG  XC1
timestamp 1695395215
transform 1 0 25926 0 1 4384
box -1593 -1520 1593 1520
use sky130_fd_pr__cap_mim_m3_1_3HBNLG  XC2
timestamp 1695395215
transform 1 0 25909 0 1 7705
box -1593 -1520 1593 1520
use sky130_fd_pr__cap_mim_m3_1_3HBNLG  XC3
timestamp 1695395215
transform 1 0 25916 0 1 11041
box -1593 -1520 1593 1520
use sky130_fd_pr__cap_mim_m3_1_3HBNLG  XC4
timestamp 1695395215
transform 1 0 25932 0 1 14223
box -1593 -1520 1593 1520
<< labels >>
rlabel metal4 27417 546 28599 8912 1 intout
port 7 nsew
rlabel metal3 17829 -2880 18431 -2293 1 opbias
port 13 nsew
rlabel metal3 10318 -1037 10833 -451 1 en
port 14 nsew
rlabel metal3 8422 860 8705 1115 1 Vtune
port 15 nsew
rlabel metal4 8164 7618 9090 8508 1 intin
port 16 nsew
rlabel metal2 7473 -5062 28559 -3197 1 VSS
port 18 nsew
rlabel metal2 7314 16078 28629 18146 1 VDD
port 17 nsew
rlabel metal3 10308 7670 11115 8500 1 sw1
port 12 nsew
rlabel metal3 10308 8735 11115 9565 1 sw2
port 11 nsew
rlabel metal3 10297 9822 11104 10652 1 rst
port 10 nsew
rlabel metal3 10286 13206 11093 14036 1 sw3
port 9 nsew
rlabel metal3 10275 14316 11082 15146 1 sw4
port 8 nsew
<< end >>
