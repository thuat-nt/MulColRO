magic
tech sky130A
magscale 1 2
timestamp 1694848836
<< pwell >>
rect -825 -260 825 260
<< nmoslvt >>
rect -629 -50 -29 50
rect 29 -50 629 50
<< ndiff >>
rect -687 38 -629 50
rect -687 -38 -675 38
rect -641 -38 -629 38
rect -687 -50 -629 -38
rect -29 38 29 50
rect -29 -38 -17 38
rect 17 -38 29 38
rect -29 -50 29 -38
rect 629 38 687 50
rect 629 -38 641 38
rect 675 -38 687 38
rect 629 -50 687 -38
<< ndiffc >>
rect -675 -38 -641 38
rect -17 -38 17 38
rect 641 -38 675 38
<< psubdiff >>
rect -789 190 -693 224
rect 693 190 789 224
rect -789 128 -755 190
rect 755 128 789 190
rect -789 -190 -755 -128
rect 755 -190 789 -128
rect -789 -224 -693 -190
rect 693 -224 789 -190
<< psubdiffcont >>
rect -693 190 693 224
rect -789 -128 -755 128
rect 755 -128 789 128
rect -693 -224 693 -190
<< poly >>
rect -629 122 -29 138
rect -629 88 -613 122
rect -45 88 -29 122
rect -629 50 -29 88
rect 29 122 629 138
rect 29 88 45 122
rect 613 88 629 122
rect 29 50 629 88
rect -629 -88 -29 -50
rect -629 -122 -613 -88
rect -45 -122 -29 -88
rect -629 -138 -29 -122
rect 29 -88 629 -50
rect 29 -122 45 -88
rect 613 -122 629 -88
rect 29 -138 629 -122
<< polycont >>
rect -613 88 -45 122
rect 45 88 613 122
rect -613 -122 -45 -88
rect 45 -122 613 -88
<< locali >>
rect -789 190 -693 224
rect 693 190 789 224
rect -789 128 -755 190
rect 755 128 789 190
rect -629 88 -613 122
rect -45 88 -29 122
rect 29 88 45 122
rect 613 88 629 122
rect -675 38 -641 54
rect -675 -54 -641 -38
rect -17 38 17 54
rect -17 -54 17 -38
rect 641 38 675 54
rect 641 -54 675 -38
rect -629 -122 -613 -88
rect -45 -122 -29 -88
rect 29 -122 45 -88
rect 613 -122 629 -88
rect -789 -190 -755 -128
rect 755 -190 789 -128
rect -789 -224 -693 -190
rect 693 -224 789 -190
<< viali >>
rect -613 88 -45 122
rect 45 88 613 122
rect -675 -38 -641 38
rect -17 -38 17 38
rect 641 -38 675 38
rect -613 -122 -45 -88
rect 45 -122 613 -88
<< metal1 >>
rect -625 122 -33 128
rect -625 88 -613 122
rect -45 88 -33 122
rect -625 82 -33 88
rect 33 122 625 128
rect 33 88 45 122
rect 613 88 625 122
rect 33 82 625 88
rect -681 38 -635 50
rect -681 -38 -675 38
rect -641 -38 -635 38
rect -681 -50 -635 -38
rect -23 38 23 50
rect -23 -38 -17 38
rect 17 -38 23 38
rect -23 -50 23 -38
rect 635 38 681 50
rect 635 -38 641 38
rect 675 -38 681 38
rect 635 -50 681 -38
rect -625 -88 -33 -82
rect -625 -122 -613 -88
rect -45 -122 -33 -88
rect -625 -128 -33 -122
rect 33 -88 625 -82
rect 33 -122 45 -88
rect 613 -122 625 -88
rect 33 -128 625 -122
<< properties >>
string FIXED_BBOX -772 -207 772 207
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 0.5 l 3.0 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
