magic
tech sky130A
magscale 1 2
timestamp 1694848836
<< nwell >>
rect -1154 -10186 1154 10186
<< pmoslvt >>
rect -958 -9967 -358 9967
rect -300 -9967 300 9967
rect 358 -9967 958 9967
<< pdiff >>
rect -1016 9955 -958 9967
rect -1016 -9955 -1004 9955
rect -970 -9955 -958 9955
rect -1016 -9967 -958 -9955
rect -358 9955 -300 9967
rect -358 -9955 -346 9955
rect -312 -9955 -300 9955
rect -358 -9967 -300 -9955
rect 300 9955 358 9967
rect 300 -9955 312 9955
rect 346 -9955 358 9955
rect 300 -9967 358 -9955
rect 958 9955 1016 9967
rect 958 -9955 970 9955
rect 1004 -9955 1016 9955
rect 958 -9967 1016 -9955
<< pdiffc >>
rect -1004 -9955 -970 9955
rect -346 -9955 -312 9955
rect 312 -9955 346 9955
rect 970 -9955 1004 9955
<< nsubdiff >>
rect -1118 10116 -1022 10150
rect 1022 10116 1118 10150
rect -1118 10054 -1084 10116
rect 1084 10054 1118 10116
rect -1118 -10116 -1084 -10054
rect 1084 -10116 1118 -10054
rect -1118 -10150 -1022 -10116
rect 1022 -10150 1118 -10116
<< nsubdiffcont >>
rect -1022 10116 1022 10150
rect -1118 -10054 -1084 10054
rect 1084 -10054 1118 10054
rect -1022 -10150 1022 -10116
<< poly >>
rect -958 10048 -358 10064
rect -958 10014 -942 10048
rect -374 10014 -358 10048
rect -958 9967 -358 10014
rect -300 10048 300 10064
rect -300 10014 -284 10048
rect 284 10014 300 10048
rect -300 9967 300 10014
rect 358 10048 958 10064
rect 358 10014 374 10048
rect 942 10014 958 10048
rect 358 9967 958 10014
rect -958 -10014 -358 -9967
rect -958 -10048 -942 -10014
rect -374 -10048 -358 -10014
rect -958 -10064 -358 -10048
rect -300 -10014 300 -9967
rect -300 -10048 -284 -10014
rect 284 -10048 300 -10014
rect -300 -10064 300 -10048
rect 358 -10014 958 -9967
rect 358 -10048 374 -10014
rect 942 -10048 958 -10014
rect 358 -10064 958 -10048
<< polycont >>
rect -942 10014 -374 10048
rect -284 10014 284 10048
rect 374 10014 942 10048
rect -942 -10048 -374 -10014
rect -284 -10048 284 -10014
rect 374 -10048 942 -10014
<< locali >>
rect -1118 10116 -1022 10150
rect 1022 10116 1118 10150
rect -1118 10054 -1084 10116
rect 1084 10054 1118 10116
rect -958 10014 -942 10048
rect -374 10014 -358 10048
rect -300 10014 -284 10048
rect 284 10014 300 10048
rect 358 10014 374 10048
rect 942 10014 958 10048
rect -1004 9955 -970 9971
rect -1004 -9971 -970 -9955
rect -346 9955 -312 9971
rect -346 -9971 -312 -9955
rect 312 9955 346 9971
rect 312 -9971 346 -9955
rect 970 9955 1004 9971
rect 970 -9971 1004 -9955
rect -958 -10048 -942 -10014
rect -374 -10048 -358 -10014
rect -300 -10048 -284 -10014
rect 284 -10048 300 -10014
rect 358 -10048 374 -10014
rect 942 -10048 958 -10014
rect -1118 -10116 -1084 -10054
rect 1084 -10116 1118 -10054
rect -1118 -10150 -1022 -10116
rect 1022 -10150 1118 -10116
<< viali >>
rect -942 10014 -374 10048
rect -284 10014 284 10048
rect 374 10014 942 10048
rect -1004 -9955 -970 9955
rect -346 -9955 -312 9955
rect 312 -9955 346 9955
rect 970 -9955 1004 9955
rect -942 -10048 -374 -10014
rect -284 -10048 284 -10014
rect 374 -10048 942 -10014
<< metal1 >>
rect -954 10048 -362 10054
rect -954 10014 -942 10048
rect -374 10014 -362 10048
rect -954 10008 -362 10014
rect -296 10048 296 10054
rect -296 10014 -284 10048
rect 284 10014 296 10048
rect -296 10008 296 10014
rect 362 10048 954 10054
rect 362 10014 374 10048
rect 942 10014 954 10048
rect 362 10008 954 10014
rect -1010 9955 -964 9967
rect -1010 -9955 -1004 9955
rect -970 -9955 -964 9955
rect -1010 -9967 -964 -9955
rect -352 9955 -306 9967
rect -352 -9955 -346 9955
rect -312 -9955 -306 9955
rect -352 -9967 -306 -9955
rect 306 9955 352 9967
rect 306 -9955 312 9955
rect 346 -9955 352 9955
rect 306 -9967 352 -9955
rect 964 9955 1010 9967
rect 964 -9955 970 9955
rect 1004 -9955 1010 9955
rect 964 -9967 1010 -9955
rect -954 -10014 -362 -10008
rect -954 -10048 -942 -10014
rect -374 -10048 -362 -10014
rect -954 -10054 -362 -10048
rect -296 -10014 296 -10008
rect -296 -10048 -284 -10014
rect 284 -10048 296 -10014
rect -296 -10054 296 -10048
rect 362 -10014 954 -10008
rect 362 -10048 374 -10014
rect 942 -10048 954 -10014
rect 362 -10054 954 -10048
<< properties >>
string FIXED_BBOX -1101 -10133 1101 10133
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 99.66666666666667 l 3.0 m 1 nf 3 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
