magic
tech sky130A
magscale 1 2
timestamp 1695461801
<< error_s >>
rect 9650 20788 10324 20801
rect 9019 20767 10324 20788
rect 9034 20625 9654 20767
rect 9704 20733 10238 20752
rect 9738 20718 10236 20733
rect 9025 20586 9654 20625
rect 8952 20500 9654 20586
rect 9025 20348 9654 20500
rect 9704 20693 10270 20699
rect 9704 20687 9738 20693
rect 10236 20687 10270 20693
rect 9704 20684 10270 20687
rect 9704 20612 9738 20684
rect 9861 20672 10113 20676
rect 9849 20653 10125 20672
rect 10075 20638 10086 20641
rect 9883 20623 10091 20638
rect 9759 20612 9840 20623
rect 9883 20619 10168 20623
rect 9704 20570 9744 20612
rect 9752 20576 9840 20612
rect 9899 20604 10086 20619
rect 10087 20576 10168 20619
rect 9752 20570 9772 20576
rect 9704 20396 9738 20570
rect 9806 20538 9840 20576
rect 10134 20538 10168 20576
rect 10075 20510 10086 20521
rect 9899 20476 10086 20510
rect 10236 20396 10270 20684
rect 9704 20362 10270 20396
rect 9025 20294 9059 20348
rect 9025 20160 9654 20294
rect 9034 19872 9654 20160
rect 9704 20242 10270 20276
rect 9704 20029 9738 20242
rect 10075 20162 10086 20173
rect 9752 20035 9754 20122
rect 9759 20100 9840 20147
rect 9899 20128 10086 20162
rect 10087 20100 10168 20147
rect 9806 20046 9840 20100
rect 10134 20063 10168 20100
rect 10126 20054 10178 20063
rect 10128 20050 10174 20054
rect 10134 20046 10168 20050
rect 9888 20041 10086 20045
rect 9899 20029 10075 20034
rect 10098 20029 10206 20035
rect 10236 20029 10270 20242
rect 9704 19995 10270 20029
rect 9704 19920 9738 19995
rect 10236 19920 10270 19995
rect 9704 19886 10270 19920
rect 9532 19268 9732 19278
rect 9504 19240 9760 19250
rect 9330 13062 10844 13076
rect 9064 13024 9088 13046
rect 9042 13000 9088 13024
rect 17152 13024 17176 13046
rect 17152 13000 17198 13024
rect 3964 11848 5144 12220
rect 9742 11572 9762 11630
rect 9770 11572 9790 11624
rect 9686 11332 10324 11572
rect 7414 11176 8294 11224
rect 7358 11120 8238 11168
rect 9742 11000 9744 11176
rect 9770 11028 9772 11148
rect 10162 11060 10196 11132
rect 10162 11056 10192 11060
rect 10218 11032 10224 11160
rect 10218 11028 10220 11032
rect 10209 10504 10624 10535
rect 6656 10499 10624 10504
rect 15280 10504 15701 10535
rect 15280 10499 20160 10504
rect 1585 10465 5421 10499
rect 6656 10470 20160 10499
rect 10209 10465 15701 10470
rect 1489 8699 1523 10403
rect 1965 10397 1999 10435
rect 5007 10413 5018 10424
rect 5030 10413 5041 10424
rect 5007 10397 5041 10413
rect 1665 10363 5341 10397
rect 1965 8699 1999 10363
rect 2068 10304 2124 10315
rect 2250 10304 2306 10315
rect 2726 10304 2782 10315
rect 2908 10304 2964 10315
rect 3384 10304 3429 10315
rect 3566 10304 3611 10315
rect 4042 10304 4087 10315
rect 4224 10304 4269 10315
rect 4700 10304 4745 10315
rect 4882 10304 4927 10315
rect 2079 10048 2800 10304
rect 2079 8699 2124 10048
rect 2140 8699 2168 9980
rect 2261 8699 2306 10048
rect 2737 8699 2782 10048
rect 2798 8699 2826 9980
rect 2854 8699 2882 9980
rect 2919 8699 2964 10304
rect 0 8665 3173 8699
rect 1489 2167 1523 8665
rect 1965 8644 1999 8665
rect 2079 8662 2124 8665
rect 2079 8644 2113 8662
rect 1603 8628 1650 8644
rect 1591 8597 1650 8628
rect 1681 8603 1728 8644
rect 1664 8597 1728 8603
rect 1965 8597 2012 8644
rect 2079 8597 2126 8644
rect 2140 8616 2168 8665
rect 2261 8662 2306 8665
rect 2737 8662 2782 8665
rect 2261 8644 2295 8662
rect 2737 8644 2771 8662
rect 2261 8597 2308 8644
rect 2339 8597 2386 8644
rect 2737 8597 2784 8644
rect 2798 8616 2826 8665
rect 2854 8616 2882 8665
rect 2919 8662 2964 8665
rect 2919 8644 2953 8662
rect 2919 8597 2966 8644
rect 2997 8597 3044 8644
rect 1591 8563 1728 8597
rect 1771 8563 2386 8597
rect 2429 8563 3044 8597
rect 1591 8557 1693 8563
rect 1591 8516 1649 8557
rect 1720 8529 1721 8563
rect 1603 8272 1637 8516
rect 1698 8504 1743 8515
rect 1603 6808 1643 8272
rect 1660 6864 1671 8216
rect 1603 2328 1637 6808
rect 1647 2652 1678 4054
rect 1703 2624 1706 4082
rect 1709 2316 1743 8504
rect 1965 2316 1999 8563
rect 2079 2328 2113 8563
rect 2261 2328 2295 8563
rect 2356 8504 2401 8515
rect 2367 6506 2401 8504
rect 2298 6498 2510 6506
rect 2298 6058 2710 6498
rect 2367 2316 2401 6058
rect 2498 6050 2710 6058
rect 2737 2328 2771 8563
rect 2919 2328 2953 8563
rect 3014 8504 3059 8515
rect 3025 6498 3059 8504
rect 3139 6506 3173 8665
rect 3361 8662 3376 9768
rect 3139 6498 3356 6506
rect 2974 6058 3356 6498
rect 2974 6050 3186 6058
rect 3025 2316 3059 6050
rect 1697 2269 1756 2316
rect 1965 2269 2012 2316
rect 2355 2269 2414 2316
rect 3013 2269 3071 2316
rect 1665 2235 3071 2269
rect 1597 2173 1620 2229
rect 1697 2219 1755 2235
rect 1709 2167 1743 2201
rect 1965 2167 1999 2235
rect 2302 2222 2413 2235
rect 2355 2220 2413 2222
rect 2330 2219 2413 2220
rect 3013 2219 3071 2235
rect 2330 2167 2361 2219
rect 3056 2204 3071 2219
rect 3139 2269 3173 6050
rect 3395 2328 3429 10304
rect 3460 4630 3488 9980
rect 3516 4630 3544 9980
rect 3460 2275 3488 4444
rect 3516 2275 3544 4444
rect 3577 2328 3611 10304
rect 3828 6498 3832 6506
rect 3840 6058 3844 6498
rect 4053 5364 4087 10304
rect 4053 5174 4098 5364
rect 4130 5174 4158 9980
rect 4186 5174 4214 9980
rect 4235 5364 4269 10304
rect 4711 8740 4745 10304
rect 4838 8740 4866 9980
rect 4893 8740 4927 10304
rect 5007 8740 5041 10363
rect 4656 8704 5553 8740
rect 6560 8704 6594 10408
rect 7036 10402 7070 10449
rect 8536 10408 8564 10428
rect 8592 10408 8620 10440
rect 9200 10408 9228 10428
rect 9256 10408 9284 10428
rect 9908 10408 9936 10428
rect 10078 10418 10089 10429
rect 10101 10418 10112 10429
rect 10078 10402 10112 10418
rect 7036 10368 10112 10402
rect 7036 8704 7070 10368
rect 7139 10318 7184 10329
rect 7321 10318 7366 10329
rect 7797 10318 7842 10329
rect 7979 10318 8024 10329
rect 8455 10318 8500 10329
rect 7150 8704 7184 10318
rect 7226 8704 7254 9980
rect 7332 8704 7366 10318
rect 7808 8704 7842 10318
rect 7878 8704 7906 9980
rect 7934 8704 7962 9980
rect 7990 8704 8024 10318
rect 4656 8670 8244 8704
rect 4656 6498 5553 8670
rect 6560 7010 6594 8670
rect 7036 8640 7070 8670
rect 7150 8640 7184 8670
rect 6674 8633 6712 8640
rect 6662 8618 6712 8633
rect 6752 8636 6790 8640
rect 6662 8602 6720 8618
rect 6752 8608 6792 8636
rect 6728 8602 6792 8608
rect 7036 8602 7074 8640
rect 7150 8602 7188 8640
rect 7226 8628 7254 8670
rect 7332 8640 7366 8670
rect 7808 8640 7842 8670
rect 7332 8602 7370 8640
rect 7410 8602 7448 8640
rect 7808 8602 7846 8640
rect 7878 8634 7906 8670
rect 7934 8634 7962 8670
rect 7990 8640 8024 8670
rect 7990 8602 8028 8640
rect 8068 8602 8106 8640
rect 6662 8568 6792 8602
rect 6842 8568 7448 8602
rect 7500 8568 8106 8602
rect 6662 8562 6764 8568
rect 6662 8530 6720 8562
rect 6784 8534 6792 8568
rect 6674 7992 6708 8530
rect 6769 8518 6814 8529
rect 6674 7164 6714 7992
rect 4316 6050 5553 6498
rect 5682 6372 6144 7010
rect 6158 6372 6620 7010
rect 6674 6942 6719 7164
rect 6674 6786 6714 6942
rect 6740 6842 6742 7936
rect 6780 7164 6814 8518
rect 6780 6942 6825 7164
rect 6830 6984 6852 7066
rect 6740 6832 6774 6842
rect 6674 6776 6774 6786
rect 6674 6504 6708 6776
rect 4235 5174 4280 5364
rect 3850 5142 4280 5174
rect 3850 5140 4269 5142
rect 3850 4642 3884 5140
rect 4053 5119 4087 5140
rect 4053 5072 4100 5119
rect 4026 5038 4100 5072
rect 4053 4990 4087 5038
rect 4092 4990 4121 4995
rect 3953 4979 3998 4990
rect 3964 4803 3998 4979
rect 4053 4979 4126 4990
rect 4130 4986 4158 5140
rect 4186 4986 4269 5140
rect 4053 4791 4087 4979
rect 4092 4803 4126 4979
rect 4092 4791 4121 4803
rect 4053 4787 4121 4791
rect 4206 4790 4269 4986
rect 4053 4744 4100 4787
rect 4026 4710 4100 4744
rect 4053 4642 4087 4710
rect 4130 4642 4158 4790
rect 4186 4642 4269 4790
rect 3850 4608 4269 4642
rect 4053 4558 4087 4608
rect 4130 4558 4158 4608
rect 4186 4558 4214 4608
rect 4235 4558 4269 4608
rect 3836 4014 4269 4558
rect 3836 3938 4280 4014
rect 4053 3796 4098 3938
rect 4053 2328 4087 3796
rect 4130 2275 4158 3938
rect 4186 2275 4214 3938
rect 4235 3796 4280 3938
rect 4235 2328 4269 3796
rect 4656 2269 5553 6050
rect 5740 6288 6090 6322
rect 5740 5808 5774 6288
rect 5932 6220 5970 6258
rect 5898 6186 5970 6220
rect 5843 6136 5888 6147
rect 5931 6136 5976 6147
rect 5854 5960 5888 6136
rect 5942 5960 5976 6136
rect 5932 5910 5970 5948
rect 5898 5876 5970 5910
rect 6056 5808 6090 6288
rect 6122 5814 6124 6356
rect 6560 6322 6594 6372
rect 6216 6288 6594 6322
rect 5740 5774 6090 5808
rect 6216 5808 6250 6288
rect 6408 6220 6446 6258
rect 6374 6186 6446 6220
rect 6319 6136 6364 6147
rect 6407 6136 6452 6147
rect 6330 5960 6364 6136
rect 6418 5960 6452 6136
rect 6408 5910 6446 5948
rect 6374 5876 6446 5910
rect 6532 5808 6594 6288
rect 6216 5774 6594 5808
rect 3139 2235 5553 2269
rect 2367 2167 2401 2201
rect 3025 2167 3059 2201
rect 3139 2167 3173 2235
rect 3460 2222 3488 2229
rect 3516 2222 3544 2229
rect 4130 2222 4158 2229
rect 4186 2222 4214 2229
rect 4656 2167 5553 2235
rect 1489 2133 5553 2167
rect 6560 2190 6594 5774
rect 6674 6192 6714 6504
rect 6732 6390 6742 6448
rect 6730 6304 6742 6390
rect 6732 6248 6742 6304
rect 6674 5814 6708 6192
rect 6768 6174 6774 6200
rect 6712 6144 6714 6174
rect 6712 6118 6774 6144
rect 6780 5814 6814 6942
rect 6674 5596 6719 5814
rect 6780 5742 6825 5814
rect 6780 5656 6894 5742
rect 6780 5596 6825 5656
rect 6674 5540 6714 5596
rect 6674 2342 6708 5540
rect 6718 2626 6746 4028
rect 6780 2330 6814 5596
rect 7036 2330 7070 8568
rect 7150 2342 7184 8568
rect 7332 2342 7366 8568
rect 7427 8518 7472 8529
rect 7438 6478 7472 8518
rect 7394 6474 7606 6478
rect 7394 6030 7796 6474
rect 7438 2330 7472 6030
rect 7584 6026 7796 6030
rect 7808 2342 7842 8568
rect 7990 2342 8024 8568
rect 8085 8518 8130 8529
rect 8096 6474 8130 8518
rect 8210 6478 8244 8670
rect 8210 6474 8444 6478
rect 8060 6030 8444 6474
rect 8060 6026 8272 6030
rect 8096 2330 8130 6026
rect 6768 2292 6826 2330
rect 7036 2292 7074 2330
rect 7426 2292 7484 2330
rect 8084 2298 8142 2330
rect 8012 2292 8142 2298
rect 8210 2292 8244 6026
rect 8466 2342 8500 10318
rect 8536 2298 8564 10362
rect 8592 2342 8620 10362
rect 8637 10318 8682 10329
rect 9113 10318 9158 10329
rect 8648 2342 8682 10318
rect 8708 6472 8920 6478
rect 8708 6030 9112 6472
rect 8900 6024 9112 6030
rect 9124 2342 9158 10318
rect 9200 2298 9228 10362
rect 9256 2298 9284 10362
rect 9295 10318 9340 10329
rect 9771 10318 9816 10329
rect 9306 2342 9340 10318
rect 9376 6460 9588 6472
rect 9376 6024 9756 6460
rect 9544 6012 9756 6024
rect 9782 2342 9816 10318
rect 9852 8578 9880 9794
rect 9852 2418 9880 4110
rect 9908 2298 9936 10362
rect 9953 10318 9998 10329
rect 9964 2342 9998 10318
rect 10078 2292 10112 10368
rect 10209 8699 10624 10465
rect 12113 10397 12147 10435
rect 13763 10413 13774 10424
rect 13786 10413 13797 10424
rect 13763 10397 13797 10413
rect 11737 10363 14173 10397
rect 10974 8699 10980 9794
rect 11017 8699 11051 8733
rect 11675 8699 11709 8733
rect 12113 8699 12147 10363
rect 12216 10304 12272 10315
rect 12322 10304 12378 10315
rect 12874 10304 12930 10315
rect 12980 10304 13036 10315
rect 13532 10304 13588 10315
rect 13638 10304 13694 10315
rect 12227 8699 12272 10304
rect 12284 8699 12295 9980
rect 12333 8699 12378 10304
rect 12885 8699 12930 10304
rect 12991 9980 13036 10304
rect 12957 8699 12970 9980
rect 12985 8699 13036 9980
rect 13543 8699 13588 10304
rect 13606 8699 13611 9980
rect 13649 8699 13694 10304
rect 13763 8699 13797 10363
rect 10209 8665 13797 8699
rect 10209 8597 10624 8665
rect 10974 8658 10980 8665
rect 11017 8644 11051 8665
rect 11675 8644 11709 8665
rect 10989 8631 11051 8644
rect 11647 8631 11709 8644
rect 10989 8603 11057 8631
rect 11647 8603 11715 8631
rect 10983 8597 11057 8603
rect 11067 8597 11085 8603
rect 11641 8597 11715 8603
rect 11725 8597 11743 8603
rect 12113 8597 12147 8665
rect 12227 8662 12272 8665
rect 12284 8664 12295 8665
rect 12333 8662 12378 8665
rect 12885 8662 12930 8665
rect 12227 8644 12267 8662
rect 12333 8644 12367 8662
rect 12227 8613 12274 8644
rect 12215 8603 12274 8613
rect 12305 8603 12367 8644
rect 12885 8644 12919 8662
rect 12957 8658 12970 8665
rect 12985 8662 13036 8665
rect 13543 8662 13588 8665
rect 12985 8644 13026 8662
rect 12885 8613 12932 8644
rect 12215 8602 12367 8603
rect 12215 8597 12274 8602
rect 12299 8597 12367 8602
rect 12873 8603 12932 8613
rect 12963 8603 13026 8644
rect 13543 8644 13577 8662
rect 13578 8644 13583 8662
rect 13543 8613 13590 8644
rect 13606 8634 13611 8665
rect 13649 8662 13694 8665
rect 13649 8644 13683 8662
rect 12873 8602 13026 8603
rect 12873 8597 12932 8602
rect 12957 8597 13025 8602
rect 13531 8597 13590 8613
rect 13621 8603 13683 8644
rect 13615 8597 13683 8603
rect 10209 8563 11057 8597
rect 11063 8563 11715 8597
rect 11721 8563 12367 8597
rect 12379 8563 13025 8597
rect 13037 8563 13683 8597
rect 10209 3498 10624 8563
rect 10983 8557 11001 8563
rect 11011 8529 11057 8563
rect 11067 8557 11085 8563
rect 11641 8557 11659 8563
rect 11669 8529 11715 8563
rect 11725 8557 11743 8563
rect 11017 3498 11051 8529
rect 11675 3698 11709 8529
rect 11654 3498 11728 3698
rect 10209 3464 10922 3498
rect 10209 2966 10624 3464
rect 10746 3396 10793 3443
rect 10708 3362 10793 3396
rect 10635 3303 10680 3314
rect 10763 3303 10808 3314
rect 10646 3127 10680 3303
rect 10774 3127 10808 3303
rect 10746 3068 10793 3115
rect 10708 3034 10793 3068
rect 10888 2966 10922 3464
rect 10209 2932 10922 2966
rect 11008 3464 11398 3498
rect 11008 3402 11051 3464
rect 11008 2966 11042 3402
rect 11222 3396 11269 3443
rect 11184 3362 11269 3396
rect 11111 3303 11156 3314
rect 11239 3303 11284 3314
rect 11122 3127 11156 3303
rect 11250 3127 11284 3303
rect 11222 3068 11269 3115
rect 11184 3034 11269 3068
rect 11364 2966 11398 3464
rect 11008 2932 11398 2966
rect 11484 3464 11874 3498
rect 11484 2966 11518 3464
rect 11564 3310 11582 3343
rect 11654 3319 11728 3464
rect 11654 3315 11743 3319
rect 11592 3314 11610 3315
rect 11654 3314 11756 3315
rect 11587 3303 11632 3314
rect 11598 3127 11632 3303
rect 11654 3127 11760 3314
rect 11654 3115 11756 3127
rect 11606 3114 11632 3115
rect 11634 3111 11743 3115
rect 11634 3086 11728 3111
rect 11654 3058 11728 3086
rect 11634 3044 11728 3058
rect 11634 2994 11724 3044
rect 11618 2980 11634 2982
rect 11675 2966 11709 2994
rect 11840 2966 11874 3464
rect 11484 2932 11874 2966
rect 10209 2882 10624 2932
rect 10209 2316 10936 2882
rect 10990 2316 11412 2882
rect 11466 2316 11888 2882
rect 10209 2292 11888 2316
rect 6736 2269 11888 2292
rect 12113 2316 12147 8563
rect 12215 8516 12273 8563
rect 12299 8557 12317 8563
rect 12327 8529 12367 8563
rect 12227 8272 12261 8516
rect 12227 6808 12267 8272
rect 12284 6864 12295 8216
rect 12227 2328 12261 6808
rect 12299 2960 12302 4054
rect 12327 2960 12330 4082
rect 12299 2652 12302 2760
rect 12327 2624 12330 2760
rect 12333 2316 12367 8529
rect 12873 8516 12931 8563
rect 12957 8557 12975 8563
rect 12985 8529 13025 8563
rect 12446 6498 12658 6506
rect 12446 6058 12808 6498
rect 12596 6050 12808 6058
rect 12885 4076 12919 8516
rect 12885 2562 12925 4076
rect 12885 2328 12919 2562
rect 12991 2316 13025 8529
rect 13531 8516 13589 8563
rect 13615 8557 13633 8563
rect 13643 8529 13683 8563
rect 13122 6050 13454 6498
rect 13543 2328 13577 8516
rect 13578 6806 13583 8214
rect 13606 6834 13611 8186
rect 13649 4098 13683 8529
rect 13643 2584 13683 4098
rect 13649 2316 13683 2584
rect 13763 6506 13797 8665
rect 15280 8704 15701 10465
rect 17184 10402 17218 10449
rect 18834 10418 18845 10429
rect 18857 10418 18868 10429
rect 18834 10402 18868 10418
rect 17184 10368 18868 10402
rect 16088 8704 16122 8738
rect 16746 8704 16780 8738
rect 17184 8704 17218 10368
rect 17287 10318 17332 10329
rect 17393 10318 17438 10329
rect 17945 10318 17990 10329
rect 18051 10318 18096 10329
rect 18603 10318 18648 10329
rect 18709 10318 18754 10329
rect 17298 9792 17332 10318
rect 17298 8704 17338 9792
rect 17364 8704 17366 9736
rect 17404 8704 17438 10318
rect 17956 8704 17990 10318
rect 18062 9810 18096 10318
rect 18028 8704 18048 9754
rect 18056 8704 18104 9810
rect 18614 9766 18648 10318
rect 18614 8704 18654 9766
rect 18672 8704 18682 9738
rect 18720 8704 18754 10318
rect 18834 8704 18868 10368
rect 15280 8670 18868 8704
rect 15280 8602 15701 8670
rect 16088 8640 16122 8670
rect 16746 8640 16780 8670
rect 16060 8636 16122 8640
rect 16718 8636 16780 8640
rect 16060 8608 16128 8636
rect 16718 8608 16786 8636
rect 16054 8602 16128 8608
rect 16138 8602 16156 8608
rect 16712 8602 16786 8608
rect 16796 8602 16814 8608
rect 17184 8602 17218 8670
rect 17298 8618 17338 8670
rect 17364 8636 17366 8670
rect 17404 8640 17438 8670
rect 17376 8636 17438 8640
rect 17364 8632 17438 8636
rect 17286 8608 17344 8618
rect 17376 8608 17438 8632
rect 17956 8640 17990 8670
rect 18028 8650 18048 8670
rect 18056 8640 18104 8670
rect 17956 8618 17994 8640
rect 17286 8602 17438 8608
rect 17944 8608 18002 8618
rect 18034 8608 18104 8640
rect 18614 8618 18654 8670
rect 18672 8636 18682 8670
rect 18720 8640 18754 8670
rect 18692 8636 18754 8640
rect 18672 8634 18754 8636
rect 17944 8602 18104 8608
rect 18602 8608 18660 8618
rect 18692 8608 18754 8634
rect 18602 8606 18754 8608
rect 18602 8602 18660 8606
rect 18686 8602 18754 8606
rect 15280 8568 16128 8602
rect 16134 8568 16786 8602
rect 16792 8568 17438 8602
rect 17450 8568 18096 8602
rect 18108 8568 18754 8602
rect 14474 6940 14864 6974
rect 13763 6406 13980 6506
rect 14474 6498 14508 6940
rect 14688 6872 14735 6919
rect 14650 6838 14735 6872
rect 14577 6779 14622 6790
rect 14705 6779 14750 6790
rect 14588 6603 14622 6779
rect 14716 6603 14750 6779
rect 14688 6544 14735 6591
rect 14650 6534 14735 6544
rect 14624 6510 14735 6534
rect 14624 6498 14714 6510
rect 14464 6470 14714 6498
rect 14464 6442 14676 6470
rect 14830 6442 14864 6940
rect 15280 6498 15701 8568
rect 16054 8562 16072 8568
rect 16082 8534 16128 8568
rect 16138 8562 16156 8568
rect 16712 8562 16730 8568
rect 16740 8534 16786 8568
rect 16796 8562 16814 8568
rect 14464 6408 14864 6442
rect 15110 6478 15701 6498
rect 13763 6274 14016 6406
rect 14464 6358 14676 6408
rect 15110 6406 15886 6478
rect 13763 6058 13980 6274
rect 12113 2269 12160 2316
rect 12321 2269 12380 2316
rect 12979 2269 13038 2316
rect 13637 2269 13695 2316
rect 6736 2262 13695 2269
rect 6736 2258 11057 2262
rect 6668 2196 6696 2252
rect 6768 2242 6826 2258
rect 6780 2190 6814 2224
rect 7036 2190 7070 2258
rect 7426 2242 7484 2258
rect 8084 2242 8142 2258
rect 8096 2227 8142 2242
rect 7402 2190 7432 2198
rect 7438 2190 7472 2224
rect 7478 2190 7510 2198
rect 8096 2190 8130 2227
rect 8210 2190 8244 2258
rect 8536 2246 8564 2252
rect 9200 2240 9228 2252
rect 9256 2246 9284 2252
rect 9908 2240 9936 2252
rect 10078 2242 10112 2258
rect 10078 2231 10089 2242
rect 10101 2231 10112 2242
rect 10209 2235 11057 2258
rect 10209 2190 10624 2235
rect 10983 2229 11001 2235
rect 11011 2201 11057 2235
rect 11067 2235 11694 2262
rect 11697 2257 11715 2262
rect 11725 2257 13695 2262
rect 11697 2242 13695 2257
rect 11067 2229 11085 2235
rect 6560 2167 10624 2190
rect 11017 2167 11051 2201
rect 11675 2197 11685 2235
rect 11699 2197 11709 2242
rect 11737 2235 13695 2242
rect 12113 2167 12147 2235
rect 12321 2219 12379 2235
rect 12926 2229 13037 2235
rect 12979 2220 13037 2229
rect 12954 2219 13037 2220
rect 13637 2219 13695 2235
rect 12954 2201 12985 2219
rect 13680 2204 13695 2219
rect 13763 2167 13797 6058
rect 14460 5738 14882 6358
rect 15038 6330 15886 6406
rect 15110 6050 15886 6330
rect 15280 6030 15886 6050
rect 14474 5140 14864 5174
rect 14474 4642 14508 5140
rect 14688 5072 14735 5119
rect 14650 5038 14735 5072
rect 14830 5112 14864 5140
rect 14577 4979 14622 4990
rect 14705 4979 14750 4990
rect 14588 4803 14622 4979
rect 14716 4803 14750 4979
rect 14688 4782 14735 4791
rect 14558 4766 14636 4782
rect 14688 4766 14768 4782
rect 14688 4754 14735 4766
rect 14586 4738 14636 4754
rect 14688 4744 14740 4754
rect 14650 4738 14740 4744
rect 14650 4710 14735 4738
rect 14830 4704 14898 5112
rect 14830 4642 14864 4704
rect 14474 4608 14864 4642
rect 14460 3938 14882 4558
rect 15280 2292 15701 6030
rect 16088 2330 16122 8534
rect 16746 7010 16780 8534
rect 16306 6372 16780 7010
rect 16340 6322 16552 6372
rect 16340 6288 16714 6322
rect 16340 6252 16552 6288
rect 16556 6252 16594 6258
rect 16340 6186 16594 6252
rect 16340 6026 16552 6186
rect 16555 6136 16600 6147
rect 16364 5808 16398 6026
rect 16478 5960 16512 6026
rect 16566 5960 16600 6136
rect 16556 5910 16594 5948
rect 16522 5876 16594 5910
rect 16680 5808 16714 6288
rect 16364 5774 16714 5808
rect 16746 2330 16780 6372
rect 16988 6330 16990 6418
rect 16060 2326 16122 2330
rect 16718 2326 16780 2330
rect 17184 2330 17218 8568
rect 17286 8530 17344 8568
rect 17370 8562 17388 8568
rect 17398 8534 17438 8568
rect 17298 7992 17332 8530
rect 17298 6776 17338 7992
rect 17364 6832 17366 7936
rect 17298 2342 17332 6776
rect 17404 2330 17438 8534
rect 17944 8530 18002 8568
rect 18028 8562 18046 8568
rect 18056 8534 18096 8568
rect 17542 6472 17754 6478
rect 17542 6030 17868 6472
rect 17656 6024 17868 6030
rect 17956 4054 17990 8530
rect 17956 2540 17996 4054
rect 17956 2342 17990 2540
rect 18062 2330 18096 8534
rect 18602 8530 18660 8568
rect 18686 8562 18704 8568
rect 18714 8534 18754 8568
rect 18614 7966 18648 8530
rect 18614 6806 18654 7966
rect 18672 6834 18682 7938
rect 18208 6460 18420 6474
rect 18208 6026 18512 6460
rect 18300 6012 18512 6026
rect 18614 2342 18648 6806
rect 18720 4090 18754 8534
rect 18714 2576 18754 4090
rect 18720 2330 18754 2576
rect 16060 2298 16128 2326
rect 16718 2298 16786 2326
rect 16054 2292 16128 2298
rect 16138 2292 16156 2298
rect 16712 2292 16786 2298
rect 16796 2292 16814 2298
rect 17184 2292 17222 2330
rect 17392 2292 17450 2330
rect 18050 2292 18108 2330
rect 18708 2292 18766 2330
rect 18834 2292 18868 8670
rect 19912 3534 19986 3678
rect 19252 2896 19714 3534
rect 19728 2896 20190 3534
rect 21290 2980 21410 3000
rect 21596 2982 21836 3534
rect 21596 2980 21886 2982
rect 21284 2952 21438 2972
rect 21596 2954 21836 2980
rect 21596 2952 21914 2954
rect 21596 2896 21836 2952
rect 19306 2812 19656 2846
rect 19306 2784 19340 2812
rect 19272 2750 19340 2784
rect 19306 2332 19340 2750
rect 19498 2744 19536 2782
rect 19464 2710 19536 2744
rect 19409 2660 19454 2671
rect 19497 2660 19542 2671
rect 19420 2484 19454 2660
rect 19508 2484 19542 2660
rect 19498 2434 19536 2472
rect 19464 2400 19536 2434
rect 19622 2332 19656 2812
rect 19306 2298 19656 2332
rect 19782 2812 20132 2846
rect 19782 2332 19816 2812
rect 19906 2760 19930 2778
rect 19974 2760 20012 2782
rect 19906 2744 20012 2760
rect 19924 2710 20012 2744
rect 19924 2694 19976 2710
rect 19930 2672 19972 2694
rect 19984 2672 19998 2676
rect 19885 2660 19918 2671
rect 19930 2660 19964 2672
rect 19896 2596 19964 2660
rect 19976 2671 20014 2672
rect 19896 2484 19970 2596
rect 19930 2472 19970 2484
rect 19976 2484 20018 2671
rect 19976 2472 20014 2484
rect 19930 2468 19972 2472
rect 19906 2450 19972 2468
rect 19974 2450 20012 2472
rect 19906 2434 20012 2450
rect 19924 2400 20012 2434
rect 19924 2384 19976 2400
rect 19930 2342 19964 2366
rect 20098 2332 20132 2812
rect 19782 2298 20132 2332
rect 15280 2258 16128 2292
rect 16134 2258 16786 2292
rect 16792 2258 19244 2292
rect 19334 2258 19902 2292
rect 15280 2190 15701 2258
rect 16054 2252 16072 2258
rect 16082 2224 16128 2258
rect 16138 2252 16156 2258
rect 16676 2252 16730 2258
rect 16740 2234 16786 2258
rect 16796 2252 16840 2258
rect 16704 2224 16812 2234
rect 16088 2190 16122 2224
rect 16746 2190 16780 2224
rect 17184 2190 17218 2258
rect 17392 2242 17450 2258
rect 18050 2242 18108 2258
rect 18708 2242 18766 2258
rect 18751 2227 18766 2242
rect 18834 2190 18868 2258
rect 15280 2167 20160 2190
rect 6560 2156 20160 2167
rect 1051 1978 1085 2012
rect 384 1944 774 1978
rect 384 1916 418 1944
rect 384 1508 452 1916
rect 598 1876 645 1923
rect 560 1842 645 1876
rect 487 1783 532 1794
rect 615 1783 660 1794
rect 498 1607 532 1783
rect 626 1607 660 1783
rect 598 1548 645 1595
rect 560 1514 645 1548
rect 384 1446 418 1508
rect 740 1446 774 1944
rect 384 1412 774 1446
rect 860 1944 1250 1978
rect 860 1446 894 1944
rect 1051 1910 1098 1923
rect 1051 1898 1108 1910
rect 1030 1842 1108 1898
rect 940 1790 958 1823
rect 1030 1799 1104 1842
rect 1030 1795 1119 1799
rect 968 1794 986 1795
rect 1030 1794 1132 1795
rect 963 1783 1008 1794
rect 974 1607 1008 1783
rect 1030 1788 1136 1794
rect 1030 1784 1142 1788
rect 1030 1607 1136 1784
rect 1030 1604 1132 1607
rect 1030 1595 1142 1604
rect 982 1594 1008 1595
rect 1010 1591 1119 1595
rect 1010 1582 1104 1591
rect 1010 1566 1108 1582
rect 1030 1538 1108 1566
rect 1010 1514 1108 1538
rect 1010 1474 1104 1514
rect 994 1460 1010 1462
rect 1030 1446 1104 1474
rect 1116 1446 1118 1591
rect 1216 1446 1250 1944
rect 860 1412 1250 1446
rect 1030 1362 1104 1412
rect -299 778 -276 852
rect -271 750 -248 852
rect 366 742 788 1362
rect 842 742 1264 1362
rect 3139 429 3173 2133
rect 4656 2097 5553 2133
rect 7438 542 7472 2156
rect 7702 1346 7706 1666
rect 7740 1346 7744 1666
rect 8096 542 8130 2156
rect 8210 452 8244 2156
rect 10209 2133 15701 2156
rect 10209 2120 10624 2133
rect 9104 1302 9344 1734
rect 8884 1282 8928 1302
rect 9104 1282 9404 1302
rect 9104 1268 9344 1282
rect 8884 1248 8894 1268
rect 9104 1248 9370 1268
rect 9104 1096 9344 1248
rect 13763 429 13797 2133
rect 15280 2097 15701 2133
rect 16088 542 16122 2156
rect 18062 542 18096 2156
rect 18834 452 18868 2156
rect 19728 1302 19968 1734
rect 19414 1282 19552 1302
rect 19728 1282 20028 1302
rect 19728 1268 19968 1282
rect 19448 1248 19518 1268
rect 19728 1248 19994 1268
rect 19728 1096 19968 1248
rect 0 0 200 44
rect -28 -28 228 -12
<< metal1 >>
rect 18616 30570 19744 30738
rect 5194 30338 5408 30390
rect 5194 30126 5242 30338
rect 5346 30126 5408 30338
rect 4402 16504 4670 16562
rect 4402 16386 4474 16504
rect 4596 16386 4670 16504
rect 4402 12478 4670 16386
rect 5194 12546 5408 30126
rect 18616 30216 18876 30570
rect 19496 30216 19744 30570
rect 6416 26036 6616 26060
rect 6416 25876 6428 26036
rect 6594 25876 6616 26036
rect 6416 25860 6616 25876
rect 5924 13738 6142 25550
rect 6464 16978 6664 16994
rect 6464 16806 6476 16978
rect 6648 16806 6664 16978
rect 6464 16794 6664 16806
rect 5914 12478 6108 12782
rect 4402 12464 6108 12478
rect 4402 12268 6114 12464
rect 5914 12264 6114 12268
rect 6544 11744 6754 12794
rect 6544 11532 6590 11744
rect 6694 11532 6754 11744
rect 6544 11480 6754 11532
rect 7414 11738 8536 22004
rect 18616 12220 19744 30216
rect 20522 20994 20722 21012
rect 20522 20832 20538 20994
rect 20706 20832 20722 20994
rect 20522 20812 20722 20832
rect 7414 11262 7642 11738
rect 8320 11262 8536 11738
rect 7414 11176 8536 11262
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
<< via1 >>
rect 5242 30126 5346 30338
rect 4474 16386 4596 16504
rect 18876 30216 19496 30570
rect 6428 25876 6594 26036
rect 6476 16806 6648 16978
rect 6590 11532 6694 11744
rect 20538 20832 20706 20994
rect 7642 11262 8320 11738
<< metal2 >>
rect 4240 30570 20872 33492
rect 4240 30338 18876 30570
rect 4240 30126 5242 30338
rect 5346 30216 18876 30338
rect 19496 30216 20872 30570
rect 5346 30126 20872 30216
rect 4240 30074 20872 30126
rect 6114 26036 10540 28732
rect 6114 25876 6428 26036
rect 6594 25876 10540 26036
rect 6114 25632 10540 25876
rect 5894 25484 6188 25538
rect 5894 25364 5976 25484
rect 6090 25364 6188 25484
rect 5894 25318 6188 25364
rect 11546 25516 11782 25550
rect 11546 25358 11580 25516
rect 11760 25358 11782 25516
rect 11546 25334 11782 25358
rect 15754 20994 20790 29664
rect 15754 20832 20538 20994
rect 20706 20832 20790 20994
rect 6130 16978 10556 19736
rect 6130 16806 6476 16978
rect 6648 16806 10556 16978
rect 6130 16636 10556 16806
rect 4384 16504 4702 16550
rect 4384 16386 4474 16504
rect 4596 16386 4702 16504
rect 4384 16330 4702 16386
rect 11578 16490 11778 16538
rect 11578 16358 11610 16490
rect 11752 16358 11778 16490
rect 11578 16288 11778 16358
rect 15754 12268 20790 20832
rect 4200 11744 20832 11840
rect 4200 11532 6590 11744
rect 6694 11738 20832 11744
rect 6694 11532 7642 11738
rect 4200 11262 7642 11532
rect 8320 11262 20832 11738
rect 4200 8422 20832 11262
<< via2 >>
rect 5976 25364 6090 25484
rect 11580 25358 11760 25516
rect 4474 16386 4596 16504
rect 11610 16358 11752 16490
<< metal3 >>
rect 5894 25516 11804 25562
rect 5894 25484 11580 25516
rect 5894 25364 5976 25484
rect 6090 25364 11580 25484
rect 5894 25358 11580 25364
rect 11760 25358 11804 25516
rect 5894 25312 11804 25358
rect 11550 16558 11810 16566
rect 4360 16504 11810 16558
rect 4360 16386 4474 16504
rect 4596 16490 11810 16504
rect 4596 16386 11610 16490
rect 4360 16358 11610 16386
rect 11752 16358 11810 16490
rect 4360 16308 11810 16358
rect 11550 16282 11810 16308
use not  not_0
timestamp 1695461801
transform 1 0 -476 0 1 1178
box 0 -578 1868 990
use not  not_1
timestamp 1695461801
transform 1 0 0 0 1 1178
box 0 -578 1868 990
use switch  switch_0
timestamp 1695461801
transform 1 0 1506 0 1 1550
box -114 -950 10510 11418
use switch  switch_1
timestamp 1695461801
transform 1 0 10262 0 1 1550
box -114 -950 10510 11418
use switch  switch_2
timestamp 1695461801
transform 1 0 1982 0 1 1550
box -114 -950 10510 11418
use switch  switch_3
timestamp 1695461801
transform 1 0 12130 0 1 1550
box -114 -950 10510 11418
use switch  switch_4
timestamp 1695461801
transform 1 0 -362 0 1 -250
box -114 -950 10510 11418
use switch  switch_5
timestamp 1695461801
transform 1 0 10262 0 1 -250
box -114 -950 10510 11418
use not  x1
timestamp 1695461801
transform 0 -1 6186 1 0 12070
box 0 -578 1868 990
use switch  x5
timestamp 1695461801
transform 0 1 8322 -1 0 29778
box -114 -950 10510 11418
use switch  x6
timestamp 1695461801
transform 0 1 8340 -1 0 20784
box -114 -950 10510 11418
<< labels >>
flabel metal1 5914 12264 6114 12464 0 FreeSans 256 0 0 0 SEL0
port 0 nsew
flabel metal1 6416 25860 6616 26060 0 FreeSans 256 0 0 0 IN0
port 3 nsew
flabel metal1 6464 16794 6664 16994 0 FreeSans 256 0 0 0 IN1
port 1 nsew
flabel metal1 20522 20812 20722 21012 0 FreeSans 256 0 0 0 OUT
port 2 nsew
rlabel metal2 4200 8422 20832 11840 1 GROUND
port 4 nsew
rlabel metal2 4240 30074 20872 33492 1 VDD
port 5 nsew
rlabel metal2 10488 9224 13228 10790 1 GROUND
rlabel metal2 10988 30990 13728 32556 1 VDD
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 SEL0
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 IN1
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 OUT
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 IN0
<< end >>
