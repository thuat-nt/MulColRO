magic
tech sky130A
magscale 1 2
timestamp 1696133064
<< pwell >>
rect -3225 -1210 3225 1210
<< nmoslvt >>
rect -3029 -1000 -29 1000
rect 29 -1000 3029 1000
<< ndiff >>
rect -3087 988 -3029 1000
rect -3087 -988 -3075 988
rect -3041 -988 -3029 988
rect -3087 -1000 -3029 -988
rect -29 988 29 1000
rect -29 -988 -17 988
rect 17 -988 29 988
rect -29 -1000 29 -988
rect 3029 988 3087 1000
rect 3029 -988 3041 988
rect 3075 -988 3087 988
rect 3029 -1000 3087 -988
<< ndiffc >>
rect -3075 -988 -3041 988
rect -17 -988 17 988
rect 3041 -988 3075 988
<< psubdiff >>
rect -3189 1140 -3093 1174
rect 3093 1140 3189 1174
rect -3189 1078 -3155 1140
rect 3155 1078 3189 1140
rect -3189 -1140 -3155 -1078
rect 3155 -1140 3189 -1078
rect -3189 -1174 -3093 -1140
rect 3093 -1174 3189 -1140
<< psubdiffcont >>
rect -3093 1140 3093 1174
rect -3189 -1078 -3155 1078
rect 3155 -1078 3189 1078
rect -3093 -1174 3093 -1140
<< poly >>
rect -3029 1072 -29 1088
rect -3029 1038 -3013 1072
rect -45 1038 -29 1072
rect -3029 1000 -29 1038
rect 29 1072 3029 1088
rect 29 1038 45 1072
rect 3013 1038 3029 1072
rect 29 1000 3029 1038
rect -3029 -1038 -29 -1000
rect -3029 -1072 -3013 -1038
rect -45 -1072 -29 -1038
rect -3029 -1088 -29 -1072
rect 29 -1038 3029 -1000
rect 29 -1072 45 -1038
rect 3013 -1072 3029 -1038
rect 29 -1088 3029 -1072
<< polycont >>
rect -3013 1038 -45 1072
rect 45 1038 3013 1072
rect -3013 -1072 -45 -1038
rect 45 -1072 3013 -1038
<< locali >>
rect -3189 1140 -3093 1174
rect 3093 1140 3189 1174
rect -3189 1078 -3155 1140
rect 3155 1078 3189 1140
rect -3029 1038 -3013 1072
rect -45 1038 -29 1072
rect 29 1038 45 1072
rect 3013 1038 3029 1072
rect -3075 988 -3041 1004
rect -3075 -1004 -3041 -988
rect -17 988 17 1004
rect -17 -1004 17 -988
rect 3041 988 3075 1004
rect 3041 -1004 3075 -988
rect -3029 -1072 -3013 -1038
rect -45 -1072 -29 -1038
rect 29 -1072 45 -1038
rect 3013 -1072 3029 -1038
rect -3189 -1140 -3155 -1078
rect 3155 -1140 3189 -1078
rect -3189 -1174 -3093 -1140
rect 3093 -1174 3189 -1140
<< viali >>
rect -3013 1038 -45 1072
rect 45 1038 3013 1072
rect -3075 -988 -3041 988
rect -17 -988 17 988
rect 3041 -988 3075 988
rect -3013 -1072 -45 -1038
rect 45 -1072 3013 -1038
<< metal1 >>
rect -3025 1072 -33 1078
rect -3025 1038 -3013 1072
rect -45 1038 -33 1072
rect -3025 1032 -33 1038
rect 33 1072 3025 1078
rect 33 1038 45 1072
rect 3013 1038 3025 1072
rect 33 1032 3025 1038
rect -3081 988 -3035 1000
rect -3081 -988 -3075 988
rect -3041 -988 -3035 988
rect -3081 -1000 -3035 -988
rect -23 988 23 1000
rect -23 -988 -17 988
rect 17 -988 23 988
rect -23 -1000 23 -988
rect 3035 988 3081 1000
rect 3035 -988 3041 988
rect 3075 -988 3081 988
rect 3035 -1000 3081 -988
rect -3025 -1038 -33 -1032
rect -3025 -1072 -3013 -1038
rect -45 -1072 -33 -1038
rect -3025 -1078 -33 -1072
rect 33 -1038 3025 -1032
rect 33 -1072 45 -1038
rect 3013 -1072 3025 -1038
rect 33 -1078 3025 -1072
<< properties >>
string FIXED_BBOX -3172 -1157 3172 1157
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 10.0 l 15.0 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
