magic
tech sky130A
magscale 1 2
timestamp 1696147843
<< locali >>
rect 476 892 1248 990
rect 476 810 528 892
rect 614 810 1248 892
rect 476 768 1248 810
rect 494 -432 1232 -360
rect 494 -518 550 -432
rect 636 -518 1232 -432
rect 494 -578 1232 -518
<< viali >>
rect 528 810 614 892
rect 550 -518 636 -432
<< metal1 >>
rect 476 892 662 990
rect 476 810 528 892
rect 614 810 662 892
rect 476 612 662 810
rect 1010 656 1082 708
rect 476 416 1008 612
rect 1102 426 1408 606
rect 994 360 1114 378
rect 994 296 1010 360
rect 1100 296 1114 360
rect 994 282 1114 296
rect 512 232 712 274
rect 512 156 614 232
rect 686 216 712 232
rect 1310 256 1408 426
rect 1668 256 1868 262
rect 686 156 714 216
rect 512 130 714 156
rect 512 74 712 130
rect 1006 78 1112 98
rect 1006 26 1030 78
rect 1086 26 1112 78
rect 1006 8 1112 26
rect 1310 70 1868 256
rect 1014 4 1090 8
rect 492 -224 1022 -30
rect 1310 -36 1408 70
rect 1668 62 1868 70
rect 1082 -216 1408 -36
rect 1310 -218 1408 -216
rect 492 -432 700 -224
rect 1020 -314 1086 -256
rect 492 -518 550 -432
rect 636 -518 700 -432
rect 492 -578 700 -518
<< via1 >>
rect 1010 296 1100 360
rect 614 156 686 232
rect 1030 26 1086 78
<< metal2 >>
rect 1024 380 1088 408
rect 984 360 1138 380
rect 984 296 1010 360
rect 1100 296 1138 360
rect 984 278 1138 296
rect 1024 250 1088 278
rect 584 232 1088 250
rect 584 156 614 232
rect 686 156 1088 232
rect 584 142 1088 156
rect 1024 88 1088 142
rect 1018 78 1098 88
rect 1018 26 1030 78
rect 1086 26 1098 78
rect 1018 14 1098 26
use sky130_fd_pr__nfet_01v8_lvt_648S5X  XM1 ~/ColRO/mag
timestamp 1695355038
transform 1 0 1053 0 1 -126
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_lvt_4QXNR3  XM10 ~/ColRO/mag
timestamp 1695355020
transform 1 0 1055 0 1 517
box -231 -319 231 319
<< labels >>
flabel metal1 512 74 712 274 0 FreeSans 256 0 0 0 in
port 1 nsew
flabel metal1 1668 62 1868 262 0 FreeSans 256 0 0 0 out
port 0 nsew
rlabel locali 846 -562 1138 -468 1 GROUND
port 3 nsew
rlabel locali 856 858 1178 968 1 VDD
port 4 nsew
<< end >>
