magic
tech sky130A
magscale 1 2
timestamp 1696521973
<< metal1 >>
rect 18242 15622 18442 15644
rect 18242 15462 18782 15622
rect 18242 15444 18442 15462
rect 30368 10020 30568 10032
rect 28176 9850 30568 10020
rect 30368 9832 30568 9850
rect 8546 9054 8746 9254
rect 15400 -10194 15600 -10176
rect 15400 -10368 15426 -10194
rect 15598 -10368 15600 -10194
rect 15400 -10376 15600 -10368
rect 38444 -10324 38644 -10310
rect 38444 -10484 38464 -10324
rect 38634 -10484 38644 -10324
rect 38444 -10510 38644 -10484
<< via1 >>
rect 15426 -10368 15598 -10194
rect 38464 -10484 38634 -10324
<< metal2 >>
rect 12744 3952 12920 3966
rect 12744 3804 12758 3952
rect 12908 3804 12920 3952
rect 12744 3788 12920 3804
rect 34400 3502 34564 3518
rect 34400 3356 34410 3502
rect 34556 3356 34564 3502
rect 34400 3344 34564 3356
rect 33838 -5848 34008 -5842
rect 33838 -6002 33848 -5848
rect 34000 -6002 34008 -5848
rect 33838 -6008 34008 -6002
rect 15376 -10160 15672 -10130
rect 15376 -10406 15386 -10160
rect 15642 -10406 15672 -10160
rect 15376 -10460 15672 -10406
rect 38434 -10324 38650 -10292
rect 38434 -10484 38464 -10324
rect 38634 -10484 38650 -10324
rect 38434 -10534 38650 -10484
<< via2 >>
rect 23046 13598 23186 13738
rect 12758 3804 12908 3952
rect 28254 3268 28488 3512
rect 29892 3316 30054 3476
rect 34410 3356 34556 3502
rect 12772 -720 12954 -534
rect 23090 -5928 23264 -5748
rect 33848 -6002 34000 -5848
rect 15386 -10194 15642 -10160
rect 15386 -10368 15426 -10194
rect 15426 -10368 15598 -10194
rect 15598 -10368 15642 -10194
rect 15386 -10406 15642 -10368
rect 23120 -10460 23336 -10226
rect 33866 -10514 34036 -10354
rect 38464 -10484 38634 -10324
rect 33870 -12134 34068 -11928
<< metal3 >>
rect 23002 13738 23246 13818
rect 23002 13598 23046 13738
rect 23186 13598 23246 13738
rect 23002 13558 23246 13598
rect 12748 3954 12916 3962
rect 12748 3798 12752 3954
rect 12910 3798 12916 3954
rect 12748 3792 12916 3798
rect 28220 3528 28514 3558
rect 28220 3252 28236 3528
rect 28500 3252 28514 3528
rect 28220 3226 28514 3252
rect 29846 3476 30122 3556
rect 29846 3316 29892 3476
rect 30054 3316 30122 3476
rect 34396 3502 34564 3518
rect 34396 3494 34410 3502
rect 34396 3356 34404 3494
rect 34556 3356 34564 3502
rect 34396 3350 34564 3356
rect 12720 -466 15648 -464
rect 12720 -534 15704 -466
rect 12720 -720 12772 -534
rect 12954 -720 15704 -534
rect 12720 -850 15704 -720
rect 12696 -11766 13060 -1960
rect 15346 -10160 15704 -850
rect 29846 -1452 30122 3316
rect 28420 -1812 30124 -1452
rect 23054 -5736 23294 -5710
rect 23054 -5930 23086 -5736
rect 23272 -5930 23294 -5736
rect 23054 -5948 23294 -5930
rect 28422 -10124 28748 -1812
rect 29846 -1814 30122 -1812
rect 33838 -5848 34010 -5840
rect 33838 -6002 33848 -5848
rect 34000 -6002 34010 -5848
rect 33838 -6008 34010 -6002
rect 28422 -10158 28746 -10124
rect 23120 -10160 28746 -10158
rect 15346 -10406 15386 -10160
rect 15642 -10226 28746 -10160
rect 15642 -10406 23120 -10226
rect 15346 -10460 23120 -10406
rect 23336 -10460 28746 -10226
rect 15346 -10506 28746 -10460
rect 23120 -10508 28746 -10506
rect 33826 -10324 38696 -10256
rect 33826 -10354 38464 -10324
rect 33826 -10514 33866 -10354
rect 34036 -10484 38464 -10354
rect 38634 -10484 38696 -10324
rect 34036 -10514 38696 -10484
rect 33826 -10598 38696 -10514
rect 12696 -12152 23382 -11766
rect 33822 -11918 34098 -11900
rect 33822 -12148 33852 -11918
rect 34076 -12148 34098 -11918
rect 12696 -12164 13060 -12152
rect 33822 -12162 34098 -12148
<< via3 >>
rect 23046 13598 23186 13738
rect 12752 3952 12910 3954
rect 12752 3804 12758 3952
rect 12758 3804 12908 3952
rect 12908 3804 12910 3952
rect 12752 3798 12910 3804
rect 28236 3512 28500 3528
rect 28236 3268 28254 3512
rect 28254 3268 28488 3512
rect 28488 3268 28500 3512
rect 28236 3252 28500 3268
rect 34404 3356 34410 3494
rect 34410 3356 34550 3494
rect 23086 -5748 23272 -5736
rect 23086 -5928 23090 -5748
rect 23090 -5928 23264 -5748
rect 23264 -5928 23272 -5748
rect 23086 -5930 23272 -5928
rect 33848 -5994 33992 -5852
rect 33852 -11928 34076 -11918
rect 33852 -12134 33870 -11928
rect 33870 -12134 34068 -11928
rect 34068 -12134 34076 -11928
rect 33852 -12148 34076 -12134
<< metal4 >>
rect 16144 16964 23294 16966
rect 16026 16716 23294 16964
rect 16028 14456 16096 16716
rect 8546 9254 11426 9256
rect 8542 9054 11426 9254
rect 8542 8212 8746 9054
rect 12706 8212 12992 8214
rect 8542 7928 12994 8212
rect 12706 3954 12992 7928
rect 17542 6118 17768 13804
rect 22986 13738 23294 16716
rect 22986 13598 23046 13738
rect 23186 13598 23294 13738
rect 22986 13516 23294 13598
rect 38620 10038 39028 10040
rect 30372 9834 39028 10038
rect 28048 6778 28610 6782
rect 21602 6470 28610 6778
rect 17542 5810 18852 6118
rect 21602 5852 21978 6470
rect 12706 3798 12752 3954
rect 12910 3798 12992 3954
rect 12706 3702 12992 3798
rect 28048 3528 28610 6470
rect 38620 3600 39028 9834
rect 28048 3252 28236 3528
rect 28500 3252 28610 3528
rect 34330 3494 39030 3600
rect 34330 3356 34404 3494
rect 34550 3356 39030 3494
rect 34330 3282 39030 3356
rect 28048 3068 28610 3252
rect 24506 -348 24574 394
rect 24506 -438 24572 -348
rect 23014 -814 24572 -438
rect 23014 -1066 23348 -814
rect 28984 -1066 29276 -1062
rect 23000 -1360 29276 -1066
rect 23014 -5736 23348 -1360
rect 23014 -5930 23086 -5736
rect 23272 -5930 23348 -5736
rect 23014 -6026 23348 -5930
rect 28984 -11894 29276 -1360
rect 38620 -5776 39028 3282
rect 33774 -5852 39030 -5776
rect 33774 -5994 33848 -5852
rect 33992 -5994 39030 -5852
rect 33774 -6080 39030 -5994
rect 28984 -11918 34172 -11894
rect 28984 -12148 33852 -11918
rect 34076 -12148 34172 -11918
rect 28984 -12178 34172 -12148
rect 28984 -12182 29276 -12178
use opamp  x1
timestamp 1696521366
transform 1 0 11486 0 1 7460
box 6068 1244 19288 9014
use switch  x2
timestamp 1696147897
transform 0 1 26630 -1 0 7734
box -53 -918 8642 11418
use switch  x3
timestamp 1696147897
transform 1 0 29621 0 1 -13774
box -53 -918 8642 11418
use switch  x4
timestamp 1696147897
transform 1 0 18873 0 1 -13684
box -53 -918 8642 11418
use switch  x5
timestamp 1696147897
transform 1 0 8529 0 1 -3974
box -53 -918 8642 11418
use sky130_fd_pr__cap_mim_m3_1_3HBNLG  XC1
timestamp 1695395215
transform 1 0 12926 0 1 11654
box -3186 -3040 3186 3040
use sky130_fd_pr__cap_mim_m3_1_3HBNLG  XC2
timestamp 1695395215
transform 1 0 21408 0 1 3220
box -3186 -3040 3186 3040
<< labels >>
flabel metal1 18242 15444 18442 15644 0 FreeSans 256 0 0 0 opbias
port 0 nsew
flabel metal1 8546 9054 8746 9254 0 FreeSans 256 0 0 0 cdsin
port 1 nsew
flabel metal1 30368 9832 30568 10032 0 FreeSans 256 0 0 0 cdsout
port 2 nsew
flabel metal1 15400 -10376 15600 -10176 0 FreeSans 256 0 0 0 sw1
port 3 nsew
flabel metal1 38444 -10510 38644 -10310 0 FreeSans 256 0 0 0 sw2
port 4 nsew
<< end >>
