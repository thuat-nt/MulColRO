magic
tech sky130A
magscale 1 2
timestamp 1695461801
<< error_p >>
rect 124848 14750 124968 14770
rect 125154 14752 125394 15304
rect 125154 14750 125444 14752
rect 124842 14722 124996 14742
rect 125154 14724 125394 14750
rect 125154 14722 125472 14724
rect 125154 14666 125394 14722
rect 72208 -8188 72328 -8168
rect 72514 -8186 72754 -7634
rect 72514 -8188 72804 -8186
rect 72202 -8216 72356 -8196
rect 72514 -8214 72754 -8188
rect 72514 -8216 72832 -8214
rect 72514 -8272 72754 -8216
<< error_s >>
rect 32926 32698 32928 32748
rect 32954 32698 32956 32776
rect 32374 32458 33012 32698
rect 38140 32654 38142 32732
rect 38168 32654 38170 32704
rect 38084 32414 38722 32654
rect 32908 32152 32928 32272
rect 32936 32146 32956 32300
rect 38140 32102 38160 32256
rect 38168 32108 38188 32228
rect 55147 28845 55181 35209
rect 55261 28941 55295 28975
rect 55919 28941 55953 28975
rect 56577 28941 56611 28975
rect 57235 28941 57269 28975
rect 57893 28941 57927 35110
rect 58551 28941 58605 28975
rect 55211 28907 55215 28941
rect 55227 28907 58605 28941
rect 55115 27035 55181 28845
rect 55257 28855 55261 28873
rect 55257 28839 55307 28855
rect 55318 28845 55336 28860
rect 55346 28845 55364 28858
rect 55859 28839 55906 28886
rect 55915 28855 55919 28873
rect 55915 28839 55965 28855
rect 56517 28845 56564 28886
rect 56508 28839 56564 28845
rect 56573 28855 56577 28873
rect 56573 28839 56623 28855
rect 56638 28845 56644 28848
rect 56666 28845 56672 28858
rect 57175 28839 57222 28886
rect 57231 28855 57235 28873
rect 57231 28839 57281 28855
rect 57833 28845 57880 28886
rect 57893 28873 57927 28907
rect 57828 28839 57880 28845
rect 57889 28855 57927 28873
rect 57889 28839 57939 28855
rect 58491 28839 58538 28886
rect 55261 28805 55906 28839
rect 55919 28805 56564 28839
rect 56577 28805 57222 28839
rect 57235 28805 57880 28839
rect 57893 28805 58538 28839
rect 55261 28758 55307 28805
rect 55217 28746 55235 28758
rect 55261 28746 55295 28758
rect 55217 27134 55295 28746
rect 55318 27458 55336 28799
rect 55346 27430 55364 28799
rect 55919 28758 55965 28805
rect 56508 28799 56529 28805
rect 56536 28771 56557 28805
rect 56577 28758 56623 28805
rect 55876 28746 55907 28757
rect 55919 28746 55953 28758
rect 56534 28746 56565 28757
rect 56577 28746 56611 28758
rect 32948 24328 32954 24340
rect 33140 24328 33148 24340
rect 32920 24300 32954 24312
rect 33140 24300 33176 24312
rect 32410 23876 32976 23910
rect 32410 23781 32444 23876
rect 32781 23796 32792 23807
rect 32605 23793 32792 23796
rect 32605 23781 32781 23793
rect 32942 23781 32976 23876
rect 32376 23747 32976 23781
rect 32410 23554 32444 23747
rect 32465 23735 32593 23747
rect 32793 23735 32890 23747
rect 32465 23734 32546 23735
rect 32793 23734 32874 23735
rect 32512 23696 32546 23734
rect 32840 23696 32874 23734
rect 32502 23670 32554 23682
rect 32781 23668 32792 23679
rect 32474 23642 32582 23654
rect 32605 23634 32792 23668
rect 32926 23654 32928 23741
rect 32942 23554 32976 23747
rect 32410 23520 32976 23554
rect 33026 23719 33646 23924
rect 37784 23722 37914 23743
rect 33026 23502 33673 23719
rect 37598 23697 37914 23722
rect 38100 23697 38506 23743
rect 37626 23669 37914 23694
rect 38100 23669 38450 23694
rect 33639 23448 33673 23502
rect 32410 23400 32976 23434
rect 32410 23112 32444 23400
rect 32781 23320 32792 23331
rect 32465 23258 32546 23305
rect 32605 23286 32792 23320
rect 32793 23258 32874 23305
rect 32512 23220 32546 23258
rect 32840 23220 32874 23258
rect 32942 23206 32976 23400
rect 32781 23192 32792 23203
rect 32908 23192 32928 23206
rect 32605 23158 32792 23192
rect 32832 23178 32928 23192
rect 32936 23192 32976 23206
rect 33026 23296 33673 23448
rect 33026 23210 33728 23296
rect 33026 23192 33673 23210
rect 32936 23172 33673 23192
rect 32942 23164 32976 23172
rect 33026 23164 33673 23172
rect 32804 23151 33673 23164
rect 32804 23150 33646 23151
rect 32908 23144 33646 23150
rect 32567 23120 32819 23123
rect 32942 23112 32976 23144
rect 32410 23089 32976 23112
rect 32410 23078 32444 23089
rect 32942 23078 32976 23089
rect 32410 23077 32976 23078
rect 32444 23063 32942 23077
rect 32410 23044 32976 23063
rect 33026 23026 33646 23144
rect 37408 23128 38028 23550
rect 38078 23502 38644 23536
rect 38078 23180 38112 23502
rect 38449 23422 38460 23433
rect 38133 23360 38214 23407
rect 38273 23388 38460 23422
rect 38461 23360 38542 23407
rect 38180 23322 38214 23360
rect 38508 23322 38542 23360
rect 38449 23294 38460 23305
rect 38273 23260 38460 23294
rect 38610 23180 38644 23502
rect 38078 23146 38644 23180
rect 37466 23074 37484 23113
rect 37784 23085 37814 23120
rect 37840 23085 37842 23120
rect 37500 23074 37518 23079
rect 37408 23028 38028 23074
rect 38140 23060 38582 23094
rect 38078 23033 38644 23060
rect 37408 23026 38088 23028
rect 37408 23012 38146 23026
rect 37408 23000 38028 23012
rect 37408 22998 38060 23000
rect 37408 22965 38118 22998
rect 37408 22931 40320 22965
rect 37408 22895 38028 22931
rect 38078 22798 38118 22931
rect 38126 22804 38146 22924
rect 38180 22897 38214 22900
rect 38508 22897 38542 22900
rect 38078 22766 38112 22798
rect 38610 22766 38644 22931
rect 55115 22173 55149 27035
rect 55217 26973 55263 27134
rect 55816 27081 55826 28480
rect 55844 27109 55854 28452
rect 55887 27134 55953 28746
rect 56545 27134 56611 28746
rect 56638 27446 56644 28799
rect 56666 27418 56672 28799
rect 57235 28758 57281 28805
rect 57828 28799 57845 28805
rect 57856 28771 57873 28805
rect 57893 28758 57939 28805
rect 57192 28746 57223 28757
rect 57235 28746 57269 28758
rect 57850 28746 57881 28757
rect 57893 28746 57927 28758
rect 55887 27122 55921 27134
rect 56545 27122 56579 27134
rect 55875 27109 55934 27122
rect 55844 27100 55934 27109
rect 55941 27100 55972 27109
rect 55875 27081 55934 27100
rect 55816 27075 55934 27081
rect 55323 27041 55934 27075
rect 55969 27075 56000 27081
rect 56533 27075 56592 27122
rect 57126 27081 57146 28486
rect 57154 27109 57174 28458
rect 57203 27134 57269 28746
rect 57861 27134 57927 28746
rect 57960 27424 57964 28799
rect 57988 27396 57992 28799
rect 58508 28746 58539 28757
rect 58551 28746 58585 28907
rect 57203 27122 57237 27134
rect 57861 27122 57895 27134
rect 57191 27109 57250 27122
rect 57154 27106 57250 27109
rect 57257 27106 57282 27109
rect 57191 27081 57250 27106
rect 57126 27078 57250 27081
rect 57285 27078 57310 27081
rect 57191 27075 57250 27078
rect 57849 27075 57908 27122
rect 58448 27081 58468 28456
rect 58476 27081 58496 28428
rect 58519 27134 58585 28746
rect 58633 28845 58651 28907
rect 58665 28845 58699 35209
rect 60218 28850 60252 35214
rect 60332 28946 60366 28980
rect 60990 28946 61024 28980
rect 61648 28946 61682 28980
rect 62306 28946 62340 28980
rect 62964 28946 62998 28980
rect 63622 28946 63676 28980
rect 60282 28912 60286 28946
rect 60298 28912 63676 28946
rect 58519 27122 58553 27134
rect 58507 27075 58565 27122
rect 55969 27072 56592 27075
rect 55981 27041 56592 27072
rect 56639 27041 57250 27075
rect 57297 27041 57908 27075
rect 57955 27041 58565 27075
rect 55875 27025 55921 27041
rect 56533 27025 56579 27041
rect 57191 27025 57237 27041
rect 57849 27025 57895 27041
rect 58507 27025 58553 27041
rect 58633 27035 58699 28845
rect 60186 27058 60252 28850
rect 60328 28860 60332 28878
rect 60328 28844 60378 28860
rect 60930 28844 60968 28882
rect 60986 28860 60990 28878
rect 60986 28844 61036 28860
rect 61588 28850 61626 28882
rect 61578 28844 61626 28850
rect 61644 28860 61648 28878
rect 61644 28844 61694 28860
rect 62246 28844 62284 28882
rect 62302 28860 62306 28878
rect 62302 28844 62352 28860
rect 62904 28844 62942 28882
rect 62960 28860 62964 28878
rect 62960 28844 63010 28860
rect 63562 28844 63600 28882
rect 60332 28810 60968 28844
rect 60990 28840 61626 28844
rect 60990 28810 61628 28840
rect 60332 28772 60378 28810
rect 60990 28772 61036 28810
rect 61578 28804 61600 28810
rect 61606 28776 61628 28810
rect 61648 28810 62284 28844
rect 62306 28810 62942 28844
rect 62964 28810 63600 28844
rect 61648 28772 61694 28810
rect 62306 28772 62352 28810
rect 62900 28804 62916 28810
rect 62928 28776 62944 28804
rect 62964 28772 63010 28810
rect 60288 28760 60306 28772
rect 60332 28760 60366 28772
rect 60947 28760 60978 28771
rect 60990 28760 61024 28772
rect 61605 28760 61636 28771
rect 61648 28760 61682 28772
rect 62263 28760 62294 28771
rect 62306 28760 62340 28772
rect 62921 28760 62952 28771
rect 62964 28760 62998 28772
rect 60288 27148 60366 28760
rect 57861 26973 57895 27025
rect 55217 26939 58565 26973
rect 55229 22269 55263 22303
rect 55887 22269 55921 22303
rect 56545 22269 56579 22303
rect 57203 22269 57237 22303
rect 57861 22269 57895 26939
rect 58519 22269 58553 22303
rect 55197 22235 58587 22269
rect 55101 20671 55149 22173
rect 55229 22183 55263 22235
rect 55887 22214 55921 22235
rect 56545 22214 56579 22235
rect 57203 22214 57237 22235
rect 57861 22214 57895 22235
rect 58519 22214 58553 22235
rect 55845 22183 55921 22214
rect 56503 22183 56579 22214
rect 57161 22183 57237 22214
rect 57819 22183 57895 22214
rect 55229 22086 55275 22183
rect 55845 22167 55933 22183
rect 56503 22167 56591 22183
rect 57161 22167 57249 22183
rect 57819 22167 57907 22183
rect 58477 22167 58553 22214
rect 58633 22173 58667 27035
rect 59880 24746 59882 24794
rect 59852 24718 59882 24738
rect 60186 22178 60220 27058
rect 60288 26996 60334 27148
rect 60886 27104 60912 28224
rect 60914 27104 60940 28196
rect 60958 27148 61024 28760
rect 61616 27148 61682 28760
rect 60958 27136 60992 27148
rect 61616 27136 61650 27148
rect 60946 27098 60996 27136
rect 61050 27104 61068 27120
rect 61604 27098 61654 27136
rect 62206 27104 62222 28206
rect 62234 27104 62250 28178
rect 62274 27148 62340 28760
rect 62932 27148 62998 28760
rect 63030 27402 63036 28804
rect 63058 27374 63064 28804
rect 63579 28760 63610 28771
rect 63622 28760 63656 28912
rect 62274 27136 62308 27148
rect 62932 27136 62966 27148
rect 62262 27098 62312 27136
rect 62920 27098 62970 27136
rect 63514 27104 63538 28208
rect 63542 27104 63566 28180
rect 63590 27148 63656 28760
rect 63704 28850 63722 28912
rect 63736 28850 63770 32670
rect 63590 27136 63624 27148
rect 63578 27098 63628 27136
rect 60394 27064 60996 27098
rect 61052 27064 61654 27098
rect 61710 27064 62312 27098
rect 62368 27064 62970 27098
rect 63026 27064 63628 27098
rect 60946 27048 60992 27064
rect 61604 27048 61650 27064
rect 62262 27048 62308 27064
rect 62920 27048 62966 27064
rect 63578 27048 63624 27064
rect 63704 27058 63770 28850
rect 64324 27786 64444 27806
rect 64630 27788 64870 28340
rect 64630 27786 64920 27788
rect 64318 27758 64472 27778
rect 64630 27760 64870 27786
rect 64630 27758 64948 27760
rect 64630 27702 64870 27758
rect 60958 26996 60992 27048
rect 60288 26962 63636 26996
rect 60300 22274 60334 22308
rect 60958 22274 60992 26962
rect 61616 22274 61650 22308
rect 62274 22274 62308 22308
rect 62932 22274 62966 22308
rect 63590 22274 63624 22308
rect 60268 22240 63658 22274
rect 55277 22133 55933 22167
rect 55935 22133 56591 22167
rect 56593 22133 57249 22167
rect 57251 22133 57907 22167
rect 57909 22133 58553 22167
rect 55853 22127 55857 22133
rect 55881 22099 55885 22133
rect 55887 22086 55933 22133
rect 56545 22086 56591 22133
rect 57169 22127 57173 22133
rect 57197 22099 57201 22133
rect 57203 22086 57249 22133
rect 57861 22086 57907 22133
rect 58485 22127 58489 22133
rect 58513 22099 58517 22133
rect 55229 22074 55263 22086
rect 55862 22074 55875 22085
rect 55887 22074 55921 22086
rect 56520 22074 56533 22085
rect 56545 22074 56579 22086
rect 57178 22074 57191 22085
rect 57203 22074 57237 22086
rect 57836 22074 57849 22085
rect 57861 22074 57895 22086
rect 58494 22074 58507 22085
rect 58519 22074 58553 22133
rect 55215 20770 55263 22074
rect 55873 20770 55921 22074
rect 56531 20770 56579 22074
rect 55101 20160 55135 20671
rect 55215 20609 55249 20770
rect 55873 20758 55907 20770
rect 56531 20758 56565 20770
rect 55251 20643 55255 20745
rect 55279 20711 55283 20717
rect 55859 20711 55907 20758
rect 56517 20711 56565 20758
rect 55275 20677 55283 20711
rect 55291 20677 55907 20711
rect 55933 20677 55941 20711
rect 55949 20677 56565 20711
rect 55279 20671 55283 20677
rect 55861 20661 55907 20677
rect 56519 20661 56565 20677
rect 55873 20609 55907 20661
rect 56531 20609 56565 20661
rect 56567 20643 56571 20745
rect 57112 20717 57114 21814
rect 57140 20717 57142 21786
rect 57189 20770 57237 22074
rect 57847 20770 57895 22074
rect 57189 20758 57223 20770
rect 57847 20758 57881 20770
rect 56595 20711 56599 20717
rect 57175 20711 57223 20758
rect 57833 20711 57881 20758
rect 56591 20677 56599 20711
rect 56607 20677 57223 20711
rect 57249 20677 57257 20711
rect 57265 20677 57881 20711
rect 56595 20671 56599 20677
rect 57112 20664 57114 20671
rect 57140 20636 57142 20671
rect 57177 20661 57223 20677
rect 57835 20661 57881 20677
rect 57189 20609 57223 20661
rect 57847 20609 57881 20661
rect 57883 20643 57887 20745
rect 58434 20717 58436 21784
rect 58462 20717 58464 21756
rect 58505 20770 58553 22074
rect 58505 20758 58539 20770
rect 57911 20711 57915 20717
rect 58491 20711 58539 20758
rect 57907 20677 57915 20711
rect 57923 20677 58539 20711
rect 57911 20671 57915 20677
rect 58434 20664 58436 20671
rect 58462 20636 58464 20671
rect 58493 20661 58539 20677
rect 58505 20609 58539 20661
rect 58619 20671 58667 22173
rect 60172 20694 60220 22178
rect 60300 22188 60334 22240
rect 60916 22206 60954 22210
rect 60300 22100 60346 22188
rect 60916 22172 60956 22206
rect 60348 22138 60956 22172
rect 60924 22132 60928 22138
rect 60952 22104 60956 22138
rect 60958 22188 60992 22240
rect 60958 22100 61004 22188
rect 61574 22172 61612 22210
rect 61006 22138 61612 22172
rect 61616 22188 61650 22240
rect 62232 22206 62270 22210
rect 61616 22100 61662 22188
rect 62232 22172 62272 22206
rect 61664 22138 62272 22172
rect 62240 22132 62244 22138
rect 62268 22104 62272 22138
rect 62274 22188 62308 22240
rect 62274 22100 62320 22188
rect 62890 22172 62928 22210
rect 62322 22138 62928 22172
rect 62932 22188 62966 22240
rect 63548 22206 63586 22210
rect 62932 22100 62978 22188
rect 63548 22172 63588 22206
rect 62980 22138 63588 22172
rect 63556 22132 63560 22138
rect 63584 22104 63588 22138
rect 60300 22088 60334 22100
rect 60933 22088 60946 22099
rect 60958 22088 60992 22100
rect 61591 22088 61604 22099
rect 61616 22088 61650 22100
rect 62249 22088 62262 22099
rect 62274 22088 62308 22100
rect 62907 22088 62920 22099
rect 62932 22088 62966 22100
rect 63565 22088 63578 22099
rect 63590 22088 63624 22240
rect 63704 22178 63738 27058
rect 60286 20784 60334 22088
rect 55203 20575 58551 20609
rect 58619 20160 58653 20671
rect 60172 20160 60206 20694
rect 60286 20632 60320 20784
rect 60322 20666 60326 20768
rect 60872 20740 60880 21552
rect 60900 20740 60908 21524
rect 60944 20784 60992 22088
rect 61602 20784 61650 22088
rect 62260 20784 62308 22088
rect 62918 20784 62966 22088
rect 60944 20772 60978 20784
rect 61602 20772 61636 20784
rect 62260 20772 62294 20784
rect 62918 20772 62952 20784
rect 60350 20734 60354 20740
rect 60930 20734 60978 20772
rect 61588 20734 61636 20772
rect 60346 20700 60354 20734
rect 60362 20700 60978 20734
rect 61004 20700 61012 20734
rect 61020 20700 61636 20734
rect 60350 20694 60354 20700
rect 60872 20688 60880 20694
rect 60900 20660 60908 20694
rect 60932 20684 60978 20700
rect 61590 20684 61636 20700
rect 60944 20632 60978 20684
rect 61602 20632 61636 20684
rect 61638 20666 61642 20768
rect 61666 20734 61670 20740
rect 62246 20734 62294 20772
rect 62904 20734 62952 20772
rect 61662 20700 61670 20734
rect 61678 20700 62294 20734
rect 62320 20700 62328 20734
rect 62336 20700 62952 20734
rect 61666 20694 61670 20700
rect 62248 20684 62294 20700
rect 62906 20684 62952 20700
rect 62260 20632 62294 20684
rect 62918 20632 62952 20684
rect 62954 20666 62958 20768
rect 63500 20740 63506 21536
rect 63528 20740 63534 21508
rect 63576 20784 63624 22088
rect 63576 20772 63610 20784
rect 62982 20734 62986 20740
rect 63562 20734 63610 20772
rect 62978 20700 62986 20734
rect 62994 20700 63610 20734
rect 62982 20694 62986 20700
rect 63500 20682 63506 20694
rect 63528 20660 63534 20694
rect 63564 20684 63610 20700
rect 63576 20632 63610 20684
rect 63690 20694 63738 22178
rect 64017 22133 64617 22164
rect 64675 22133 65056 22164
rect 63937 21752 63960 22114
rect 63983 22099 65022 22130
rect 63965 21752 63988 22086
rect 64158 21906 64548 21940
rect 64158 21408 64192 21906
rect 64372 21838 64419 21885
rect 64334 21804 64419 21838
rect 64261 21745 64306 21756
rect 64389 21745 64434 21756
rect 64272 21569 64306 21745
rect 64400 21569 64434 21745
rect 64372 21510 64419 21557
rect 64334 21476 64419 21510
rect 64514 21408 64548 21906
rect 64158 21374 64548 21408
rect 64634 21906 65024 21940
rect 64634 21408 64668 21906
rect 64848 21838 64895 21885
rect 64810 21804 64895 21838
rect 64737 21745 64782 21756
rect 64865 21745 64910 21756
rect 64748 21569 64782 21745
rect 64876 21569 64910 21745
rect 64848 21510 64895 21557
rect 64810 21476 64895 21510
rect 64990 21408 65024 21906
rect 64634 21374 65024 21408
rect 60274 20598 63622 20632
rect 63690 20160 63724 20694
rect 63933 20622 63934 20708
rect 63971 20584 63972 20746
rect 64140 20704 64562 21324
rect 64616 20704 65038 21324
rect 37381 14445 37415 14454
rect 37376 14411 37449 14420
rect 37518 14030 38138 14452
rect 38284 14438 38658 14467
rect 38188 14404 38754 14438
rect 38188 14082 38222 14404
rect 38559 14324 38570 14335
rect 38243 14262 38324 14309
rect 38383 14290 38570 14324
rect 38571 14262 38652 14309
rect 38290 14224 38324 14262
rect 38618 14224 38652 14262
rect 38559 14196 38570 14207
rect 38383 14162 38570 14196
rect 38720 14082 38754 14404
rect 60944 14112 60978 20160
rect 73090 15268 73124 16594
rect 73170 15268 73178 15458
rect 73198 15302 73206 15486
rect 73198 15268 73228 15302
rect 64144 15234 64534 15268
rect 64144 14736 64178 15234
rect 64358 15166 64405 15213
rect 64320 15132 64405 15166
rect 64247 15073 64292 15084
rect 64375 15073 64420 15084
rect 64258 14897 64292 15073
rect 64386 14897 64420 15073
rect 64358 14838 64405 14885
rect 64320 14804 64405 14838
rect 64500 14736 64534 15234
rect 64144 14702 64534 14736
rect 64620 15234 65010 15268
rect 72996 15234 73290 15268
rect 64620 15206 64654 15234
rect 64620 14798 64688 15206
rect 64834 15166 64881 15213
rect 64796 15132 64881 15166
rect 64723 15073 64768 15084
rect 64851 15073 64896 15084
rect 64734 14897 64768 15073
rect 64862 14897 64896 15073
rect 64834 14838 64881 14885
rect 64796 14804 64881 14838
rect 64620 14736 64654 14798
rect 64976 14736 65010 15234
rect 73090 15200 73124 15234
rect 73090 15132 73148 15200
rect 73090 14872 73124 15132
rect 73142 14881 73158 15089
rect 73170 15085 73178 15234
rect 73198 15139 73206 15234
rect 73222 15139 73238 15234
rect 73170 15080 73182 15085
rect 73170 15073 73176 15080
rect 73166 14897 73176 15073
rect 73170 14881 73176 14897
rect 73192 14910 73242 15139
rect 73192 14885 73250 14910
rect 73090 14804 73148 14872
rect 73090 14770 73124 14804
rect 73150 14770 73154 14846
rect 73034 14750 73154 14770
rect 73090 14742 73124 14750
rect 73178 14742 73182 14874
rect 73028 14736 73182 14742
rect 73194 14736 73250 14885
rect 73256 14736 73290 15234
rect 64620 14702 65010 14736
rect 72996 14702 73290 14736
rect 73376 15234 73766 15268
rect 73376 14736 73410 15234
rect 73590 15166 73637 15213
rect 73552 15132 73637 15166
rect 73479 15073 73524 15084
rect 73607 15073 73652 15084
rect 73490 14897 73524 15073
rect 73618 14897 73652 15073
rect 73428 14736 73448 14884
rect 73590 14838 73637 14885
rect 73552 14804 73637 14838
rect 73732 14736 73766 15234
rect 73376 14702 73766 14736
rect 105810 15234 106200 15268
rect 105810 14736 105844 15234
rect 106024 15166 106071 15213
rect 105986 15132 106071 15166
rect 105913 15073 105958 15084
rect 106041 15073 106086 15084
rect 105924 14897 105958 15073
rect 106052 14897 106086 15073
rect 106024 14838 106071 14885
rect 105986 14804 106071 14838
rect 106166 14736 106200 15234
rect 105810 14702 106200 14736
rect 106286 15234 106676 15268
rect 106286 15206 106320 15234
rect 106286 14798 106354 15206
rect 106500 15166 106547 15213
rect 106462 15132 106547 15166
rect 106389 15073 106434 15084
rect 106517 15073 106562 15084
rect 106400 14897 106434 15073
rect 106528 14897 106562 15073
rect 106500 14838 106547 14885
rect 106462 14804 106547 14838
rect 106286 14736 106320 14798
rect 106642 14736 106676 15234
rect 114700 14750 114820 14770
rect 115006 14752 115246 15304
rect 115006 14750 115296 14752
rect 106286 14702 106676 14736
rect 114694 14722 114848 14742
rect 115006 14724 115246 14750
rect 115006 14722 115324 14724
rect 73090 14652 73124 14702
rect 73194 14700 73250 14702
rect 73130 14652 73250 14700
rect 115006 14666 115246 14722
rect 115635 14666 115722 15558
rect 38188 14048 38754 14082
rect 64126 14039 64548 14652
rect 64033 14005 64601 14039
rect 64602 14032 65024 14652
rect 73054 14288 73304 14652
rect 73358 14288 73780 14652
rect 73120 14238 73154 14248
rect 73508 14238 73542 14248
rect 73596 14238 73630 14248
rect 73136 14204 73188 14214
rect 73474 14204 73664 14214
rect 73102 14170 73126 14204
rect 73136 14136 73160 14204
rect 73234 14102 73268 14114
rect 73012 14068 73268 14102
rect 73394 14102 73428 14114
rect 73710 14102 73744 14114
rect 73394 14068 73744 14102
rect 105792 14039 106214 14652
rect 105699 14005 106267 14039
rect 106268 14032 106690 14652
rect 37398 13803 37415 13862
rect 37436 13775 37453 13824
rect 37518 13775 38138 13976
rect 38188 13928 38754 13962
rect 38188 13854 38222 13928
rect 38566 13878 38599 13882
rect 38720 13878 38754 13928
rect 73212 13890 73216 13980
rect 73240 13906 73244 13952
rect 38566 13859 38972 13878
rect 38559 13858 38972 13859
rect 38559 13854 38570 13858
rect 38188 13816 38228 13854
rect 38559 13850 38571 13854
rect 38720 13850 38754 13858
rect 38559 13848 38944 13850
rect 38243 13826 38324 13833
rect 38236 13816 38324 13826
rect 38178 13802 38186 13808
rect 38188 13796 38222 13816
rect 38243 13796 38324 13816
rect 38383 13830 38944 13848
rect 38383 13814 38570 13830
rect 38571 13796 38652 13830
rect 38720 13796 38754 13830
rect 38188 13775 38844 13796
rect 37436 13742 38138 13775
rect 38154 13742 40320 13775
rect 37436 13741 40320 13742
rect 37518 13591 38138 13741
rect 38188 13729 38844 13741
rect 38190 13722 38844 13729
rect 38208 13700 38228 13708
rect 38236 13706 38256 13708
rect 38367 13707 38575 13720
rect 38371 13695 38571 13707
rect 38188 13668 38222 13695
rect 38367 13686 38575 13695
rect 38371 13674 38571 13686
rect 38720 13668 38754 13695
rect 114148 13682 114160 13964
rect 114182 13716 114194 13938
rect 38333 13660 38609 13661
rect 38222 13627 38720 13660
rect 38222 13593 38720 13606
rect 25336 3874 25356 3932
rect 25364 3874 25384 3926
rect 25280 3634 25918 3874
rect 25336 3302 25338 3478
rect 25364 3330 25366 3450
rect 25144 2576 25344 2602
rect 25116 2548 25372 2574
rect 30942 1948 32294 1972
rect 43792 1052 43826 1854
rect 44450 1052 44484 1854
rect 43342 680 44522 1052
rect 30636 556 32641 584
rect 32687 556 32700 584
rect 40828 404 40886 434
rect 40862 370 40886 400
rect 43792 0 43826 680
rect 44450 0 44484 680
rect 26262 -542 30394 -540
rect 24381 -544 30394 -542
rect 24381 -615 30683 -544
rect 24381 -645 32600 -615
rect 920 -703 3348 -669
rect 844 -805 857 -771
rect 878 -782 891 -737
rect 974 -752 1537 -733
rect 1551 -752 2195 -733
rect 2209 -752 2853 -733
rect 2867 -752 3294 -733
rect 177 -1200 200 -1000
rect 205 -1228 228 -972
rect 177 -1600 200 -1400
rect 205 -1628 228 -1372
rect 177 -2000 200 -1800
rect 205 -2028 228 -1772
rect 177 -2400 200 -2200
rect 205 -2428 228 -2172
rect 930 -2510 954 -1158
rect 177 -2800 200 -2600
rect 205 -2828 228 -2572
rect 177 -3200 200 -3000
rect 205 -3228 228 -2972
rect 974 -3050 1008 -752
rect 2893 -782 2939 -765
rect 1112 -786 1499 -782
rect 1589 -786 2157 -782
rect 2247 -786 2815 -782
rect 2893 -786 3156 -782
rect 1100 -805 1515 -786
rect 1573 -805 2173 -786
rect 2231 -805 2831 -786
rect 2889 -805 3168 -786
rect 2893 -811 2970 -805
rect 2865 -820 2970 -814
rect 1134 -839 3134 -820
rect 1150 -843 3118 -839
rect 1489 -852 1599 -843
rect 2147 -852 2257 -843
rect 2805 -852 2915 -843
rect 1150 -854 3165 -852
rect 1515 -901 1573 -854
rect 2173 -901 2231 -854
rect 2831 -901 2889 -854
rect 1077 -913 1122 -902
rect 1088 -2889 1122 -913
rect 1527 -2901 1561 -901
rect 2185 -1696 2219 -901
rect 2164 -1832 2234 -1696
rect 1922 -1946 2336 -1832
rect 2164 -2152 2234 -1946
rect 2185 -2901 2219 -2152
rect 2843 -2901 2877 -901
rect 3135 -913 3180 -902
rect 3146 -2889 3180 -913
rect 1515 -2948 1574 -2901
rect 2173 -2948 2232 -2901
rect 2831 -2948 2890 -2901
rect 3118 -2948 3165 -2901
rect 1150 -2982 3165 -2948
rect 1515 -2998 1573 -2982
rect 2173 -2998 2231 -2982
rect 2831 -2998 2889 -2982
rect 1527 -3050 1561 -3016
rect 2185 -3050 2219 -3016
rect 2843 -3050 2877 -3016
rect 3260 -3050 3294 -752
rect 5168 -1890 5202 -760
rect 5282 -1890 5316 -1856
rect 5940 -1890 5974 -1856
rect 6598 -1890 6632 -1856
rect 7256 -1890 7290 -1856
rect 7914 -1890 7948 -1856
rect 8572 -1890 8606 -1856
rect 8686 -1890 8720 -760
rect 24381 -783 30683 -645
rect 32749 -651 32783 -635
rect 30719 -670 32749 -669
rect 30753 -703 32749 -670
rect 30685 -747 30787 -731
rect 30857 -747 31501 -733
rect 31515 -747 32159 -733
rect 32173 -747 32783 -733
rect 34008 -765 34040 -752
rect 34064 -765 34068 -724
rect 26648 -834 30008 -830
rect 30719 -834 30753 -765
rect 34306 -796 34307 -633
rect 36876 -664 36910 -236
rect 36990 -664 37024 -630
rect 37648 -664 37682 -630
rect 37762 -664 37796 -236
rect 38066 -664 38100 -236
rect 38180 -664 38214 -630
rect 38838 -664 38872 -630
rect 38952 -664 38986 -236
rect 35886 -698 39246 -664
rect 36876 -794 36910 -698
rect 37642 -728 37644 -724
rect 36978 -794 37230 -728
rect 37244 -766 37694 -728
rect 37282 -794 37694 -766
rect 37762 -794 37796 -698
rect 38066 -794 38100 -698
rect 38168 -794 38546 -728
rect 38560 -766 38884 -728
rect 38598 -794 38884 -766
rect 38952 -794 38986 -698
rect 39376 -794 39396 -610
rect 40262 -794 40296 -776
rect 34008 -830 34040 -811
rect 34064 -830 34068 -811
rect 26648 -864 31892 -834
rect 29094 -868 31892 -864
rect 28998 -916 29009 -905
rect 29021 -916 29032 -905
rect 28998 -932 29032 -916
rect 28998 -936 29270 -932
rect 29360 -936 29928 -932
rect 30070 -936 30104 -898
rect 23548 -1370 23910 -962
rect 28998 -966 30104 -936
rect 28688 -1006 28720 -972
rect 28688 -1024 28714 -1006
rect 28744 -1024 28748 -972
rect 23374 -1516 23910 -1370
rect 25434 -1516 25684 -1370
rect 4666 -1924 9794 -1890
rect 5168 -2378 5202 -1924
rect 5282 -1961 5320 -1954
rect 5270 -1976 5320 -1961
rect 5940 -1976 5978 -1954
rect 6598 -1976 6636 -1954
rect 7256 -1976 7294 -1954
rect 7914 -1976 7952 -1954
rect 8572 -1961 8610 -1954
rect 8572 -1976 8618 -1961
rect 5270 -1992 5328 -1976
rect 5928 -1992 5986 -1976
rect 6586 -1992 6644 -1976
rect 7244 -1992 7302 -1976
rect 7902 -1992 7960 -1976
rect 8524 -1986 8544 -1978
rect 8560 -1992 8618 -1976
rect 5270 -2026 8618 -1992
rect 5270 -2064 5328 -2026
rect 5928 -2064 5986 -2026
rect 6586 -2064 6644 -2026
rect 7244 -2064 7302 -2026
rect 7902 -2064 7960 -2026
rect 4616 -2392 5230 -2378
rect 5168 -2406 5202 -2392
rect 4644 -2448 5230 -2406
rect 5168 -3004 5202 -2448
rect 5282 -2864 5316 -2064
rect 5940 -2864 5974 -2064
rect 6598 -2864 6632 -2064
rect 7256 -2864 7290 -2064
rect 7914 -2864 7948 -2064
rect 8524 -2534 8544 -2032
rect 8560 -2064 8618 -2026
rect 8572 -2864 8606 -2064
rect 5270 -2902 5328 -2864
rect 5928 -2902 5986 -2864
rect 6586 -2902 6644 -2864
rect 7244 -2902 7302 -2864
rect 7902 -2902 7960 -2864
rect 8560 -2902 8618 -2864
rect 5270 -2936 8618 -2902
rect 5270 -2952 5328 -2936
rect 5928 -2952 5986 -2936
rect 6586 -2952 6644 -2936
rect 7244 -2952 7302 -2936
rect 7902 -2952 7960 -2936
rect 8560 -2952 8618 -2936
rect 5270 -2967 5285 -2952
rect 8603 -2967 8618 -2952
rect 5282 -3004 5316 -2970
rect 5940 -3004 5974 -2970
rect 6598 -3004 6632 -2970
rect 7256 -3004 7290 -2970
rect 7914 -3004 7948 -2970
rect 8572 -3004 8606 -2970
rect 8686 -3004 8720 -1924
rect 22518 -2010 22540 -1770
rect 23548 -2018 23910 -1516
rect 25498 -1630 25652 -1516
rect 24512 -2010 24628 -1988
rect 24556 -2015 24602 -2010
rect 25214 -2015 25260 -1988
rect 25850 -2004 25944 -1988
rect 25852 -2012 25942 -2004
rect 25872 -2015 25918 -2012
rect 24484 -2038 24656 -2016
rect 24528 -2043 24630 -2038
rect 25186 -2043 25288 -2016
rect 25822 -2032 25972 -2016
rect 25824 -2040 25970 -2032
rect 25844 -2043 25946 -2040
rect 27982 -2230 28016 -1025
rect 28616 -1190 28714 -1024
rect 28616 -1204 28694 -1190
rect 28614 -1374 28782 -1204
rect 28022 -1832 28642 -1410
rect 28658 -1848 28674 -1390
rect 28998 -1424 29032 -966
rect 29174 -970 29742 -966
rect 29832 -970 30104 -966
rect 29286 -1017 29344 -1013
rect 29944 -1017 30002 -1013
rect 29101 -1029 29146 -1018
rect 29287 -1025 29332 -1017
rect 29112 -1424 29146 -1029
rect 28692 -1458 29258 -1424
rect 28692 -1780 28726 -1458
rect 28998 -1538 29032 -1458
rect 29112 -1521 29146 -1458
rect 29224 -1517 29258 -1458
rect 29298 -1426 29332 -1025
rect 29759 -1029 29804 -1018
rect 29945 -1025 29990 -1017
rect 29298 -1517 29343 -1426
rect 29770 -1505 29804 -1029
rect 29956 -1517 29990 -1025
rect 29063 -1538 29074 -1527
rect 28747 -1600 28828 -1553
rect 28887 -1572 29074 -1538
rect 28794 -1638 28828 -1600
rect 28998 -1666 29032 -1572
rect 29075 -1600 29156 -1553
rect 29224 -1564 29448 -1517
rect 29742 -1564 29789 -1517
rect 29944 -1564 30002 -1517
rect 29158 -1598 29789 -1564
rect 29832 -1598 30002 -1564
rect 29122 -1654 29156 -1600
rect 29063 -1666 29074 -1655
rect 29224 -1666 29258 -1598
rect 29286 -1614 29344 -1598
rect 29944 -1614 30002 -1598
rect 29298 -1666 29332 -1614
rect 29987 -1629 30002 -1614
rect 30070 -1666 30104 -970
rect 30464 -1370 30468 -1017
rect 30719 -1308 30753 -868
rect 30833 -905 30880 -889
rect 30821 -936 30880 -905
rect 31058 -936 31105 -889
rect 31491 -920 31538 -889
rect 31479 -936 31538 -920
rect 31716 -936 31763 -889
rect 30821 -970 31105 -936
rect 31148 -970 31763 -936
rect 30821 -1017 30879 -970
rect 31479 -1017 31537 -970
rect 30719 -1336 30778 -1308
rect 30410 -1380 30420 -1370
rect 30406 -1510 30420 -1380
rect 30410 -1512 30420 -1510
rect 30464 -1380 30482 -1370
rect 30464 -1510 30486 -1380
rect 30464 -1512 30482 -1510
rect 30464 -1517 30468 -1512
rect 30719 -1666 30753 -1336
rect 30833 -1517 30867 -1017
rect 31075 -1029 31120 -1018
rect 31086 -1505 31120 -1029
rect 31491 -1274 31525 -1017
rect 31733 -1029 31778 -1018
rect 31292 -1336 31588 -1274
rect 31491 -1517 31525 -1336
rect 31744 -1380 31778 -1029
rect 31734 -1450 31786 -1380
rect 31618 -1506 31786 -1450
rect 31618 -1517 31754 -1506
rect 30821 -1564 30880 -1517
rect 31058 -1564 31105 -1517
rect 31479 -1564 31538 -1517
rect 31618 -1564 31763 -1517
rect 30821 -1598 31105 -1564
rect 31148 -1598 31763 -1564
rect 30821 -1614 30879 -1598
rect 31479 -1614 31537 -1598
rect 30821 -1629 30836 -1614
rect 31554 -1642 31576 -1604
rect 31582 -1614 31604 -1604
rect 31858 -1666 31892 -868
rect 28887 -1700 31892 -1666
rect 32510 -841 32806 -830
rect 32841 -841 33464 -830
rect 32510 -852 32795 -841
rect 32841 -852 33453 -841
rect 33499 -852 34088 -830
rect 32510 -864 34088 -852
rect 29224 -1780 29258 -1700
rect 28692 -1814 29258 -1780
rect 28560 -1962 28568 -1932
rect 28588 -1962 28596 -1960
rect 28716 -2162 28732 -1962
rect 28744 -2190 28760 -1934
rect 29298 -2230 29332 -1700
rect 30070 -2230 30104 -1700
rect 30719 -2230 30753 -1700
rect 32510 -2162 32544 -864
rect 32746 -932 33852 -885
rect 33912 -932 33959 -885
rect 32686 -966 33301 -932
rect 33344 -966 33959 -932
rect 32613 -1025 32658 -1014
rect 32624 -2001 32658 -1025
rect 32666 -2014 32718 -972
rect 32722 -2014 32746 -972
rect 32795 -1013 32853 -966
rect 33453 -1013 33511 -966
rect 32807 -2013 32841 -1013
rect 33271 -1025 33316 -1014
rect 33282 -2001 33316 -1025
rect 33465 -2013 33499 -1013
rect 33929 -1025 33974 -1014
rect 33940 -2001 33974 -1025
rect 32795 -2060 32854 -2013
rect 33254 -2060 33301 -2013
rect 33453 -2060 33512 -2013
rect 33912 -2060 33959 -2013
rect 34008 -2014 34040 -864
rect 34054 -926 34088 -864
rect 34054 -2014 34096 -926
rect 34560 -1210 34561 -796
rect 35344 -1196 35362 -1020
rect 35754 -1210 36210 -796
rect 34214 -1234 36210 -1210
rect 32686 -2094 33301 -2060
rect 33344 -2094 33959 -2060
rect 32795 -2110 32853 -2094
rect 33453 -2110 33511 -2094
rect 34008 -2162 34040 -2152
rect 34054 -2162 34088 -2014
rect 32510 -2196 34088 -2162
rect 24412 -2234 26062 -2230
rect 17792 -2902 20074 -2506
rect 14894 -2936 20074 -2902
rect 4666 -3038 9794 -3004
rect 974 -3084 3294 -3050
rect 914 -3348 3685 -3312
rect 5168 -3348 5202 -3038
rect 5282 -3348 5316 -3314
rect 5940 -3348 5974 -3314
rect 6598 -3348 6632 -3314
rect 7256 -3348 7290 -3314
rect 7914 -3348 7948 -3314
rect 8572 -3348 8606 -3314
rect 8686 -3348 8720 -3038
rect 17792 -3074 20074 -2936
rect 17792 -3348 20100 -3312
rect 177 -3600 200 -3400
rect 205 -3628 228 -3372
rect 914 -3382 20100 -3348
rect 914 -4034 3685 -3382
rect 5168 -3462 5202 -3382
rect 5282 -3462 5316 -3382
rect 5940 -3462 5974 -3382
rect 6598 -3462 6632 -3382
rect 7256 -3462 7290 -3382
rect 7914 -3462 7948 -3382
rect 8572 -3462 8606 -3382
rect 8686 -3462 8720 -3382
rect 11250 -3444 11298 -3428
rect 5168 -3496 8720 -3462
rect 5168 -3920 5202 -3496
rect 5282 -3920 5316 -3496
rect 5328 -3508 5329 -3507
rect 5927 -3508 5928 -3507
rect 5327 -3509 5328 -3508
rect 5928 -3509 5929 -3508
rect 5327 -3908 5328 -3907
rect 5928 -3908 5929 -3907
rect 5328 -3909 5329 -3908
rect 5927 -3909 5928 -3908
rect 5940 -3920 5974 -3496
rect 5986 -3508 5987 -3507
rect 6585 -3508 6586 -3507
rect 5985 -3509 5986 -3508
rect 6586 -3509 6587 -3508
rect 5985 -3908 5986 -3907
rect 6586 -3908 6587 -3907
rect 5986 -3909 5987 -3908
rect 6585 -3909 6586 -3908
rect 6598 -3920 6632 -3496
rect 6644 -3508 6645 -3507
rect 7243 -3508 7244 -3507
rect 6643 -3509 6644 -3508
rect 7244 -3509 7245 -3508
rect 6643 -3908 6644 -3907
rect 7244 -3908 7245 -3907
rect 6644 -3909 6645 -3908
rect 7243 -3909 7244 -3908
rect 7256 -3920 7290 -3496
rect 7302 -3508 7303 -3507
rect 7901 -3508 7902 -3507
rect 7301 -3509 7302 -3508
rect 7902 -3509 7903 -3508
rect 7301 -3908 7302 -3907
rect 7902 -3908 7903 -3907
rect 7302 -3909 7303 -3908
rect 7901 -3909 7902 -3908
rect 7914 -3920 7948 -3496
rect 7960 -3508 7961 -3507
rect 8559 -3508 8560 -3507
rect 7959 -3509 7960 -3508
rect 8560 -3509 8561 -3508
rect 7959 -3908 7960 -3907
rect 8560 -3908 8561 -3907
rect 7960 -3909 7961 -3908
rect 8559 -3909 8560 -3908
rect 8572 -3920 8606 -3496
rect 8686 -3920 8720 -3496
rect 5168 -3954 8720 -3920
rect 11098 -3477 11124 -3450
rect 11250 -3462 11264 -3444
rect 11272 -3462 11298 -3450
rect 11128 -3477 11132 -3474
rect 11098 -3919 11132 -3477
rect 11264 -3477 11268 -3474
rect 11272 -3477 11318 -3462
rect 11264 -3496 11318 -3477
rect 11162 -3908 11196 -3508
rect 11200 -3908 11234 -3508
rect 11264 -3886 11298 -3496
rect 11098 -3942 11124 -3919
rect 11128 -3942 11132 -3919
rect 11250 -3919 11298 -3886
rect 11250 -3920 11268 -3919
rect 11264 -3942 11268 -3920
rect 11272 -3920 11298 -3919
rect 11010 -3954 11124 -3942
rect 5168 -4034 5202 -3954
rect 5282 -4034 5316 -3954
rect 5940 -4034 5974 -3954
rect 6598 -4034 6632 -3954
rect 7256 -4034 7290 -3954
rect 7914 -4034 7948 -3954
rect 8572 -4034 8606 -3954
rect 8686 -4034 8720 -3954
rect 11098 -3966 11124 -3954
rect 11272 -3954 11318 -3920
rect 17792 -3944 20100 -3382
rect 20370 -3938 21482 -3312
rect 11272 -3966 11298 -3954
rect 11044 -3988 11098 -3976
rect 914 -4068 20160 -4034
rect 20298 -4068 21326 -4066
rect 914 -4104 3685 -4068
rect 5168 -8916 5202 -4068
rect 8686 -8916 8720 -4068
rect 24440 -4108 24474 -2362
rect 26516 -2506 30140 -2230
rect 30683 -2500 32824 -2230
rect 26516 -3944 30248 -2506
rect 30518 -2624 32824 -2500
rect 30518 -2952 32841 -2624
rect 32848 -2914 32879 -2662
rect 30518 -3938 32824 -2952
rect 22776 -4142 26232 -4108
rect 24440 -4210 24474 -4142
rect 24542 -4210 24576 -4142
rect 24740 -4210 24778 -4172
rect 25398 -4210 25436 -4172
rect 26056 -4210 26094 -4172
rect 24440 -4244 24778 -4210
rect 24830 -4244 25436 -4210
rect 25488 -4244 26094 -4210
rect 22788 -4288 22834 -4282
rect 22788 -4294 22860 -4288
rect 22794 -4306 22860 -4294
rect 22828 -4694 22860 -4306
rect 22828 -5798 22834 -4694
rect 22884 -4722 22888 -4260
rect 24104 -4294 24150 -4282
rect 24104 -4306 24144 -4294
rect 23512 -5742 23526 -5496
rect 23540 -5798 23582 -5496
rect 24104 -5542 24128 -4634
rect 24440 -5784 24474 -4244
rect 24542 -4326 24576 -4244
rect 24734 -4270 24836 -4254
rect 25392 -4260 25494 -4254
rect 25362 -4270 25520 -4260
rect 26050 -4270 26152 -4254
rect 24614 -4282 24615 -4281
rect 24613 -4283 24614 -4282
rect 24762 -4283 24808 -4282
rect 25420 -4283 25466 -4282
rect 26078 -4283 26124 -4282
rect 24757 -4294 24808 -4283
rect 25415 -4288 25466 -4283
rect 24762 -4298 24808 -4294
rect 25390 -4298 25492 -4288
rect 26073 -4294 26124 -4283
rect 26078 -4298 26124 -4294
rect 24756 -4342 24757 -4341
rect 24755 -4343 24756 -4342
rect 24768 -4354 24802 -4298
rect 24813 -4342 24814 -4341
rect 25414 -4342 25415 -4341
rect 24814 -4343 24815 -4342
rect 25413 -4343 25414 -4342
rect 25426 -4354 25460 -4298
rect 25471 -4342 25472 -4341
rect 26072 -4342 26073 -4341
rect 25472 -4343 25473 -4342
rect 26071 -4343 26072 -4342
rect 26084 -4354 26118 -4298
rect 26198 -4354 26232 -4142
rect 24504 -4416 24576 -4378
rect 24626 -4388 26232 -4354
rect 24755 -4400 24756 -4399
rect 24756 -4401 24757 -4400
rect 24542 -4984 24576 -4416
rect 24756 -5000 24757 -4999
rect 24755 -5001 24756 -5000
rect 24768 -5012 24802 -4388
rect 24814 -4400 24815 -4399
rect 25413 -4400 25414 -4399
rect 24813 -4401 24814 -4400
rect 25414 -4401 25415 -4400
rect 24813 -5000 24814 -4999
rect 25414 -5000 25415 -4999
rect 24814 -5001 24815 -5000
rect 25413 -5001 25414 -5000
rect 25426 -5012 25460 -4388
rect 25472 -4400 25473 -4399
rect 26071 -4400 26072 -4399
rect 25471 -4401 25472 -4400
rect 26072 -4401 26073 -4400
rect 25471 -5000 25472 -4999
rect 26072 -5000 26073 -4999
rect 25472 -5001 25473 -5000
rect 26071 -5001 26072 -5000
rect 26084 -5012 26118 -4388
rect 26198 -5012 26232 -4388
rect 24504 -5074 24576 -5036
rect 24626 -5046 26232 -5012
rect 24755 -5058 24756 -5057
rect 24756 -5059 24757 -5058
rect 24542 -5642 24576 -5074
rect 24756 -5658 24757 -5657
rect 24755 -5659 24756 -5658
rect 24768 -5670 24802 -5046
rect 24814 -5058 24815 -5057
rect 25413 -5058 25414 -5057
rect 24813 -5059 24814 -5058
rect 25414 -5059 25415 -5058
rect 24813 -5658 24814 -5657
rect 25414 -5658 25415 -5657
rect 24814 -5659 24815 -5658
rect 25413 -5659 25414 -5658
rect 25426 -5670 25460 -5046
rect 25472 -5058 25473 -5057
rect 26071 -5058 26072 -5057
rect 25471 -5059 25472 -5058
rect 26072 -5059 26073 -5058
rect 25471 -5658 25472 -5657
rect 26072 -5658 26073 -5657
rect 25472 -5659 25473 -5658
rect 26071 -5659 26072 -5658
rect 26084 -5670 26118 -5046
rect 26198 -5670 26232 -5046
rect 26516 -5232 30140 -3944
rect 30683 -4072 32824 -3938
rect 34008 -4072 34040 -2196
rect 34064 -4072 34068 -2196
rect 34560 -2234 34561 -1234
rect 35754 -2234 36210 -1234
rect 30683 -4108 34307 -4072
rect 35790 -4108 35824 -2234
rect 36562 -2670 36596 -850
rect 36632 -2518 36654 -1414
rect 36664 -1462 40296 -794
rect 40688 -1110 40698 -752
rect 40831 -771 41500 -633
rect 41518 -765 41546 -752
rect 41574 -765 41602 -752
rect 41668 -771 44931 -633
rect 45074 -706 45098 400
rect 45108 -740 45132 434
rect 40831 -805 44931 -771
rect 40688 -1324 40716 -1110
rect 40688 -1330 40698 -1324
rect 36664 -1532 40288 -1462
rect 36562 -2700 36602 -2670
rect 36664 -2682 39378 -1532
rect 39440 -1714 39444 -1532
rect 40218 -1714 40252 -1532
rect 40831 -1540 41500 -805
rect 40867 -1714 40901 -1540
rect 40981 -1714 41015 -1680
rect 41343 -1714 41377 -1540
rect 41457 -1714 41491 -1540
rect 41518 -1714 41546 -811
rect 41574 -1464 41602 -811
rect 41668 -853 44931 -805
rect 41628 -864 44931 -853
rect 41639 -1544 44931 -864
rect 45102 -1334 45104 -752
rect 41639 -1652 41673 -1544
rect 41639 -1714 41684 -1652
rect 36628 -2698 39378 -2682
rect 36622 -2700 39378 -2698
rect 30683 -4120 36380 -4108
rect 30500 -4142 36380 -4120
rect 30500 -4154 34307 -4142
rect 30500 -4354 30534 -4154
rect 30683 -4222 34307 -4154
rect 30676 -4256 34307 -4222
rect 30580 -4270 30682 -4266
rect 30608 -4295 30654 -4294
rect 30603 -4298 30654 -4295
rect 30603 -4306 30648 -4298
rect 30614 -4354 30648 -4306
rect 30652 -4348 30670 -4298
rect 30683 -4354 34307 -4256
rect 30466 -4388 34307 -4354
rect 30500 -5012 30534 -4388
rect 30614 -5012 30648 -4388
rect 30652 -4486 30670 -4394
rect 30652 -5006 30654 -4934
rect 30659 -5000 30660 -4999
rect 30660 -5001 30661 -5000
rect 30683 -5012 34307 -4388
rect 34912 -4796 35374 -4158
rect 35598 -4184 35670 -4172
rect 35636 -4222 35708 -4210
rect 35536 -4382 35564 -4250
rect 35538 -4586 35564 -4578
rect 30466 -5046 34307 -5012
rect 28000 -5442 28034 -5232
rect 28114 -5290 28148 -5232
rect 28772 -5290 28806 -5232
rect 28744 -5340 28782 -5302
rect 28176 -5374 28782 -5340
rect 28886 -5442 28920 -5232
rect 28000 -5476 28920 -5442
rect 29190 -5442 29224 -5232
rect 29304 -5290 29338 -5232
rect 29962 -5290 29996 -5232
rect 29934 -5340 29972 -5302
rect 29366 -5374 29972 -5340
rect 30076 -5442 30110 -5232
rect 29190 -5476 30110 -5442
rect 29362 -5586 29912 -5584
rect 29390 -5614 29884 -5612
rect 30500 -5670 30534 -5046
rect 30614 -5670 30648 -5046
rect 30652 -5138 30654 -5052
rect 30660 -5058 30661 -5057
rect 30659 -5059 30660 -5058
rect 30652 -5664 30654 -5586
rect 30659 -5658 30660 -5657
rect 30660 -5659 30661 -5658
rect 30683 -5670 34307 -5046
rect 24626 -5704 34307 -5670
rect 24768 -5784 24802 -5704
rect 25426 -5784 25460 -5704
rect 26084 -5784 26118 -5704
rect 26198 -5784 26232 -5704
rect 30500 -5784 30534 -5704
rect 30614 -5784 30648 -5704
rect 30652 -5784 30654 -5710
rect 30683 -5784 34307 -5704
rect 24440 -5818 34307 -5784
rect 20268 -6684 20292 -5990
rect 20302 -6684 20326 -6024
rect 25342 -6202 25360 -5818
rect 25398 -6202 25416 -5870
rect 24582 -6290 25130 -6256
rect 24582 -6572 24616 -6290
rect 24768 -6370 24802 -6290
rect 24944 -6370 24955 -6359
rect 24646 -6414 24718 -6376
rect 24684 -6448 24718 -6414
rect 24768 -6404 24955 -6370
rect 24755 -6416 24756 -6415
rect 24756 -6417 24757 -6416
rect 24756 -6446 24757 -6445
rect 24755 -6447 24756 -6446
rect 24768 -6458 24802 -6404
rect 24956 -6414 25028 -6376
rect 24814 -6416 24815 -6415
rect 24813 -6417 24814 -6416
rect 24813 -6446 24814 -6445
rect 24814 -6447 24815 -6446
rect 24944 -6458 24955 -6447
rect 24994 -6448 25028 -6414
rect 24768 -6492 24955 -6458
rect 24768 -6572 24802 -6492
rect 25096 -6572 25130 -6290
rect 24582 -6606 25130 -6572
rect 25180 -6664 25818 -6202
rect 25342 -6678 25360 -6664
rect 25398 -6678 25416 -6664
rect 24582 -6766 25130 -6732
rect 24582 -7048 24616 -6766
rect 24768 -6846 24802 -6766
rect 24944 -6846 24955 -6835
rect 24646 -6886 24718 -6852
rect 24768 -6880 24955 -6846
rect 24646 -6890 24726 -6886
rect 24684 -6924 24726 -6890
rect 24755 -6892 24756 -6891
rect 24756 -6893 24757 -6892
rect 24756 -6922 24757 -6921
rect 24755 -6923 24756 -6922
rect 24700 -6940 24726 -6924
rect 24756 -6942 24762 -6928
rect 24768 -6934 24802 -6880
rect 24956 -6890 25028 -6852
rect 24814 -6892 24815 -6891
rect 24813 -6893 24814 -6892
rect 24813 -6922 24814 -6921
rect 24814 -6923 24815 -6922
rect 24808 -6934 24862 -6928
rect 24944 -6934 24955 -6923
rect 24994 -6924 25028 -6890
rect 24768 -6968 24955 -6934
rect 24768 -7048 24802 -6968
rect 25096 -7048 25130 -6766
rect 24582 -7082 25130 -7048
rect 25180 -7140 25818 -6678
rect 26078 -6868 26080 -5854
rect 26198 -7560 26232 -5818
rect 30500 -5972 30534 -5818
rect 30652 -5894 30654 -5818
rect 30683 -5854 34307 -5818
rect 30683 -6104 31456 -5854
rect 9274 -8188 9394 -8168
rect 9580 -8186 9820 -7634
rect 9580 -8188 9870 -8186
rect 9268 -8216 9422 -8196
rect 9580 -8214 9820 -8188
rect 9580 -8216 9898 -8214
rect 9580 -8272 9820 -8216
rect 30833 -8840 30867 -6104
rect 31457 -7612 31462 -6024
rect 31491 -7612 31496 -5990
rect 31632 -6096 32624 -5854
rect 32149 -8840 32183 -6096
rect 32792 -6774 34307 -5854
rect 34916 -6146 34950 -4796
rect 34970 -4880 35320 -4846
rect 34970 -5354 35004 -4880
rect 35090 -4948 35200 -4910
rect 35128 -4982 35200 -4948
rect 35073 -5032 35129 -5021
rect 35161 -5032 35217 -5021
rect 35084 -5208 35129 -5032
rect 35172 -5208 35217 -5032
rect 35090 -5258 35200 -5220
rect 35128 -5292 35200 -5258
rect 34966 -5360 35004 -5354
rect 35286 -5360 35320 -4880
rect 34966 -5394 35320 -5360
rect 34966 -5572 34984 -5394
rect 34916 -6376 34956 -6146
rect 34964 -6374 34984 -6174
rect 35484 -6376 35508 -5572
rect 35540 -5812 35564 -5572
rect 35574 -6376 35608 -4294
rect 35618 -4586 35640 -4578
rect 35790 -6376 35824 -4142
rect 35892 -4210 36128 -4172
rect 36204 -4210 36242 -4172
rect 35892 -4244 36242 -4210
rect 35892 -4282 35950 -4244
rect 35904 -6376 35949 -4282
rect 36221 -4294 36266 -4283
rect 34916 -6398 36046 -6376
rect 34916 -6402 36006 -6398
rect 34916 -6774 34950 -6402
rect 35484 -6596 35508 -6402
rect 35574 -6774 35608 -6402
rect 35790 -6774 35824 -6402
rect 35904 -6774 35949 -6402
rect 36232 -6596 36266 -4294
rect 36232 -6774 36277 -6596
rect 36346 -6774 36380 -4142
rect 36562 -6774 36596 -2700
rect 36628 -2808 39378 -2700
rect 36628 -2938 36634 -2808
rect 36664 -3916 39378 -2808
rect 39430 -1748 41684 -1714
rect 39430 -1848 39464 -1748
rect 40104 -1800 40150 -1769
rect 40092 -1816 40150 -1800
rect 39482 -1848 39486 -1841
rect 39430 -1904 39486 -1848
rect 39606 -1850 40150 -1816
rect 40184 -1850 40190 -1816
rect 40092 -1897 40150 -1850
rect 40218 -1875 40252 -1748
rect 40833 -1850 40848 -1816
rect 39430 -3046 39464 -1904
rect 39480 -2228 39486 -1904
rect 39508 -2200 39514 -1904
rect 39533 -1909 39578 -1898
rect 39482 -2953 39486 -2228
rect 39544 -2885 39578 -1909
rect 39684 -2434 39876 -2382
rect 40104 -2434 40138 -1897
rect 39660 -2502 40138 -2434
rect 40104 -2897 40138 -2502
rect 40140 -2682 40172 -2318
rect 40196 -2682 40200 -1897
rect 40140 -2892 40200 -2682
rect 40218 -2851 40270 -1875
rect 40202 -2885 40270 -2851
rect 40140 -2897 40172 -2892
rect 40196 -2897 40200 -2892
rect 40092 -2944 40172 -2897
rect 39606 -2978 40150 -2944
rect 40092 -2994 40172 -2978
rect 40106 -3009 40172 -2994
rect 40106 -3046 40138 -3009
rect 40140 -3046 40172 -3009
rect 40218 -3046 40252 -2885
rect 40867 -3046 40901 -1748
rect 40981 -1785 41028 -1769
rect 40969 -1816 41028 -1785
rect 41343 -1816 41377 -1748
rect 41457 -1769 41491 -1748
rect 41457 -1782 41504 -1769
rect 41518 -1782 41546 -1748
rect 41457 -1800 41546 -1782
rect 41445 -1816 41546 -1800
rect 40906 -1850 40939 -1816
rect 40969 -1850 41546 -1816
rect 40969 -1897 41027 -1850
rect 40981 -2318 41015 -1897
rect 40981 -2897 41026 -2318
rect 41343 -2897 41377 -1850
rect 41445 -1897 41503 -1850
rect 41518 -1897 41546 -1850
rect 41632 -1776 41684 -1748
rect 41457 -2318 41491 -1897
rect 41518 -1898 41558 -1897
rect 41507 -1909 41558 -1898
rect 41518 -2318 41558 -1909
rect 41457 -2897 41502 -2318
rect 41518 -2885 41563 -2318
rect 41574 -2688 41586 -1869
rect 41518 -2897 41558 -2892
rect 40969 -2910 41504 -2897
rect 41518 -2910 41546 -2897
rect 40922 -2978 40939 -2944
rect 40969 -2978 41546 -2910
rect 41574 -2925 41586 -2892
rect 41632 -2973 41700 -1776
rect 40969 -2994 41027 -2978
rect 40969 -3009 40984 -2994
rect 40981 -3046 41015 -3012
rect 41343 -3046 41377 -2978
rect 41445 -2994 41503 -2978
rect 41457 -3046 41502 -2994
rect 41518 -3046 41546 -2978
rect 41628 -2984 41700 -2973
rect 42115 -2318 42149 -1544
rect 41632 -3046 41684 -2984
rect 39430 -3080 41684 -3046
rect 39440 -3916 39444 -3080
rect 40106 -3528 40138 -3080
rect 40140 -3494 40172 -3080
rect 40218 -3916 40252 -3080
rect 40867 -3626 40901 -3080
rect 36664 -3950 40320 -3916
rect 36664 -4018 39378 -3950
rect 39440 -4002 39444 -3950
rect 39446 -4002 39493 -3971
rect 39434 -4018 39493 -4002
rect 39934 -4018 39981 -3971
rect 40104 -4002 40150 -3971
rect 40092 -4018 40150 -4002
rect 36664 -4052 39981 -4018
rect 40024 -4052 40150 -4018
rect 36664 -4058 39378 -4052
rect 39434 -4058 39492 -4052
rect 40092 -4058 40150 -4052
rect 36664 -4640 39388 -4058
rect 39396 -4099 39492 -4058
rect 39396 -4599 39444 -4099
rect 39446 -4599 39480 -4099
rect 39951 -4111 39996 -4100
rect 39962 -4587 39996 -4111
rect 39396 -4640 39493 -4599
rect 36664 -4646 39378 -4640
rect 39434 -4646 39493 -4640
rect 39934 -4646 39981 -4599
rect 40024 -4640 40038 -4058
rect 40052 -4099 40150 -4058
rect 40052 -4599 40094 -4099
rect 40104 -4599 40138 -4099
rect 40218 -4280 40252 -3950
rect 40168 -4308 40344 -4280
rect 40168 -4326 40288 -4308
rect 40168 -4342 40344 -4326
rect 40052 -4640 40150 -4599
rect 40092 -4646 40150 -4640
rect 36664 -4680 39981 -4646
rect 40024 -4680 40150 -4646
rect 36664 -4748 39378 -4680
rect 39434 -4696 39492 -4680
rect 40092 -4696 40150 -4680
rect 39440 -4748 39444 -4696
rect 40135 -4711 40150 -4696
rect 40218 -4748 40252 -4342
rect 40288 -4344 40344 -4342
rect 36664 -4782 40320 -4748
rect 36664 -5232 39378 -4782
rect 39440 -4800 39444 -4782
rect 39418 -5008 39444 -4800
rect 39440 -5013 39444 -5008
rect 40218 -5100 40252 -4782
rect 40831 -4818 41058 -3626
rect 32792 -7668 36852 -6774
rect 32792 -7692 34307 -7668
rect 35790 -8916 35824 -7668
rect 35904 -8826 35938 -7668
rect 36562 -8826 36596 -7668
rect 37178 -7816 37192 -7134
rect 40867 -7380 40901 -4818
rect 39896 -8188 40016 -8168
rect 40202 -8186 40442 -7634
rect 40202 -8188 40492 -8186
rect 39890 -8216 40044 -8196
rect 40202 -8214 40442 -8188
rect 40202 -8216 40520 -8214
rect 40202 -8272 40442 -8216
rect 40831 -8272 40918 -7380
rect 40867 -8939 40901 -8272
rect 41343 -8899 41377 -3080
rect 41457 -3386 41502 -3080
rect 41448 -3420 41502 -3386
rect 41518 -3420 41546 -3080
rect 41639 -3420 41684 -3080
rect 42115 -3420 42160 -2318
rect 42176 -3420 42204 -1544
rect 42232 -3420 42260 -1544
rect 42297 -2318 42331 -1544
rect 42297 -3420 42342 -2318
rect 42773 -3420 42807 -1544
rect 42838 -3420 42866 -1544
rect 42894 -3420 42922 -1544
rect 42955 -3420 42989 -1544
rect 41386 -3454 42989 -3420
rect 41386 -4752 41420 -3454
rect 41457 -3460 41502 -3454
rect 41518 -3460 41546 -3454
rect 41457 -3475 41546 -3460
rect 41639 -3475 41684 -3454
rect 42115 -3460 42160 -3454
rect 42176 -3460 42204 -3454
rect 42115 -3475 42204 -3460
rect 42232 -3475 42260 -3454
rect 42297 -3475 42342 -3454
rect 42773 -3475 42807 -3454
rect 41457 -3494 42590 -3475
rect 41457 -3604 41491 -3494
rect 41494 -3516 42590 -3494
rect 42773 -3488 42820 -3475
rect 42773 -3506 42822 -3488
rect 41500 -3522 42164 -3516
rect 42173 -3522 42590 -3516
rect 42761 -3522 42822 -3506
rect 41500 -3562 41546 -3522
rect 41550 -3556 42164 -3522
rect 41550 -3562 41574 -3556
rect 41494 -3604 41546 -3562
rect 41457 -3606 41546 -3604
rect 41457 -3615 41564 -3606
rect 41457 -4718 41491 -3615
rect 41500 -3846 41564 -3615
rect 41500 -4591 41546 -3846
rect 41574 -3874 41592 -3578
rect 41639 -3636 41684 -3556
rect 42103 -3562 42160 -3556
rect 42180 -3562 42204 -3522
rect 42208 -3556 42822 -3522
rect 42208 -3562 42260 -3556
rect 42103 -3603 42204 -3562
rect 42115 -3636 42204 -3603
rect 41494 -4644 41546 -4591
rect 41639 -4603 41673 -3636
rect 42115 -4603 42149 -3636
rect 42158 -4330 42204 -3636
rect 42232 -4274 42260 -3562
rect 42297 -3636 42342 -3556
rect 42761 -3603 42807 -3556
rect 42838 -3599 42866 -3454
rect 42773 -3604 42807 -3603
rect 42816 -3604 42866 -3599
rect 42773 -3606 42866 -3604
rect 42894 -3550 42922 -3454
rect 42930 -3482 42989 -3454
rect 42930 -3550 42998 -3482
rect 42894 -3606 42998 -3550
rect 42773 -3615 42888 -3606
rect 42232 -4330 42276 -4274
rect 42158 -4591 42220 -4330
rect 42152 -4598 42220 -4591
rect 42232 -4598 42248 -4330
rect 42152 -4603 42204 -4598
rect 41522 -4690 41546 -4644
rect 41550 -4650 41574 -4644
rect 41639 -4650 41686 -4603
rect 42103 -4644 42204 -4603
rect 42232 -4644 42276 -4598
rect 42103 -4650 42164 -4644
rect 41550 -4684 42164 -4650
rect 41550 -4690 41574 -4684
rect 41448 -4730 41491 -4718
rect 41494 -4730 41546 -4690
rect 41448 -4746 41546 -4730
rect 41448 -4752 41502 -4746
rect 41518 -4752 41546 -4746
rect 41639 -4730 41673 -4684
rect 41676 -4730 42088 -4684
rect 42103 -4700 42149 -4684
rect 42180 -4690 42204 -4644
rect 42208 -4650 42276 -4644
rect 42297 -4603 42331 -3636
rect 42773 -4603 42807 -3615
rect 42816 -3954 42888 -3615
rect 42894 -3954 42916 -3606
rect 42930 -3954 42998 -3606
rect 42816 -4603 42866 -3954
rect 42297 -4650 42344 -4603
rect 42761 -4607 42866 -4603
rect 42761 -4616 42820 -4607
rect 42761 -4650 42822 -4616
rect 42208 -4684 42822 -4650
rect 42208 -4690 42260 -4684
rect 41639 -4752 42088 -4730
rect 42115 -4730 42149 -4700
rect 42152 -4730 42204 -4690
rect 42115 -4746 42204 -4730
rect 42115 -4752 42160 -4746
rect 42176 -4752 42204 -4746
rect 42232 -4752 42260 -4690
rect 42297 -4730 42331 -4684
rect 42297 -4752 42342 -4730
rect 42352 -4752 42734 -4684
rect 42761 -4700 42807 -4684
rect 42773 -4730 42807 -4700
rect 42773 -4752 42818 -4730
rect 42838 -4752 42866 -4607
rect 42894 -4010 42998 -3954
rect 42894 -4752 42922 -4010
rect 42930 -4690 42998 -4010
rect 43206 -4670 43210 -4662
rect 42930 -4730 42989 -4690
rect 42930 -4752 43000 -4730
rect 41386 -4786 43000 -4752
rect 41457 -5262 41502 -4786
rect 41457 -8840 41491 -5262
rect 41518 -8893 41546 -4786
rect 41639 -5110 42088 -4786
rect 41639 -5262 41684 -5110
rect 41876 -5118 42088 -5110
rect 42115 -5262 42160 -4786
rect 41639 -8840 41673 -5262
rect 42115 -8840 42149 -5262
rect 42176 -8893 42204 -4786
rect 42232 -8893 42260 -4786
rect 42297 -5262 42342 -4786
rect 42352 -5110 42734 -4786
rect 42352 -5118 42564 -5110
rect 42773 -5262 42818 -4786
rect 42297 -8840 42331 -5262
rect 42773 -8840 42807 -5262
rect 42838 -8893 42866 -4786
rect 42894 -8893 42922 -4786
rect 42955 -5262 43000 -4786
rect 43218 -5110 43222 -4670
rect 43431 -4730 43465 -1544
rect 43508 -3418 43536 -1544
rect 43564 -3418 43592 -1544
rect 43613 -3418 43647 -1544
rect 44089 -3418 44123 -1544
rect 44216 -3418 44244 -1544
rect 44271 -3418 44305 -1544
rect 44385 -3418 44419 -1544
rect 44747 -3418 44781 -3384
rect 44861 -3418 44895 -1544
rect 43472 -3452 44954 -3418
rect 43472 -4730 43506 -3452
rect 43508 -3606 43536 -3452
rect 43564 -3602 43592 -3452
rect 43613 -3520 43647 -3452
rect 44089 -3473 44123 -3452
rect 44216 -3473 44244 -3452
rect 44089 -3504 44136 -3473
rect 44077 -3520 44136 -3504
rect 44216 -3520 44263 -3473
rect 43613 -3554 44263 -3520
rect 44271 -3520 44305 -3452
rect 44385 -3520 44419 -3452
rect 44747 -3504 44793 -3473
rect 44735 -3520 44793 -3504
rect 44271 -3554 44793 -3520
rect 43613 -3602 43647 -3554
rect 44077 -3601 44135 -3554
rect 43564 -3606 43647 -3602
rect 43575 -3613 43647 -3606
rect 43586 -3862 43647 -3613
rect 43431 -4750 43506 -4730
rect 43508 -4750 43536 -3862
rect 43564 -4589 43647 -3862
rect 43564 -4750 43592 -4589
rect 43613 -4648 43647 -4589
rect 44089 -4601 44123 -3601
rect 44077 -4648 44136 -4601
rect 44160 -4642 44188 -3560
rect 44216 -3602 44244 -3560
rect 44271 -3602 44305 -3554
rect 44216 -4589 44305 -3602
rect 44216 -4601 44244 -4589
rect 44216 -4648 44263 -4601
rect 43613 -4682 44263 -4648
rect 44271 -4648 44305 -4589
rect 44385 -4648 44419 -3554
rect 44735 -3601 44793 -3554
rect 44861 -3520 44895 -3452
rect 44861 -3563 44890 -3520
rect 44747 -4601 44781 -3601
rect 44735 -4648 44793 -4601
rect 44271 -4682 44793 -4648
rect 44861 -4639 44895 -3563
rect 44902 -4605 44929 -3597
rect 45576 -3904 45610 -516
rect 46348 -603 46382 -599
rect 46342 -628 46382 -603
rect 47006 -628 47040 -599
rect 47664 -628 47698 -599
rect 48322 -628 48356 -599
rect 48980 -628 49014 -599
rect 45902 -664 49164 -628
rect 56050 -664 57423 -633
rect 45902 -698 49870 -664
rect 56050 -669 60480 -664
rect 51111 -698 60480 -669
rect 45902 -766 49164 -698
rect 51111 -703 57423 -698
rect 49286 -760 49314 -734
rect 49456 -750 49467 -739
rect 49479 -750 49490 -739
rect 49456 -766 49490 -750
rect 45902 -800 49490 -766
rect 45902 -839 49164 -800
rect 49172 -839 49194 -834
rect 45042 -4194 45050 -4140
rect 45540 -4158 45776 -3904
rect 45536 -4194 45776 -4158
rect 45902 -4194 49194 -839
rect 44861 -4658 44890 -4639
rect 43613 -4730 43647 -4682
rect 43613 -4750 43658 -4730
rect 43694 -4750 44076 -4682
rect 44077 -4698 44135 -4682
rect 44089 -4730 44123 -4698
rect 44089 -4750 44134 -4730
rect 44216 -4750 44244 -4688
rect 44271 -4730 44305 -4682
rect 44271 -4750 44316 -4730
rect 44340 -4750 44552 -4682
rect 44735 -4698 44793 -4682
rect 44830 -4682 44890 -4658
rect 44830 -4684 44895 -4682
rect 44778 -4713 44793 -4698
rect 44664 -4738 44678 -4732
rect 44664 -4744 44741 -4738
rect 44747 -4750 44781 -4716
rect 44861 -4738 44895 -4684
rect 44938 -4732 44942 -4688
rect 44787 -4744 44942 -4738
rect 44861 -4750 44895 -4744
rect 43431 -4784 44954 -4750
rect 45096 -4760 45104 -4194
rect 45536 -4228 49194 -4194
rect 45536 -4296 45776 -4228
rect 45786 -4296 45833 -4249
rect 45536 -4330 45833 -4296
rect 45536 -4577 45776 -4330
rect 45803 -4389 45848 -4378
rect 45814 -4565 45848 -4389
rect 45536 -4603 45833 -4577
rect 45536 -4616 45776 -4603
rect 45536 -4634 45790 -4616
rect 45536 -4650 45786 -4634
rect 45902 -4650 49194 -4228
rect 45536 -4684 49194 -4650
rect 43431 -5262 43476 -4784
rect 42955 -8840 42989 -5262
rect 43431 -8840 43465 -5262
rect 43508 -8893 43536 -4784
rect 43564 -8893 43592 -4784
rect 43613 -5262 43658 -4784
rect 43694 -5118 44076 -4784
rect 44089 -5262 44134 -4784
rect 43613 -8840 43647 -5262
rect 44089 -8840 44123 -5262
rect 44216 -8893 44244 -4784
rect 44271 -5262 44316 -4784
rect 44340 -4894 44638 -4784
rect 44340 -5118 44552 -4894
rect 44271 -8840 44305 -5262
rect 44385 -8899 44419 -5118
rect 41343 -8933 44419 -8899
rect 41343 -8949 41377 -8933
rect 41518 -8946 41546 -8939
rect 42176 -8946 42204 -8939
rect 42232 -8946 42260 -8939
rect 42838 -8946 42866 -8939
rect 42894 -8946 42922 -8939
rect 43508 -8946 43536 -8939
rect 43564 -8946 43592 -8939
rect 44216 -8946 44244 -8939
rect 41343 -8960 41354 -8949
rect 41366 -8960 41377 -8949
rect 44385 -8949 44419 -8933
rect 44861 -8939 44895 -4784
rect 45082 -4820 45086 -4810
rect 45136 -4950 45156 -4714
rect 45164 -4978 45184 -4686
rect 45536 -4692 45776 -4684
rect 45232 -4712 45352 -4710
rect 45536 -4712 45828 -4692
rect 45902 -4704 49194 -4684
rect 45838 -4712 49194 -4704
rect 45536 -4720 45776 -4712
rect 45536 -4726 45834 -4720
rect 45204 -4740 45380 -4738
rect 45536 -4752 45866 -4726
rect 45902 -4730 49194 -4712
rect 49206 -4730 49228 -800
rect 45902 -4752 49205 -4730
rect 45536 -4786 49205 -4752
rect 45536 -4796 45776 -4786
rect 45902 -4810 49205 -4786
rect 45558 -4822 49205 -4810
rect 45938 -4942 45972 -4822
rect 46080 -4892 46092 -4822
rect 46108 -4864 46120 -4822
rect 45256 -4990 45332 -4988
rect 45228 -5018 45360 -5016
rect 45238 -5240 45348 -5220
rect 45276 -5278 45310 -5258
rect 45910 -5298 45972 -4942
rect 46082 -4948 46092 -4892
rect 46110 -4920 46120 -4864
rect 45938 -6376 45972 -5298
rect 46414 -6376 46448 -4822
rect 46528 -5262 46573 -4822
rect 46604 -5194 46632 -4994
rect 46710 -5262 46755 -4822
rect 46772 -5138 47174 -4822
rect 46962 -5142 47174 -5138
rect 47186 -5262 47231 -4822
rect 46528 -6376 46562 -5262
rect 46604 -6376 46632 -5394
rect 45102 -6398 46670 -6376
rect 45102 -6402 46632 -6398
rect 45938 -8916 45972 -6402
rect 46414 -8876 46448 -6402
rect 46528 -8826 46562 -6402
rect 46604 -8826 46632 -6402
rect 46710 -8826 46744 -5262
rect 47186 -8826 47220 -5262
rect 47256 -8810 47284 -4822
rect 47312 -8810 47340 -4822
rect 47368 -5262 47413 -4822
rect 47438 -5138 47822 -4822
rect 47438 -5142 47650 -5138
rect 47844 -5262 47889 -4822
rect 47368 -8826 47402 -5262
rect 47844 -8826 47878 -5262
rect 47914 -8870 47942 -4822
rect 47970 -8826 47998 -4822
rect 48026 -5262 48071 -4822
rect 48086 -5138 48490 -4822
rect 48278 -5144 48490 -5138
rect 48502 -5262 48547 -4822
rect 48026 -8826 48060 -5262
rect 48502 -8826 48536 -5262
rect 48578 -8870 48606 -4822
rect 48634 -8870 48662 -4822
rect 48684 -5262 48729 -4822
rect 48754 -5144 49134 -4822
rect 48922 -5156 49134 -5144
rect 49160 -5262 49205 -4822
rect 48684 -8826 48718 -5262
rect 49160 -8826 49194 -5262
rect 49206 -5298 49228 -5262
rect 49286 -8870 49314 -806
rect 49331 -850 49387 -839
rect 49342 -5298 49387 -850
rect 49342 -8826 49376 -5298
rect 49456 -8876 49490 -800
rect 51015 -7380 51049 -765
rect 53835 -771 53869 -733
rect 54533 -755 54544 -744
rect 54556 -755 54567 -744
rect 54533 -771 54567 -755
rect 53835 -805 54567 -771
rect 49856 -7670 49864 -7616
rect 50979 -7634 51066 -7380
rect 49874 -8272 50002 -7634
rect 50012 -8053 50020 -7853
rect 50350 -8168 50590 -7634
rect 50826 -7670 51066 -7634
rect 51129 -7670 51190 -7636
rect 50826 -7704 51252 -7670
rect 50044 -8188 50164 -8168
rect 50350 -8188 50640 -8168
rect 50826 -8186 51066 -7704
rect 51096 -7738 51112 -7734
rect 51068 -7766 51084 -7762
rect 51068 -7812 51088 -7766
rect 51068 -7814 51084 -7812
rect 51096 -7840 51116 -7738
rect 51117 -7806 51123 -7725
rect 51096 -7842 51112 -7840
rect 51129 -7865 51163 -7704
rect 51104 -8041 51163 -7865
rect 51110 -8124 51114 -8098
rect 51117 -8134 51123 -8053
rect 51129 -8168 51163 -8041
rect 50826 -8188 51096 -8186
rect 50350 -8196 50590 -8188
rect 50038 -8216 50192 -8196
rect 50350 -8216 50668 -8196
rect 50690 -8214 50714 -8196
rect 50826 -8202 51066 -8188
rect 51129 -8202 51190 -8168
rect 51218 -8202 51252 -7704
rect 50718 -8214 50742 -8208
rect 50350 -8272 50590 -8216
rect 50826 -8236 51252 -8202
rect 50826 -8272 51066 -8236
rect 49932 -8418 49966 -8272
rect 51015 -8286 51049 -8272
rect 49928 -8774 49966 -8418
rect 50008 -8470 50198 -8468
rect 50036 -8498 50082 -8496
rect 50124 -8498 50170 -8496
rect 46114 -8910 49790 -8876
rect 46414 -8926 46448 -8910
rect 47914 -8922 47942 -8916
rect 46414 -8937 46425 -8926
rect 46437 -8937 46448 -8926
rect 48578 -8928 48606 -8916
rect 48634 -8922 48662 -8916
rect 49286 -8928 49314 -8916
rect 49456 -8926 49490 -8910
rect 49932 -8916 49966 -8774
rect 50979 -8906 51266 -8286
rect 53835 -8899 53869 -805
rect 53938 -864 53983 -853
rect 54408 -864 54453 -853
rect 53949 -8840 53983 -864
rect 54168 -4670 54380 -4662
rect 54012 -5110 54380 -4670
rect 54012 -5118 54224 -5110
rect 54419 -8840 54453 -864
rect 54533 -1158 54567 -805
rect 55945 -839 55972 -737
rect 55973 -811 56000 -765
rect 54533 -2510 54570 -1158
rect 54533 -8899 54567 -2510
rect 55244 -4228 55634 -4194
rect 55244 -4726 55278 -4228
rect 55458 -4296 55505 -4249
rect 55420 -4330 55505 -4296
rect 55347 -4389 55392 -4378
rect 55475 -4389 55520 -4378
rect 55358 -4565 55392 -4389
rect 55486 -4565 55520 -4389
rect 55458 -4624 55505 -4577
rect 55420 -4658 55505 -4624
rect 55478 -4662 55484 -4658
rect 55490 -4698 55496 -4662
rect 55600 -4726 55634 -4228
rect 55244 -4760 55634 -4726
rect 55230 -5430 55652 -4810
rect 55923 -5426 55957 -864
rect 56000 -2504 56002 -1152
rect 56000 -4578 56018 -4004
rect 56050 -4704 57423 -703
rect 58906 -766 58940 -719
rect 59604 -750 59615 -739
rect 59627 -750 59638 -739
rect 59604 -766 59638 -750
rect 58906 -800 59638 -766
rect 58090 -1808 58226 -1698
rect 58090 -1834 58242 -1808
rect 58150 -2266 58242 -1834
rect 58028 -4696 58490 -4158
rect 56050 -4960 57432 -4704
rect 57446 -4932 57488 -4732
rect 58028 -4762 58638 -4696
rect 58028 -4796 58700 -4762
rect 58148 -4846 58174 -4812
rect 58426 -4838 58700 -4796
rect 58426 -4846 58638 -4838
rect 58086 -4880 58638 -4846
rect 55858 -5512 55957 -5426
rect 55808 -6376 55834 -5572
rect 55836 -6376 55862 -5572
rect 55923 -6376 55957 -5512
rect 56000 -5572 56002 -5024
rect 56050 -6376 57423 -4960
rect 58086 -5360 58120 -4880
rect 58174 -4986 58208 -4880
rect 58278 -4948 58316 -4910
rect 58228 -4982 58242 -4948
rect 58244 -4982 58316 -4948
rect 58174 -5018 58214 -4986
rect 58224 -4990 58242 -4986
rect 58278 -4990 58300 -4986
rect 58306 -5018 58328 -4986
rect 58174 -5032 58208 -5018
rect 58220 -5032 58234 -5021
rect 58277 -5032 58322 -5021
rect 58174 -5208 58234 -5032
rect 58288 -5208 58322 -5032
rect 58402 -5144 58638 -4880
rect 58798 -4920 58802 -4720
rect 58826 -4948 58830 -4692
rect 58174 -5222 58208 -5208
rect 58278 -5222 58316 -5220
rect 58174 -5326 58214 -5222
rect 58228 -5308 58242 -5250
rect 58278 -5258 58322 -5222
rect 58244 -5292 58322 -5258
rect 58278 -5308 58294 -5292
rect 58148 -5336 58214 -5326
rect 58306 -5336 58322 -5292
rect 58148 -5360 58208 -5336
rect 58402 -5360 58436 -5144
rect 58086 -5394 58436 -5360
rect 58798 -5572 58822 -5024
rect 58826 -5320 58850 -4996
rect 58826 -5600 58854 -5320
rect 58832 -5606 58854 -5600
rect 58278 -6374 58280 -6174
rect 55250 -6402 57423 -6376
rect 58306 -6402 58308 -6146
rect 55244 -7800 55318 -7470
rect 55244 -7954 55450 -7800
rect 55244 -8124 55318 -7954
rect 55808 -8893 55834 -6402
rect 55836 -8893 55862 -6402
rect 55923 -8840 55957 -6402
rect 49456 -8937 49467 -8926
rect 49479 -8937 49490 -8926
rect 44385 -8960 44396 -8949
rect 44408 -8960 44419 -8949
rect 40963 -9035 44799 -9001
rect 46034 -9012 49870 -8978
rect 52440 -9001 53410 -8900
rect 53835 -8933 54567 -8899
rect 53835 -8949 53869 -8933
rect 53835 -8960 53846 -8949
rect 53858 -8960 53869 -8949
rect 54533 -8949 54567 -8933
rect 55808 -8946 55834 -8939
rect 54533 -8960 54544 -8949
rect 54556 -8960 54567 -8949
rect 55836 -8974 55862 -8939
rect 56050 -8978 57423 -6402
rect 57474 -8536 57488 -7134
rect 58278 -7974 58290 -7774
rect 58306 -8002 58318 -7746
rect 58768 -8600 58794 -7142
rect 58796 -8572 58822 -7170
rect 58902 -8572 58904 -7170
rect 58906 -8876 58940 -800
rect 59009 -850 59054 -839
rect 59479 -850 59524 -839
rect 59020 -8826 59054 -850
rect 59264 -4708 59476 -4690
rect 59070 -5138 59476 -4708
rect 59070 -5156 59282 -5138
rect 59490 -8826 59524 -850
rect 59604 -1414 59638 -800
rect 59604 -2518 59656 -1414
rect 59604 -8876 59638 -2518
rect 59688 -7698 59712 -7540
rect 59726 -7660 59750 -7578
rect 60022 -8272 60484 -7634
rect 60498 -8272 60960 -7634
rect 63031 -7670 63065 -765
rect 63107 -7660 63108 -7578
rect 63145 -7636 63146 -7540
rect 63145 -7670 63206 -7636
rect 62974 -7704 63268 -7670
rect 63031 -7772 63065 -7704
rect 63038 -7815 63065 -7772
rect 63133 -7806 63139 -7725
rect 62997 -8057 63026 -7849
rect 63031 -8091 63065 -7815
rect 63145 -7865 63179 -7704
rect 63120 -8041 63179 -7865
rect 63038 -8134 63065 -8091
rect 63126 -8124 63130 -8098
rect 63133 -8134 63139 -8053
rect 63031 -8168 63065 -8134
rect 63145 -8168 63179 -8041
rect 63012 -8188 63112 -8168
rect 63031 -8196 63065 -8188
rect 63006 -8202 63112 -8196
rect 63145 -8202 63206 -8168
rect 63234 -8202 63268 -7704
rect 62974 -8236 63268 -8202
rect 63354 -7704 63744 -7670
rect 63354 -8202 63388 -7704
rect 63568 -7772 63615 -7725
rect 63530 -7806 63615 -7772
rect 63457 -7865 63502 -7854
rect 63585 -7865 63630 -7854
rect 63468 -8041 63502 -7865
rect 63596 -8041 63630 -7865
rect 63568 -8100 63615 -8053
rect 63530 -8134 63615 -8100
rect 63710 -8202 63744 -7704
rect 63354 -8236 63744 -8202
rect 63892 -8214 63902 -7864
rect 63920 -8214 63930 -7836
rect 63026 -8248 63065 -8236
rect 63031 -8286 63065 -8248
rect 60336 -8322 60364 -8288
rect 60076 -8356 60426 -8322
rect 59712 -8830 59726 -8808
rect 60076 -8836 60110 -8356
rect 60268 -8424 60306 -8386
rect 60234 -8458 60306 -8424
rect 60266 -8466 60288 -8462
rect 60179 -8508 60224 -8497
rect 60244 -8500 60252 -8470
rect 60294 -8494 60316 -8462
rect 60336 -8470 60346 -8458
rect 60272 -8497 60280 -8496
rect 60302 -8497 60312 -8494
rect 60267 -8508 60312 -8497
rect 60190 -8684 60224 -8508
rect 60278 -8684 60312 -8508
rect 60302 -8696 60312 -8684
rect 60268 -8700 60312 -8696
rect 60268 -8734 60306 -8700
rect 60336 -8722 60350 -8470
rect 60336 -8734 60346 -8722
rect 60234 -8768 60306 -8734
rect 60358 -8802 60370 -8356
rect 60336 -8826 60370 -8802
rect 60358 -8830 60370 -8826
rect 60392 -8836 60426 -8356
rect 59674 -8870 59690 -8842
rect 58906 -8910 59638 -8876
rect 59646 -8876 59662 -8870
rect 59646 -8898 59666 -8876
rect 59658 -8910 59666 -8898
rect 58906 -8926 58940 -8910
rect 58906 -8937 58917 -8926
rect 58929 -8937 58940 -8926
rect 59604 -8926 59638 -8910
rect 59604 -8937 59615 -8926
rect 59627 -8937 59638 -8926
rect 59692 -8944 59700 -8842
rect 60076 -8870 60426 -8836
rect 60552 -8356 60902 -8322
rect 60552 -8836 60586 -8356
rect 60744 -8424 60782 -8386
rect 60710 -8458 60782 -8424
rect 60655 -8508 60700 -8497
rect 60743 -8508 60788 -8497
rect 60666 -8684 60700 -8508
rect 60754 -8684 60788 -8508
rect 60744 -8734 60782 -8696
rect 60710 -8768 60782 -8734
rect 60868 -8836 60902 -8356
rect 60552 -8870 60902 -8836
rect 59740 -8902 60308 -8876
rect 59740 -8910 60310 -8902
rect 60358 -8944 60374 -8870
rect 60386 -8916 60402 -8870
rect 62995 -8906 63282 -8286
rect 63336 -8906 63758 -8286
rect 63892 -8688 63902 -8400
rect 63920 -8716 63930 -8400
rect 63167 -8967 63194 -8906
rect 63195 -8939 63222 -8906
rect 56050 -9001 60480 -8978
rect 51111 -9012 60480 -9001
rect 51111 -9035 57423 -9012
rect 52440 -9071 53410 -9035
rect 56050 -9048 57423 -9035
rect 52884 -9332 52956 -9324
rect 62080 -9332 62152 -9324
rect 52884 -9334 52952 -9332
rect 62080 -9334 62148 -9332
rect 47080 -9822 47084 -9502
rect 47118 -9822 47122 -9502
rect 62162 -9552 62182 -9373
rect 62162 -9573 62192 -9552
rect 62128 -9912 62186 -9910
rect 62102 -9946 62152 -9944
<< pdiodelvtc >>
rect 36628 -2808 36736 -2682
<< locali >>
rect 15024 33870 16026 33956
rect 15024 32316 15094 33870
rect 15952 32316 16026 33870
rect 15024 12840 16026 32316
rect 35070 14078 36124 14218
rect 35070 13732 35278 14078
rect 35988 13732 36124 14078
rect 35070 13152 36124 13732
rect 35070 9588 36820 13152
rect 35070 4060 36124 9588
rect 47350 5426 50654 5440
rect 47350 4492 50706 5426
rect 19378 -6684 20292 3040
rect 35048 2518 36128 4060
rect 35048 1920 37074 2518
rect 35048 -6596 36128 1920
rect 40140 -3316 42584 -2318
rect 40140 -3376 42588 -3316
rect 40140 -3494 42590 -3376
rect 41500 -3636 42590 -3494
rect 49206 -5298 50706 4492
rect 18628 -6810 21072 -6684
rect 18628 -7506 18770 -6810
rect 20886 -7506 21072 -6810
rect 18628 -7688 21072 -7506
rect 33864 -6774 37084 -6596
rect 33864 -7668 34260 -6774
rect 36852 -7668 37084 -6774
rect 33864 -7816 37084 -7668
<< viali >>
rect 15094 32316 15952 33870
rect 35278 13732 35988 14078
rect 18770 -7506 20886 -6810
rect 34260 -7668 36852 -6774
<< metal1 >>
rect 15054 33870 16000 33918
rect 15054 32316 15094 33870
rect 15952 32316 16000 33870
rect 15054 32232 16000 32316
rect 22946 32740 24126 32954
rect 22946 32406 23126 32740
rect 23972 32406 24126 32740
rect 22946 31358 24126 32406
rect 46946 32772 48150 32880
rect 46946 32248 47056 32772
rect 48054 32248 48150 32772
rect 22934 22368 24150 23238
rect 22916 13726 24116 14248
rect 34120 14078 36970 31590
rect 46946 31404 48150 32248
rect 46934 21856 48162 23084
rect 34120 13732 35278 14078
rect 35988 13732 36970 14078
rect 22916 13712 33790 13726
rect 22916 13504 33816 13712
rect 34120 13528 36970 13732
rect 33204 13126 33816 13504
rect 33178 12720 34640 13126
rect 47028 12590 48112 14026
rect 23816 4806 24178 5548
rect 22950 2730 24178 4806
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
rect 0 -2400 200 -2200
rect 0 -2800 200 -2600
rect 0 -3200 200 -3000
rect 0 -3600 200 -3400
rect 18628 -6810 21072 -6684
rect 18628 -7506 18770 -6810
rect 20886 -7506 21072 -6810
rect 18628 -7688 21072 -7506
rect 33864 -6774 37084 -6596
rect 33864 -7668 34260 -6774
rect 36852 -7668 37084 -6774
rect 33864 -7816 37084 -7668
<< via1 >>
rect 15094 32316 15952 33870
rect 23126 32406 23972 32740
rect 47056 32248 48054 32772
rect 22222 6310 22362 6456
rect 23548 -2018 23910 -962
rect 18770 -7506 20886 -6810
rect 34260 -7668 36852 -6774
<< metal2 >>
rect 14628 33870 57258 36292
rect 14628 32316 15094 33870
rect 15952 32772 57258 33870
rect 15952 32740 47056 32772
rect 15952 32406 23126 32740
rect 23972 32406 47056 32740
rect 15952 32316 47056 32406
rect 14628 32248 47056 32316
rect 48054 32248 57258 32772
rect 14628 32156 57258 32248
rect 16718 9180 17114 9292
rect 16718 8572 16762 9180
rect 17070 8572 17114 9180
rect 16718 8460 17114 8572
rect 22200 6456 22376 6472
rect 22200 6310 22222 6456
rect 22362 6310 22376 6456
rect 22200 6290 22376 6310
rect 31452 3880 39416 31570
rect 43930 18196 56166 18372
rect 43930 17776 55314 18196
rect 56030 17776 56166 18196
rect 43930 17516 56166 17776
rect 16844 2090 17410 2230
rect 16844 1868 16970 2090
rect 17302 1868 17410 2090
rect 16844 1720 17410 1868
rect 23430 -962 26630 2892
rect 23430 -2018 23548 -962
rect 23910 -2018 26630 -962
rect 23430 -4916 26630 -2018
rect 36202 -2642 36780 3880
rect 22856 -6432 26660 -4916
rect 14582 -6774 57212 -6432
rect 14582 -6810 34260 -6774
rect 14582 -7506 18770 -6810
rect 20886 -7506 34260 -6810
rect 14582 -7668 34260 -7506
rect 36852 -7668 57212 -6774
rect 14582 -10568 57212 -7668
<< via2 >>
rect 30942 27254 31096 27416
rect 26260 23556 27224 24248
rect 30930 18268 31106 18436
rect 26148 14606 27300 15542
rect 16762 8572 17070 9180
rect 25368 8598 25938 9180
rect 27202 8670 27364 8830
rect 21122 6370 21222 6454
rect 22236 6330 22348 6438
rect 39996 27186 40162 27404
rect 44146 27008 44952 27430
rect 39952 17902 40124 18066
rect 55314 17776 56030 18196
rect 40068 8796 40228 8974
rect 44222 8624 45018 9066
rect 16970 1868 17302 2090
rect 27102 -1626 27260 -1470
rect 31500 -1652 31890 -1280
rect 41928 -2498 42036 -2434
rect 37518 -4376 37628 -4258
<< metal3 >>
rect 20550 29986 22164 30292
rect 20550 28896 40436 29986
rect 20550 28632 22164 28896
rect 20572 27644 22186 28072
rect 20572 27416 31334 27644
rect 20572 27254 30942 27416
rect 31096 27254 31334 27416
rect 20572 26824 31334 27254
rect 39788 27404 40430 28896
rect 39788 27186 39996 27404
rect 40162 27186 40430 27404
rect 39788 27068 40430 27186
rect 44044 27430 45012 27488
rect 44044 27008 44146 27430
rect 44952 27008 45012 27430
rect 44044 26942 45012 27008
rect 20572 26412 22186 26824
rect 26150 24248 27368 24346
rect 26150 23556 26260 24248
rect 27224 23556 27368 24248
rect 26150 23446 27368 23556
rect 20594 20878 22208 21304
rect 20594 20000 40506 20878
rect 20594 19644 22208 20000
rect 20616 18664 22230 19130
rect 20616 18436 31258 18664
rect 20616 18268 30930 18436
rect 31106 18268 31258 18436
rect 20616 17856 31258 18268
rect 39654 18066 40490 20000
rect 39654 17902 39952 18066
rect 40124 17902 40490 18066
rect 20616 17470 22230 17856
rect 39654 17780 40490 17902
rect 55248 18196 56070 18248
rect 55248 17776 55314 18196
rect 56030 17776 56070 18196
rect 55248 17704 56070 17776
rect 20616 15340 22230 17000
rect 26094 15542 27478 15704
rect 20932 12410 21958 15340
rect 26094 14606 26148 15542
rect 27300 14606 27478 15542
rect 26094 14498 27478 14606
rect 20932 11616 40604 12410
rect 16744 9180 17092 9258
rect 16744 8572 16762 9180
rect 17070 8572 17092 9180
rect 16744 8506 17092 8572
rect 25252 9180 25996 9236
rect 25252 8598 25368 9180
rect 25938 8598 25996 9180
rect 39810 8974 40588 11616
rect 25252 8518 25996 8598
rect 27126 8830 27436 8888
rect 27126 8670 27202 8830
rect 27364 8670 27436 8830
rect 20890 6454 21304 6548
rect 27126 6498 27436 8670
rect 39810 8796 40068 8974
rect 40228 8796 40588 8974
rect 39810 8628 40588 8796
rect 44166 9066 45096 9160
rect 44166 8624 44222 9066
rect 45018 8624 45096 9066
rect 44166 8552 45096 8624
rect 20890 6370 21122 6454
rect 21222 6370 21304 6454
rect 16844 2090 17410 2230
rect 16844 1868 16970 2090
rect 17302 1868 17410 2090
rect 16844 1720 17410 1868
rect 20890 -902 21304 6370
rect 22180 6438 27460 6498
rect 22180 6330 22236 6438
rect 22348 6330 27460 6438
rect 22180 6258 27460 6330
rect 20636 -1196 21666 -902
rect 31352 -1108 32016 -1102
rect 20636 -1238 22676 -1196
rect 20636 -1848 22884 -1238
rect 24072 -1470 27316 -1238
rect 24072 -1626 27102 -1470
rect 27260 -1626 27316 -1470
rect 24072 -1848 27316 -1626
rect 31352 -1280 32018 -1108
rect 31352 -1652 31500 -1280
rect 31890 -1652 32018 -1280
rect 20636 -1924 22676 -1848
rect 31352 -1894 32018 -1652
rect 31368 -1896 32018 -1894
rect 20636 -2074 21666 -1924
rect 41868 -2234 42188 -2158
rect 41868 -2552 41898 -2234
rect 42136 -2552 42188 -2234
rect 41868 -2564 42188 -2552
rect 35964 -4114 37728 -4064
rect 35954 -4258 37728 -4114
rect 35954 -4376 37518 -4258
rect 37628 -4376 37728 -4258
rect 35954 -4586 37728 -4376
rect 35658 -4606 37728 -4586
rect 35658 -5760 36862 -4606
<< via3 >>
rect 44146 27008 44952 27430
rect 26260 23556 27224 24248
rect 55362 17824 55974 18154
rect 26148 14606 27300 15542
rect 16792 8698 17056 9048
rect 25490 8630 25844 9028
rect 44222 8624 45018 9066
rect 41898 -2434 42136 -2234
rect 41898 -2498 41928 -2434
rect 41928 -2498 42036 -2434
rect 42036 -2498 42136 -2434
rect 41898 -2552 42136 -2498
<< metal4 >>
rect 43928 27430 50272 27584
rect 43928 27008 44146 27430
rect 44952 27008 50272 27430
rect 43928 26774 50272 27008
rect 26058 24248 50282 24536
rect 26058 23556 26260 24248
rect 27224 23556 50282 24248
rect 26058 23260 50282 23556
rect 54812 18154 57228 31570
rect 54772 17824 55362 18154
rect 55974 17824 57228 18154
rect 16328 15236 18180 17016
rect 25976 15542 50196 15820
rect 16720 9332 17814 15236
rect 25976 14606 26148 15542
rect 27300 14606 50196 15542
rect 25976 14396 50196 14606
rect 16682 9048 26064 9332
rect 16682 8698 16792 9048
rect 17056 9028 26064 9048
rect 17056 8698 25490 9028
rect 16682 8630 25490 8698
rect 25844 8630 26064 9028
rect 16682 8386 26064 8630
rect 44038 9066 50258 9232
rect 44038 8624 44222 9066
rect 45018 8624 50258 9066
rect 44038 8436 50258 8624
rect 54812 6018 57228 17824
rect 54834 1498 57198 6018
rect 53568 1454 57198 1498
rect 46982 1092 57198 1454
rect 46982 1082 54970 1092
rect 53568 1048 54970 1082
rect 31368 -1646 42344 -1066
rect 31368 -1868 42348 -1646
rect 41794 -2234 42348 -1868
rect 41794 -2552 41898 -2234
rect 42136 -2552 42348 -2234
rect 41794 -2600 42348 -2552
use curr_mir  curr_mir_0
timestamp 1695461801
transform 1 0 72116 0 1 7240
box 0 -400 11334 10390
use curr_mir  curr_mir_1
timestamp 1695461801
transform 1 0 10148 0 1 -10168
box 0 -400 11334 10390
use curr_mir  curr_mir_2
timestamp 1695461801
transform 1 0 0 0 1 -10168
box 0 -400 11334 10390
use not  not_0
timestamp 1695461801
transform 1 0 20522 0 1 6220
box 0 -578 1868 990
use not  not_1
timestamp 1695461801
transform 1 0 61066 0 1 -9990
box 0 -578 1868 990
use not  not_2
timestamp 1695461801
transform 1 0 51870 0 1 -9990
box 0 -578 1868 990
use opamp  opamp_0
timestamp 1695461801
transform 1 0 77382 0 1 11126
box 0 -1200 19288 9014
use opamp  opamp_1
timestamp 1695461801
transform 1 0 21482 0 1 -9368
box 0 -1200 19288 9014
use opamp  opamp_2
timestamp 1695461801
transform 1 0 11334 0 1 -9368
box 0 -1200 19288 9014
use switch  switch_0
timestamp 1695461801
transform 1 0 55118 0 1 13320
box -114 -950 10510 11418
use switch  switch_1
timestamp 1695461801
transform 1 0 63874 0 1 13320
box -114 -950 10510 11418
use switch  switch_2
timestamp 1695461801
transform 1 0 96784 0 1 13320
box -114 -950 10510 11418
use switch  switch_3
timestamp 1695461801
transform 1 0 105540 0 1 13320
box -114 -950 10510 11418
use switch  switch_4
timestamp 1695461801
transform 1 0 115688 0 1 13320
box -114 -950 10510 11418
use switch  switch_5
timestamp 1695461801
transform 1 0 55132 0 1 19992
box -114 -950 10510 11418
use switch  switch_6
timestamp 1695461801
transform 1 0 55164 0 1 26356
box -114 -950 10510 11418
use switch  switch_7
timestamp 1695461801
transform 1 0 114 0 1 -9618
box -114 -950 10510 11418
use switch  switch_8
timestamp 1695461801
transform 1 0 40884 0 1 -9618
box -114 -950 10510 11418
use switch  switch_9
timestamp 1695461801
transform 1 0 51032 0 1 -9618
box -114 -950 10510 11418
use switch  switch_10
timestamp 1695461801
transform 1 0 63048 0 1 -9618
box -114 -950 10510 11418
use switch  switch_11
timestamp 1695461801
transform 1 0 30736 0 1 -9618
box -114 -950 10510 11418
use switch  switch_12
timestamp 1695461801
transform 1 0 41360 0 1 -9618
box -114 -950 10510 11418
use switch  switch_13
timestamp 1695461801
transform 1 0 53852 0 1 -9618
box -114 -950 10510 11418
use switch  x1
timestamp 1695461801
transform 0 1 36806 1 0 4546
box -114 -950 10510 11418
use switch  x2
timestamp 1695461801
transform 0 1 23934 -1 0 13086
box -114 -950 10510 11418
use curr_mir  x3
timestamp 1695461801
transform 0 -1 25426 1 0 1738
box 0 -400 11334 10390
use opamp  x4
timestamp 1695461801
transform 1 0 30358 0 -1 3752
box 0 -1200 19288 9014
use switch  x5
timestamp 1695461801
transform 0 1 36696 1 0 13644
box -114 -950 10510 11418
use switch  x6
timestamp 1695461801
transform 0 1 23834 -1 0 2788
box -114 -950 10510 11418
use not  x7
timestamp 1695461801
transform 1 0 113706 0 1 12948
box 0 -578 1868 990
use switch  x8
timestamp 1695461801
transform 0 1 36738 1 0 22948
box -114 -950 10510 11418
use switch  x9
timestamp 1695461801
transform 0 -1 34358 1 0 14018
box -114 -950 10510 11418
use switch  x10
timestamp 1695461801
transform 0 -1 34358 1 0 22992
box -114 -950 10510 11418
use sky130_fd_pr__cap_mim_m3_1_3HBNLG  XC1
timestamp 1695395215
transform 1 0 51818 0 1 9140
box -3186 -3040 3186 3040
use sky130_fd_pr__cap_mim_m3_1_3HBNLG  XC2
timestamp 1695395215
transform 1 0 51818 0 1 15410
box -3186 -3040 3186 3040
use sky130_fd_pr__cap_mim_m3_1_3HBNLG  XC3
timestamp 1695395215
transform 1 0 51832 0 1 22082
box -3186 -3040 3186 3040
use sky130_fd_pr__cap_mim_m3_1_3HBNLG  XC4
timestamp 1695395215
transform 1 0 51864 0 1 28446
box -3186 -3040 3186 3040
<< labels >>
rlabel metal4 54834 1092 57198 17824 1 intout
port 7 nsew
rlabel metal3 20550 28632 22164 30292 1 sw4
port 8 nsew
rlabel metal3 20572 26412 22186 28072 1 sw3
port 9 nsew
rlabel metal3 20594 19644 22208 21304 1 rst
port 10 nsew
rlabel metal3 20616 17470 22230 19130 1 sw2
port 11 nsew
rlabel metal3 20616 15340 22230 17000 1 sw1
port 12 nsew
rlabel metal3 35658 -5760 36862 -4586 1 opbias
port 13 nsew
rlabel metal3 20636 -2074 21666 -902 1 en
port 14 nsew
rlabel metal3 16844 1720 17410 2230 1 Vtune
port 15 nsew
rlabel metal4 16328 15236 18180 17016 1 intin
port 16 nsew
rlabel metal2 14628 32156 57258 36292 1 VDD
port 17 nsew
rlabel metal2 14582 -10568 57212 -6432 1 GROUND
port 18 nsew
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 sw2
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 sw1
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 intin
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 intout
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 opbias
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 en
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 256 0 0 0 Vtune
port 6 nsew
flabel metal1 0 -2800 200 -2600 0 FreeSans 256 0 0 0 rst
flabel metal1 0 -3200 200 -3000 0 FreeSans 256 0 0 0 sw4
flabel metal1 0 -3600 200 -3400 0 FreeSans 256 0 0 0 sw3
<< end >>
