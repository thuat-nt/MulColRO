magic
tech sky130A
magscale 1 2
timestamp 1695698273
<< error_s >>
rect 55147 28845 55181 35209
rect 55261 28941 55295 28975
rect 55919 28941 55953 28975
rect 56577 28941 56611 28975
rect 57235 28941 57269 28975
rect 57893 28941 57927 35110
rect 58551 28941 58605 28975
rect 55211 28907 55215 28941
rect 55227 28907 58605 28941
rect 55115 27035 55181 28845
rect 55257 28855 55261 28873
rect 55257 28839 55307 28855
rect 55318 28845 55336 28860
rect 55346 28845 55364 28858
rect 55859 28839 55906 28886
rect 55915 28855 55919 28873
rect 55915 28839 55965 28855
rect 56517 28845 56564 28886
rect 56508 28839 56564 28845
rect 56573 28855 56577 28873
rect 56573 28839 56623 28855
rect 56638 28845 56644 28848
rect 56666 28845 56672 28858
rect 57175 28839 57222 28886
rect 57231 28855 57235 28873
rect 57231 28839 57281 28855
rect 57833 28845 57880 28886
rect 57893 28873 57927 28907
rect 57828 28839 57880 28845
rect 57889 28855 57927 28873
rect 57889 28839 57939 28855
rect 58491 28839 58538 28886
rect 55261 28805 55906 28839
rect 55919 28805 56564 28839
rect 56577 28805 57222 28839
rect 57235 28805 57880 28839
rect 57893 28805 58538 28839
rect 55261 28758 55307 28805
rect 55217 28746 55235 28758
rect 55261 28746 55295 28758
rect 55217 27134 55295 28746
rect 55318 27458 55336 28799
rect 55346 27430 55364 28799
rect 55919 28758 55965 28805
rect 56508 28799 56529 28805
rect 56536 28771 56557 28805
rect 56577 28758 56623 28805
rect 55876 28746 55907 28757
rect 55919 28746 55953 28758
rect 56534 28746 56565 28757
rect 56577 28746 56611 28758
rect 37878 23697 38134 23706
rect 37906 23669 38106 23678
rect 32410 23400 32976 23434
rect 32410 23112 32444 23400
rect 32781 23320 32792 23331
rect 32465 23258 32546 23305
rect 32605 23286 32792 23320
rect 32793 23258 32874 23305
rect 32512 23220 32546 23258
rect 32565 23220 32821 23226
rect 32840 23220 32874 23258
rect 32565 23206 32822 23220
rect 32781 23198 32792 23203
rect 32593 23192 32793 23198
rect 32593 23178 32794 23192
rect 32832 23178 32928 23192
rect 32605 23158 32792 23178
rect 32942 23164 32976 23400
rect 32804 23150 32976 23164
rect 32567 23120 32819 23123
rect 32942 23112 32976 23150
rect 32410 23089 32976 23112
rect 32410 23078 32444 23089
rect 32942 23078 32976 23089
rect 32410 23077 32976 23078
rect 32444 23063 32942 23077
rect 32410 23044 32976 23063
rect 33026 23026 33646 23448
rect 37500 23074 37516 23076
rect 37408 22965 38028 23074
rect 38140 23060 38582 23094
rect 38078 23033 38644 23060
rect 37408 22931 40320 22965
rect 37408 22895 38028 22931
rect 38078 22766 38112 22931
rect 38180 22897 38214 22900
rect 38508 22897 38542 22900
rect 38610 22766 38644 22931
rect 55115 22173 55149 27035
rect 55217 26973 55263 27134
rect 55816 27081 55826 28480
rect 55844 27109 55854 28452
rect 55887 27134 55953 28746
rect 56545 27134 56611 28746
rect 56638 27446 56644 28799
rect 56666 27418 56672 28799
rect 57235 28758 57281 28805
rect 57828 28799 57845 28805
rect 57856 28771 57873 28805
rect 57893 28758 57939 28805
rect 57192 28746 57223 28757
rect 57235 28746 57269 28758
rect 57850 28746 57881 28757
rect 57893 28746 57927 28758
rect 55887 27122 55921 27134
rect 56545 27122 56579 27134
rect 55875 27109 55934 27122
rect 55844 27100 55934 27109
rect 55941 27100 55972 27109
rect 55875 27081 55934 27100
rect 55816 27075 55934 27081
rect 55323 27041 55934 27075
rect 55969 27075 56000 27081
rect 56533 27075 56592 27122
rect 57126 27081 57146 28486
rect 57154 27109 57174 28458
rect 57203 27134 57269 28746
rect 57861 27134 57927 28746
rect 57960 27424 57964 28799
rect 57988 27396 57992 28799
rect 58508 28746 58539 28757
rect 58551 28746 58585 28907
rect 57203 27122 57237 27134
rect 57861 27122 57895 27134
rect 57191 27109 57250 27122
rect 57154 27106 57250 27109
rect 57257 27106 57282 27109
rect 57191 27081 57250 27106
rect 57126 27078 57250 27081
rect 57285 27078 57310 27081
rect 57191 27075 57250 27078
rect 57849 27075 57908 27122
rect 58448 27081 58468 28456
rect 58476 27081 58496 28428
rect 58519 27134 58585 28746
rect 58633 28845 58651 28907
rect 58665 28845 58699 35209
rect 60218 28850 60252 35214
rect 60332 28946 60366 28980
rect 60990 28946 61024 28980
rect 61648 28946 61682 28980
rect 62306 28946 62340 28980
rect 62964 28946 62998 28980
rect 63622 28946 63676 28980
rect 60282 28912 60286 28946
rect 60298 28912 63676 28946
rect 58519 27122 58553 27134
rect 58507 27075 58565 27122
rect 55969 27072 56592 27075
rect 55981 27041 56592 27072
rect 56639 27041 57250 27075
rect 57297 27041 57908 27075
rect 57955 27041 58565 27075
rect 55875 27025 55921 27041
rect 56533 27025 56579 27041
rect 57191 27025 57237 27041
rect 57849 27025 57895 27041
rect 58507 27025 58553 27041
rect 58633 27035 58699 28845
rect 60186 27058 60252 28850
rect 60328 28860 60332 28878
rect 60328 28844 60378 28860
rect 60930 28844 60968 28882
rect 60986 28860 60990 28878
rect 60986 28844 61036 28860
rect 61588 28850 61626 28882
rect 61578 28844 61626 28850
rect 61644 28860 61648 28878
rect 61644 28844 61694 28860
rect 62246 28844 62284 28882
rect 62302 28860 62306 28878
rect 62302 28844 62352 28860
rect 62904 28844 62942 28882
rect 62960 28860 62964 28878
rect 62960 28844 63010 28860
rect 63562 28844 63600 28882
rect 60332 28810 60968 28844
rect 60990 28840 61626 28844
rect 60990 28810 61628 28840
rect 60332 28772 60378 28810
rect 60990 28772 61036 28810
rect 61578 28804 61600 28810
rect 61606 28776 61628 28810
rect 61648 28810 62284 28844
rect 62306 28810 62942 28844
rect 62964 28810 63600 28844
rect 61648 28772 61694 28810
rect 62306 28772 62352 28810
rect 62900 28804 62916 28810
rect 62928 28776 62944 28804
rect 62964 28772 63010 28810
rect 60288 28760 60306 28772
rect 60332 28760 60366 28772
rect 60947 28760 60978 28771
rect 60990 28760 61024 28772
rect 61605 28760 61636 28771
rect 61648 28760 61682 28772
rect 62263 28760 62294 28771
rect 62306 28760 62340 28772
rect 62921 28760 62952 28771
rect 62964 28760 62998 28772
rect 60288 27148 60366 28760
rect 57861 26973 57895 27025
rect 55217 26939 58565 26973
rect 55229 22269 55263 22303
rect 55887 22269 55921 22303
rect 56545 22269 56579 22303
rect 57203 22269 57237 22303
rect 57861 22269 57895 26939
rect 58519 22269 58553 22303
rect 55197 22235 58587 22269
rect 55101 20671 55149 22173
rect 55229 22183 55263 22235
rect 55887 22214 55921 22235
rect 56545 22214 56579 22235
rect 57203 22214 57237 22235
rect 57861 22214 57895 22235
rect 58519 22214 58553 22235
rect 55845 22183 55921 22214
rect 56503 22183 56579 22214
rect 57161 22183 57237 22214
rect 57819 22183 57895 22214
rect 55229 22086 55275 22183
rect 55845 22167 55933 22183
rect 56503 22167 56591 22183
rect 57161 22167 57249 22183
rect 57819 22167 57907 22183
rect 58477 22167 58553 22214
rect 58633 22173 58667 27035
rect 59880 24746 59882 24794
rect 59852 24718 59882 24738
rect 60186 22178 60220 27058
rect 60288 26996 60334 27148
rect 60886 27104 60912 28224
rect 60914 27104 60940 28196
rect 60958 27148 61024 28760
rect 61616 27148 61682 28760
rect 60958 27136 60992 27148
rect 61616 27136 61650 27148
rect 60946 27098 60996 27136
rect 61050 27104 61068 27120
rect 61604 27098 61654 27136
rect 62206 27104 62222 28206
rect 62234 27104 62250 28178
rect 62274 27148 62340 28760
rect 62932 27148 62998 28760
rect 63030 27402 63036 28804
rect 63058 27374 63064 28804
rect 63579 28760 63610 28771
rect 63622 28760 63656 28912
rect 62274 27136 62308 27148
rect 62932 27136 62966 27148
rect 62262 27098 62312 27136
rect 62920 27098 62970 27136
rect 63514 27104 63538 28208
rect 63542 27104 63566 28180
rect 63590 27148 63656 28760
rect 63704 28850 63722 28912
rect 63736 28850 63770 32670
rect 63590 27136 63624 27148
rect 63578 27098 63628 27136
rect 60394 27064 60996 27098
rect 61052 27064 61654 27098
rect 61710 27064 62312 27098
rect 62368 27064 62970 27098
rect 63026 27064 63628 27098
rect 60946 27048 60992 27064
rect 61604 27048 61650 27064
rect 62262 27048 62308 27064
rect 62920 27048 62966 27064
rect 63578 27048 63624 27064
rect 63704 27058 63770 28850
rect 60958 26996 60992 27048
rect 60288 26962 63636 26996
rect 60300 22274 60334 22308
rect 60958 22274 60992 26962
rect 61616 22274 61650 22308
rect 62274 22274 62308 22308
rect 62932 22274 62966 22308
rect 63590 22274 63624 22308
rect 60268 22240 63658 22274
rect 55277 22133 55933 22167
rect 55935 22133 56591 22167
rect 56593 22133 57249 22167
rect 57251 22133 57907 22167
rect 57909 22133 58553 22167
rect 55853 22127 55857 22133
rect 55881 22099 55885 22133
rect 55887 22086 55933 22133
rect 56545 22086 56591 22133
rect 57169 22127 57173 22133
rect 57197 22099 57201 22133
rect 57203 22086 57249 22133
rect 57861 22086 57907 22133
rect 58485 22127 58489 22133
rect 58513 22099 58517 22133
rect 55229 22074 55263 22086
rect 55862 22074 55875 22085
rect 55887 22074 55921 22086
rect 56520 22074 56533 22085
rect 56545 22074 56579 22086
rect 57178 22074 57191 22085
rect 57203 22074 57237 22086
rect 57836 22074 57849 22085
rect 57861 22074 57895 22086
rect 58494 22074 58507 22085
rect 58519 22074 58553 22133
rect 55215 20770 55263 22074
rect 55873 20770 55921 22074
rect 56531 20770 56579 22074
rect 55101 20160 55135 20671
rect 55215 20609 55249 20770
rect 55873 20758 55907 20770
rect 56531 20758 56565 20770
rect 55251 20643 55255 20745
rect 55279 20711 55283 20717
rect 55859 20711 55907 20758
rect 56517 20711 56565 20758
rect 55275 20677 55283 20711
rect 55291 20677 55907 20711
rect 55933 20677 55941 20711
rect 55949 20677 56565 20711
rect 55279 20671 55283 20677
rect 55861 20661 55907 20677
rect 56519 20661 56565 20677
rect 55873 20609 55907 20661
rect 56531 20609 56565 20661
rect 56567 20643 56571 20745
rect 57112 20717 57114 21814
rect 57140 20717 57142 21786
rect 57189 20770 57237 22074
rect 57847 20770 57895 22074
rect 57189 20758 57223 20770
rect 57847 20758 57881 20770
rect 56595 20711 56599 20717
rect 57175 20711 57223 20758
rect 57833 20711 57881 20758
rect 56591 20677 56599 20711
rect 56607 20677 57223 20711
rect 57249 20677 57257 20711
rect 57265 20677 57881 20711
rect 56595 20671 56599 20677
rect 57112 20664 57114 20671
rect 57140 20636 57142 20671
rect 57177 20661 57223 20677
rect 57835 20661 57881 20677
rect 57189 20609 57223 20661
rect 57847 20609 57881 20661
rect 57883 20643 57887 20745
rect 58434 20717 58436 21784
rect 58462 20717 58464 21756
rect 58505 20770 58553 22074
rect 58505 20758 58539 20770
rect 57911 20711 57915 20717
rect 58491 20711 58539 20758
rect 57907 20677 57915 20711
rect 57923 20677 58539 20711
rect 57911 20671 57915 20677
rect 58434 20664 58436 20671
rect 58462 20636 58464 20671
rect 58493 20661 58539 20677
rect 58505 20609 58539 20661
rect 58619 20671 58667 22173
rect 60172 20694 60220 22178
rect 60300 22188 60334 22240
rect 60916 22206 60954 22210
rect 60300 22100 60346 22188
rect 60916 22172 60956 22206
rect 60348 22138 60956 22172
rect 60924 22132 60928 22138
rect 60952 22104 60956 22138
rect 60958 22188 60992 22240
rect 60958 22100 61004 22188
rect 61574 22172 61612 22210
rect 61006 22138 61612 22172
rect 61616 22188 61650 22240
rect 62232 22206 62270 22210
rect 61616 22100 61662 22188
rect 62232 22172 62272 22206
rect 61664 22138 62272 22172
rect 62240 22132 62244 22138
rect 62268 22104 62272 22138
rect 62274 22188 62308 22240
rect 62274 22100 62320 22188
rect 62890 22172 62928 22210
rect 62322 22138 62928 22172
rect 62932 22188 62966 22240
rect 63548 22206 63586 22210
rect 62932 22100 62978 22188
rect 63548 22172 63588 22206
rect 62980 22138 63588 22172
rect 63556 22132 63560 22138
rect 63584 22104 63588 22138
rect 60300 22088 60334 22100
rect 60933 22088 60946 22099
rect 60958 22088 60992 22100
rect 61591 22088 61604 22099
rect 61616 22088 61650 22100
rect 62249 22088 62262 22099
rect 62274 22088 62308 22100
rect 62907 22088 62920 22099
rect 62932 22088 62966 22100
rect 63565 22088 63578 22099
rect 63590 22088 63624 22240
rect 63704 22178 63738 27058
rect 60286 20784 60334 22088
rect 55203 20575 58551 20609
rect 58619 20160 58653 20671
rect 60172 20160 60206 20694
rect 60286 20632 60320 20784
rect 60322 20666 60326 20768
rect 60872 20740 60880 21552
rect 60900 20740 60908 21524
rect 60944 20784 60992 22088
rect 61602 20784 61650 22088
rect 62260 20784 62308 22088
rect 62918 20784 62966 22088
rect 60944 20772 60978 20784
rect 61602 20772 61636 20784
rect 62260 20772 62294 20784
rect 62918 20772 62952 20784
rect 60350 20734 60354 20740
rect 60930 20734 60978 20772
rect 61588 20734 61636 20772
rect 60346 20700 60354 20734
rect 60362 20700 60978 20734
rect 61004 20700 61012 20734
rect 61020 20700 61636 20734
rect 60350 20694 60354 20700
rect 60872 20688 60880 20694
rect 60900 20660 60908 20694
rect 60932 20684 60978 20700
rect 61590 20684 61636 20700
rect 60944 20632 60978 20684
rect 61602 20632 61636 20684
rect 61638 20666 61642 20768
rect 61666 20734 61670 20740
rect 62246 20734 62294 20772
rect 62904 20734 62952 20772
rect 61662 20700 61670 20734
rect 61678 20700 62294 20734
rect 62320 20700 62328 20734
rect 62336 20700 62952 20734
rect 61666 20694 61670 20700
rect 62248 20684 62294 20700
rect 62906 20684 62952 20700
rect 62260 20632 62294 20684
rect 62918 20632 62952 20684
rect 62954 20666 62958 20768
rect 63500 20740 63506 21536
rect 63528 20740 63534 21508
rect 63576 20784 63624 22088
rect 63576 20772 63610 20784
rect 62982 20734 62986 20740
rect 63562 20734 63610 20772
rect 62978 20700 62986 20734
rect 62994 20700 63610 20734
rect 62982 20694 62986 20700
rect 63500 20682 63506 20694
rect 63528 20660 63534 20694
rect 63564 20684 63610 20700
rect 63576 20632 63610 20684
rect 63690 20694 63738 22178
rect 64017 22133 64580 22164
rect 63937 21752 63960 22114
rect 63983 22099 64546 22130
rect 63965 21752 63988 22086
rect 64158 21906 64548 21940
rect 64158 21408 64192 21906
rect 64372 21838 64419 21885
rect 64334 21804 64419 21838
rect 64261 21745 64306 21756
rect 64389 21745 64434 21756
rect 64272 21569 64306 21745
rect 64400 21569 64434 21745
rect 64372 21510 64419 21557
rect 64334 21476 64419 21510
rect 64514 21408 64548 21906
rect 64158 21374 64548 21408
rect 60274 20598 63622 20632
rect 63690 20160 63724 20694
rect 63933 20622 63934 20708
rect 63971 20584 63972 20746
rect 64140 20704 64562 21324
rect 60944 14112 60978 20160
rect 73090 15268 73124 16594
rect 73204 15268 73228 15302
rect 64144 15234 64534 15268
rect 72996 15234 73290 15268
rect 64144 14736 64178 15234
rect 64358 15166 64405 15213
rect 64320 15132 64405 15166
rect 64247 15073 64292 15084
rect 64375 15073 64420 15084
rect 64258 14897 64292 15073
rect 64386 14897 64420 15073
rect 64358 14838 64405 14885
rect 64320 14804 64405 14838
rect 64500 14736 64534 15234
rect 73090 15200 73124 15234
rect 73090 15132 73148 15200
rect 73222 15139 73238 15234
rect 73090 14872 73124 15132
rect 73142 14881 73158 15089
rect 73170 15085 73176 15089
rect 73170 15074 73182 15085
rect 73170 15073 73176 15074
rect 73166 14897 73176 15073
rect 73170 14881 73176 14897
rect 73192 14885 73242 15139
rect 73090 14804 73148 14872
rect 73090 14736 73124 14804
rect 73150 14750 73154 14846
rect 73178 14736 73182 14874
rect 73204 14859 73214 14885
rect 73204 14847 73210 14859
rect 73222 14770 73238 14885
rect 73204 14736 73238 14770
rect 73256 14736 73290 15234
rect 105810 15234 106200 15268
rect 64144 14702 64534 14736
rect 72996 14702 73290 14736
rect 73428 14724 73448 15074
rect 105810 14736 105844 15234
rect 106024 15166 106071 15213
rect 105986 15132 106071 15166
rect 105913 15073 105958 15084
rect 106041 15073 106086 15084
rect 105924 14897 105958 15073
rect 106052 14897 106086 15073
rect 106024 14838 106071 14885
rect 105986 14804 106071 14838
rect 106166 14736 106200 15234
rect 105810 14702 106200 14736
rect 73090 14652 73124 14702
rect 64126 14032 64548 14652
rect 73054 14288 73304 14652
rect 73428 14466 73448 14538
rect 73428 14354 73448 14420
rect 73120 14238 73154 14248
rect 73136 14204 73188 14214
rect 73102 14170 73126 14204
rect 73136 14136 73160 14204
rect 73234 14102 73268 14114
rect 73012 14068 73268 14102
rect 105792 14032 106214 14652
rect 37518 13591 38138 13976
rect 38188 13928 38754 13962
rect 38188 13796 38222 13928
rect 38343 13858 38380 13882
rect 38560 13859 38599 13882
rect 38559 13858 38599 13859
rect 38559 13854 38570 13858
rect 38243 13796 38324 13833
rect 38371 13830 38380 13854
rect 38559 13848 38571 13854
rect 38383 13833 38571 13848
rect 38383 13830 38652 13833
rect 38383 13814 38570 13830
rect 38571 13796 38652 13830
rect 38720 13796 38754 13928
rect 38188 13775 38844 13796
rect 38154 13741 38844 13775
rect 38188 13729 38844 13741
rect 38190 13722 38844 13729
rect 38367 13707 38575 13720
rect 38371 13695 38571 13707
rect 38188 13668 38222 13695
rect 38367 13686 38575 13695
rect 38371 13674 38571 13686
rect 38720 13668 38754 13695
rect 114148 13682 114160 13964
rect 114182 13716 114194 13938
rect 38333 13660 38609 13661
rect 38222 13627 38720 13660
rect 38222 13593 38720 13606
<< pdiodelvtc >>
rect 36628 -2808 36736 -2682
<< locali >>
rect 15024 33870 16026 33956
rect 15024 32316 15094 33870
rect 15952 32316 16026 33870
rect 15024 12840 16026 32316
rect 35070 14078 36124 14218
rect 35070 13732 35278 14078
rect 35988 13732 36124 14078
rect 35070 13152 36124 13732
rect 35070 9588 36820 13152
rect 35070 4060 36124 9588
rect 47350 5426 50654 5440
rect 47350 4492 50706 5426
rect 19378 -6684 20292 3040
rect 35048 2518 36128 4060
rect 35048 1920 37074 2518
rect 35048 -6596 36128 1920
rect 40140 -3316 42584 -2318
rect 40140 -3376 42588 -3316
rect 40140 -3494 42590 -3376
rect 41500 -3636 42590 -3494
rect 49206 -5298 50706 4492
rect 18628 -6810 21072 -6684
rect 18628 -7506 18770 -6810
rect 20886 -7506 21072 -6810
rect 18628 -7688 21072 -7506
rect 33864 -6774 37084 -6596
rect 33864 -7668 34260 -6774
rect 36852 -7668 37084 -6774
rect 33864 -7816 37084 -7668
<< viali >>
rect 15094 32316 15952 33870
rect 35278 13732 35988 14078
rect 18770 -7506 20886 -6810
rect 34260 -7668 36852 -6774
<< metal1 >>
rect 15054 33870 16000 33918
rect 15054 32316 15094 33870
rect 15952 32316 16000 33870
rect 15054 32232 16000 32316
rect 22946 32740 24126 32954
rect 22946 32406 23126 32740
rect 23972 32406 24126 32740
rect 22946 31358 24126 32406
rect 46946 32772 48150 32880
rect 46946 32248 47056 32772
rect 48054 32248 48150 32772
rect 22934 22368 24150 23238
rect 22916 13726 24116 14248
rect 34120 14078 36970 31590
rect 46946 31404 48150 32248
rect 46934 21856 48162 23084
rect 34120 13732 35278 14078
rect 35988 13732 36970 14078
rect 22916 13712 33790 13726
rect 22916 13504 33816 13712
rect 34120 13528 36970 13732
rect 33204 13126 33816 13504
rect 33178 12720 34640 13126
rect 47028 12590 48112 14026
rect 23816 4806 24178 5548
rect 22950 2730 24178 4806
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
rect 0 -2400 200 -2200
rect 0 -2800 200 -2600
rect 0 -3200 200 -3000
rect 0 -3600 200 -3400
rect 18628 -6810 21072 -6684
rect 18628 -7506 18770 -6810
rect 20886 -7506 21072 -6810
rect 18628 -7688 21072 -7506
rect 33864 -6774 37084 -6596
rect 33864 -7668 34260 -6774
rect 36852 -7668 37084 -6774
rect 33864 -7816 37084 -7668
<< via1 >>
rect 15094 32316 15952 33870
rect 23126 32406 23972 32740
rect 47056 32248 48054 32772
rect 22222 6310 22362 6456
rect 23548 -2018 23910 -962
rect 18770 -7506 20886 -6810
rect 34260 -7668 36852 -6774
<< metal2 >>
rect 14628 33870 57258 36292
rect 14628 32316 15094 33870
rect 15952 32772 57258 33870
rect 15952 32740 47056 32772
rect 15952 32406 23126 32740
rect 23972 32406 47056 32740
rect 15952 32316 47056 32406
rect 14628 32248 47056 32316
rect 48054 32248 57258 32772
rect 14628 32156 57258 32248
rect 16718 9180 17114 9292
rect 16718 8572 16762 9180
rect 17070 8572 17114 9180
rect 16718 8460 17114 8572
rect 22200 6456 22376 6472
rect 22200 6310 22222 6456
rect 22362 6310 22376 6456
rect 22200 6290 22376 6310
rect 31452 3880 39416 31570
rect 43930 18196 56166 18372
rect 43930 17776 55314 18196
rect 56030 17776 56166 18196
rect 43930 17516 56166 17776
rect 16844 2090 17410 2230
rect 16844 1868 16970 2090
rect 17302 1868 17410 2090
rect 16844 1720 17410 1868
rect 23430 -962 26630 2892
rect 23430 -2018 23548 -962
rect 23910 -2018 26630 -962
rect 23430 -4916 26630 -2018
rect 36202 -2642 36780 3880
rect 22856 -6432 26660 -4916
rect 14582 -6774 57212 -6432
rect 14582 -6810 34260 -6774
rect 14582 -7506 18770 -6810
rect 20886 -7506 34260 -6810
rect 14582 -7668 34260 -7506
rect 36852 -7668 57212 -6774
rect 14582 -10568 57212 -7668
<< via2 >>
rect 30942 27254 31096 27416
rect 26260 23556 27224 24248
rect 30930 18268 31106 18436
rect 26148 14606 27300 15542
rect 16762 8572 17070 9180
rect 25368 8598 25938 9180
rect 27202 8670 27364 8830
rect 21122 6370 21222 6454
rect 22236 6330 22348 6438
rect 39996 27186 40162 27404
rect 44146 27008 44952 27430
rect 39952 17902 40124 18066
rect 55314 17776 56030 18196
rect 40068 8796 40228 8974
rect 44222 8624 45018 9066
rect 16970 1868 17302 2090
rect 27102 -1626 27260 -1470
rect 31500 -1652 31890 -1280
rect 41928 -2498 42036 -2434
rect 37518 -4376 37628 -4258
<< metal3 >>
rect 20550 29986 22164 30292
rect 20550 28896 40436 29986
rect 20550 28632 22164 28896
rect 20572 27644 22186 28072
rect 20572 27416 31334 27644
rect 20572 27254 30942 27416
rect 31096 27254 31334 27416
rect 20572 26824 31334 27254
rect 39788 27404 40430 28896
rect 39788 27186 39996 27404
rect 40162 27186 40430 27404
rect 39788 27068 40430 27186
rect 44044 27430 45012 27488
rect 44044 27008 44146 27430
rect 44952 27008 45012 27430
rect 44044 26942 45012 27008
rect 20572 26412 22186 26824
rect 26150 24248 27368 24346
rect 26150 23556 26260 24248
rect 27224 23556 27368 24248
rect 26150 23446 27368 23556
rect 20594 20878 22208 21304
rect 20594 20000 40506 20878
rect 20594 19644 22208 20000
rect 20616 18664 22230 19130
rect 20616 18436 31258 18664
rect 20616 18268 30930 18436
rect 31106 18268 31258 18436
rect 20616 17856 31258 18268
rect 39654 18066 40490 20000
rect 39654 17902 39952 18066
rect 40124 17902 40490 18066
rect 20616 17470 22230 17856
rect 39654 17780 40490 17902
rect 55248 18196 56070 18248
rect 55248 17776 55314 18196
rect 56030 17776 56070 18196
rect 55248 17704 56070 17776
rect 20616 15340 22230 17000
rect 26094 15542 27478 15704
rect 20932 12410 21958 15340
rect 26094 14606 26148 15542
rect 27300 14606 27478 15542
rect 26094 14498 27478 14606
rect 20932 11616 40604 12410
rect 16744 9180 17092 9258
rect 16744 8572 16762 9180
rect 17070 8572 17092 9180
rect 16744 8506 17092 8572
rect 25252 9180 25996 9236
rect 25252 8598 25368 9180
rect 25938 8598 25996 9180
rect 39810 8974 40588 11616
rect 25252 8518 25996 8598
rect 27126 8830 27436 8888
rect 27126 8670 27202 8830
rect 27364 8670 27436 8830
rect 20890 6454 21304 6548
rect 27126 6498 27436 8670
rect 39810 8796 40068 8974
rect 40228 8796 40588 8974
rect 39810 8628 40588 8796
rect 44166 9066 45096 9160
rect 44166 8624 44222 9066
rect 45018 8624 45096 9066
rect 44166 8552 45096 8624
rect 20890 6370 21122 6454
rect 21222 6370 21304 6454
rect 16844 2090 17410 2230
rect 16844 1868 16970 2090
rect 17302 1868 17410 2090
rect 16844 1720 17410 1868
rect 20890 -902 21304 6370
rect 22180 6438 27460 6498
rect 22180 6330 22236 6438
rect 22348 6330 27460 6438
rect 22180 6258 27460 6330
rect 20636 -1196 21666 -902
rect 31352 -1108 32016 -1102
rect 20636 -1238 22676 -1196
rect 20636 -1848 22884 -1238
rect 24072 -1470 27316 -1238
rect 24072 -1626 27102 -1470
rect 27260 -1626 27316 -1470
rect 24072 -1848 27316 -1626
rect 31352 -1280 32018 -1108
rect 31352 -1652 31500 -1280
rect 31890 -1652 32018 -1280
rect 20636 -1924 22676 -1848
rect 31352 -1894 32018 -1652
rect 31368 -1896 32018 -1894
rect 20636 -2074 21666 -1924
rect 41868 -2234 42188 -2158
rect 41868 -2552 41898 -2234
rect 42136 -2552 42188 -2234
rect 41868 -2564 42188 -2552
rect 35964 -4114 37728 -4064
rect 35954 -4258 37728 -4114
rect 35954 -4376 37518 -4258
rect 37628 -4376 37728 -4258
rect 35954 -4586 37728 -4376
rect 35658 -4606 37728 -4586
rect 35658 -5760 36862 -4606
<< via3 >>
rect 44146 27008 44952 27430
rect 26260 23556 27224 24248
rect 55362 17824 55974 18154
rect 26148 14606 27300 15542
rect 16792 8698 17056 9048
rect 25490 8630 25844 9028
rect 44222 8624 45018 9066
rect 41898 -2434 42136 -2234
rect 41898 -2498 41928 -2434
rect 41928 -2498 42036 -2434
rect 42036 -2498 42136 -2434
rect 41898 -2552 42136 -2498
<< metal4 >>
rect 43928 27430 50272 27584
rect 43928 27008 44146 27430
rect 44952 27008 50272 27430
rect 43928 26774 50272 27008
rect 26058 24248 50282 24536
rect 26058 23556 26260 24248
rect 27224 23556 50282 24248
rect 26058 23260 50282 23556
rect 54812 18154 57228 31570
rect 54772 17824 55362 18154
rect 55974 17824 57228 18154
rect 16328 15236 18180 17016
rect 25976 15542 50196 15820
rect 16720 9332 17814 15236
rect 25976 14606 26148 15542
rect 27300 14606 50196 15542
rect 25976 14396 50196 14606
rect 16682 9048 26064 9332
rect 16682 8698 16792 9048
rect 17056 9028 26064 9048
rect 17056 8698 25490 9028
rect 16682 8630 25490 8698
rect 25844 8630 26064 9028
rect 16682 8386 26064 8630
rect 44038 9066 50258 9232
rect 44038 8624 44222 9066
rect 45018 8624 50258 9066
rect 44038 8436 50258 8624
rect 54812 6018 57228 17824
rect 54834 1498 57198 6018
rect 53568 1454 57198 1498
rect 46982 1092 57198 1454
rect 46982 1082 54970 1092
rect 53568 1048 54970 1082
rect 31368 -1646 42344 -1066
rect 31368 -1868 42348 -1646
rect 41794 -2234 42348 -1868
rect 41794 -2552 41898 -2234
rect 42136 -2552 42348 -2234
rect 41794 -2600 42348 -2552
use curr_mir  curr_mir_0
timestamp 1695698273
transform 1 0 72116 0 1 7240
box 0 -400 11334 10390
use not  not_0
timestamp 1695698273
transform 1 0 20522 0 1 6220
box 0 -578 1868 990
use opamp  opamp_0
timestamp 1695698273
transform 1 0 77382 0 1 11126
box 0 -1200 19288 9014
use switch  switch_0
timestamp 1695698273
transform 1 0 55118 0 1 13320
box -114 -950 10034 11418
use switch  switch_1
timestamp 1695698273
transform 1 0 63874 0 1 13320
box -114 -950 10034 11418
use switch  switch_2
timestamp 1695698273
transform 1 0 96784 0 1 13320
box -114 -950 10034 11418
use switch  switch_3
timestamp 1695698273
transform 1 0 105540 0 1 13320
box -114 -950 10034 11418
use switch  switch_4
timestamp 1695698273
transform 1 0 115688 0 1 13320
box -114 -950 10034 11418
use switch  switch_5
timestamp 1695698273
transform 1 0 55132 0 1 19992
box -114 -950 10034 11418
use switch  switch_6
timestamp 1695698273
transform 1 0 55164 0 1 26356
box -114 -950 10034 11418
use switch  x1
timestamp 1695698273
transform 0 1 36806 1 0 4546
box -114 -950 10034 11418
use switch  x2
timestamp 1695698273
transform 0 1 23934 -1 0 13086
box -114 -950 10034 11418
use curr_mir  x3
timestamp 1695698273
transform 0 -1 25426 1 0 1738
box 0 -400 11334 10390
use opamp  x4
timestamp 1695698273
transform 1 0 30358 0 -1 3752
box 0 -1200 19288 9014
use switch  x5
timestamp 1695698273
transform 0 1 36696 1 0 13644
box -114 -950 10034 11418
use switch  x6
timestamp 1695698273
transform 0 1 23834 -1 0 2788
box -114 -950 10034 11418
use not  x7
timestamp 1695698273
transform 1 0 113706 0 1 12948
box 0 -578 1868 990
use switch  x8
timestamp 1695698273
transform 0 1 36738 1 0 22948
box -114 -950 10034 11418
use switch  x9
timestamp 1695698273
transform 0 -1 34358 1 0 14018
box -114 -950 10034 11418
use switch  x10
timestamp 1695698273
transform 0 -1 34358 1 0 22992
box -114 -950 10034 11418
use sky130_fd_pr__cap_mim_m3_1_3HBNLG  XC1
timestamp 1695395215
transform 1 0 51818 0 1 9140
box -3186 -3040 3186 3040
use sky130_fd_pr__cap_mim_m3_1_3HBNLG  XC2
timestamp 1695395215
transform 1 0 51818 0 1 15410
box -3186 -3040 3186 3040
use sky130_fd_pr__cap_mim_m3_1_3HBNLG  XC3
timestamp 1695395215
transform 1 0 51832 0 1 22082
box -3186 -3040 3186 3040
use sky130_fd_pr__cap_mim_m3_1_3HBNLG  XC4
timestamp 1695395215
transform 1 0 51864 0 1 28446
box -3186 -3040 3186 3040
<< labels >>
rlabel metal4 54834 1092 57198 17824 1 intout
port 7 nsew
rlabel metal3 20550 28632 22164 30292 1 sw4
port 8 nsew
rlabel metal3 20572 26412 22186 28072 1 sw3
port 9 nsew
rlabel metal3 20594 19644 22208 21304 1 rst
port 10 nsew
rlabel metal3 20616 17470 22230 19130 1 sw2
port 11 nsew
rlabel metal3 20616 15340 22230 17000 1 sw1
port 12 nsew
rlabel metal3 35658 -5760 36862 -4586 1 opbias
port 13 nsew
rlabel metal3 20636 -2074 21666 -902 1 en
port 14 nsew
rlabel metal3 16844 1720 17410 2230 1 Vtune
port 15 nsew
rlabel metal4 16328 15236 18180 17016 1 intin
port 16 nsew
rlabel metal2 14628 32156 57258 36292 1 VDD
port 17 nsew
rlabel metal2 14582 -10568 57212 -6432 1 GROUND
port 18 nsew
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 sw2
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 sw1
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 intin
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 intout
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 opbias
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 en
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 256 0 0 0 Vtune
port 6 nsew
flabel metal1 0 -2800 200 -2600 0 FreeSans 256 0 0 0 rst
flabel metal1 0 -3200 200 -3000 0 FreeSans 256 0 0 0 sw4
flabel metal1 0 -3600 200 -3400 0 FreeSans 256 0 0 0 sw3
<< end >>
