magic
tech sky130A
timestamp 1695803704
<< metal1 >>
rect 3660 5583 9473 5591
rect 3660 5461 9480 5583
rect 3663 5287 9480 5461
rect 3265 4979 3365 4986
rect 3265 4898 3277 4979
rect 3357 4898 3365 4979
rect 3265 4886 3365 4898
rect 2815 3854 2915 3865
rect 2815 3778 2833 3854
rect 2906 3778 2915 3854
rect 2815 3765 2915 3778
rect 8930 1863 9030 1866
rect 8927 1770 8932 1863
rect 9027 1770 9032 1863
rect 8930 1766 9030 1770
rect 3138 1278 7659 1734
rect 3092 1165 7692 1278
rect 3138 1163 7659 1165
<< via1 >>
rect 3277 4898 3357 4979
rect 2833 3778 2906 3854
rect 8932 1770 9027 1863
<< metal2 >>
rect 3184 5108 3446 5154
rect 3184 4780 3224 5108
rect 3415 4983 3446 5108
rect 3415 4892 3651 4983
rect 3415 4780 3446 4892
rect 3184 4728 3446 4780
rect 2926 4055 3020 4056
rect 2926 3963 3128 4055
rect 5778 4036 5849 4041
rect 2823 3854 2911 3863
rect 2823 3778 2833 3854
rect 2906 3778 2911 3854
rect 2823 3770 2911 3778
rect 2926 1625 3020 3963
rect 5778 3960 5849 3965
rect 2925 1431 3020 1625
rect 8328 1866 8430 2189
rect 8932 1866 9027 1868
rect 8328 1863 9030 1866
rect 8328 1770 8932 1863
rect 9027 1770 9030 1863
rect 8328 1766 9030 1770
rect 8328 1431 8430 1766
rect 8932 1765 9027 1766
rect 2925 1340 8430 1431
rect 2925 1339 8262 1340
<< via2 >>
rect 3224 4979 3415 5108
rect 3224 4898 3277 4979
rect 3277 4898 3357 4979
rect 3357 4898 3415 4979
rect 3224 4780 3415 4898
rect 5778 3965 5849 4036
rect 2833 3778 2906 3854
<< metal3 >>
rect 3126 5108 3494 5186
rect 3126 4780 3224 5108
rect 3415 4780 3494 5108
rect 3126 4693 3494 4780
rect 5769 4036 5861 4053
rect 5769 3965 5778 4036
rect 5849 3965 5861 4036
rect 5769 3961 5861 3965
rect 2820 3854 2912 3864
rect 2820 3778 2833 3854
rect 2906 3778 2912 3854
rect 2820 3768 2912 3778
<< via3 >>
rect 5778 3965 5849 4036
rect 2833 3778 2906 3854
<< metal4 >>
rect 5775 4036 5866 4047
rect 5775 3965 5778 4036
rect 5849 3965 5866 4036
rect 5775 3861 5866 3965
rect 2824 3854 5866 3861
rect 2824 3778 2833 3854
rect 2906 3778 5866 3854
rect 2824 3764 5866 3778
use opamp  x1
timestamp 1695803704
transform 1 0 0 0 1 900
box 3034 622 9644 4507
<< labels >>
flabel metal1 2815 3765 2915 3865 0 FreeSans 128 0 0 0 in
port 1 nsew
flabel metal1 3265 4886 3365 4986 0 FreeSans 128 0 0 0 opbias
port 0 nsew
flabel metal1 8930 1766 9030 1866 0 FreeSans 128 0 0 0 out
port 2 nsew
rlabel metal1 3660 5461 9473 5591 1 VDD
port 3 nsew
rlabel metal1 3092 1165 7692 1278 1 GROUND
port 4 nsew
<< end >>
