magic
tech sky130A
magscale 1 2
timestamp 1695378092
<< nwell >>
rect -1483 -469 1483 469
<< pmoslvt >>
rect -1287 -250 -687 250
rect -629 -250 -29 250
rect 29 -250 629 250
rect 687 -250 1287 250
<< pdiff >>
rect -1345 238 -1287 250
rect -1345 -238 -1333 238
rect -1299 -238 -1287 238
rect -1345 -250 -1287 -238
rect -687 238 -629 250
rect -687 -238 -675 238
rect -641 -238 -629 238
rect -687 -250 -629 -238
rect -29 238 29 250
rect -29 -238 -17 238
rect 17 -238 29 238
rect -29 -250 29 -238
rect 629 238 687 250
rect 629 -238 641 238
rect 675 -238 687 238
rect 629 -250 687 -238
rect 1287 238 1345 250
rect 1287 -238 1299 238
rect 1333 -238 1345 238
rect 1287 -250 1345 -238
<< pdiffc >>
rect -1333 -238 -1299 238
rect -675 -238 -641 238
rect -17 -238 17 238
rect 641 -238 675 238
rect 1299 -238 1333 238
<< nsubdiff >>
rect -1447 399 -1351 433
rect 1351 399 1447 433
rect -1447 337 -1413 399
rect 1413 337 1447 399
rect -1447 -399 -1413 -337
rect 1413 -399 1447 -337
rect -1447 -433 -1351 -399
rect 1351 -433 1447 -399
<< nsubdiffcont >>
rect -1351 399 1351 433
rect -1447 -337 -1413 337
rect 1413 -337 1447 337
rect -1351 -433 1351 -399
<< poly >>
rect -1287 331 -687 347
rect -1287 297 -1271 331
rect -703 297 -687 331
rect -1287 250 -687 297
rect -629 331 -29 347
rect -629 297 -613 331
rect -45 297 -29 331
rect -629 250 -29 297
rect 29 331 629 347
rect 29 297 45 331
rect 613 297 629 331
rect 29 250 629 297
rect 687 331 1287 347
rect 687 297 703 331
rect 1271 297 1287 331
rect 687 250 1287 297
rect -1287 -297 -687 -250
rect -1287 -331 -1271 -297
rect -703 -331 -687 -297
rect -1287 -347 -687 -331
rect -629 -297 -29 -250
rect -629 -331 -613 -297
rect -45 -331 -29 -297
rect -629 -347 -29 -331
rect 29 -297 629 -250
rect 29 -331 45 -297
rect 613 -331 629 -297
rect 29 -347 629 -331
rect 687 -297 1287 -250
rect 687 -331 703 -297
rect 1271 -331 1287 -297
rect 687 -347 1287 -331
<< polycont >>
rect -1271 297 -703 331
rect -613 297 -45 331
rect 45 297 613 331
rect 703 297 1271 331
rect -1271 -331 -703 -297
rect -613 -331 -45 -297
rect 45 -331 613 -297
rect 703 -331 1271 -297
<< locali >>
rect -1447 399 -1351 433
rect 1351 399 1447 433
rect -1447 337 -1413 399
rect 1413 337 1447 399
rect -1287 297 -1271 331
rect -703 297 -687 331
rect -629 297 -613 331
rect -45 297 -29 331
rect 29 297 45 331
rect 613 297 629 331
rect 687 297 703 331
rect 1271 297 1287 331
rect -1333 238 -1299 254
rect -1333 -254 -1299 -238
rect -675 238 -641 254
rect -675 -254 -641 -238
rect -17 238 17 254
rect -17 -254 17 -238
rect 641 238 675 254
rect 641 -254 675 -238
rect 1299 238 1333 254
rect 1299 -254 1333 -238
rect -1287 -331 -1271 -297
rect -703 -331 -687 -297
rect -629 -331 -613 -297
rect -45 -331 -29 -297
rect 29 -331 45 -297
rect 613 -331 629 -297
rect 687 -331 703 -297
rect 1271 -331 1287 -297
rect -1447 -399 -1413 -337
rect 1413 -399 1447 -337
rect -1447 -433 -1351 -399
rect 1351 -433 1447 -399
<< viali >>
rect -1271 297 -703 331
rect -613 297 -45 331
rect 45 297 613 331
rect 703 297 1271 331
rect -1333 -238 -1299 238
rect -675 -238 -641 238
rect -17 -238 17 238
rect 641 -238 675 238
rect 1299 -238 1333 238
rect -1271 -331 -703 -297
rect -613 -331 -45 -297
rect 45 -331 613 -297
rect 703 -331 1271 -297
<< metal1 >>
rect -1283 331 -691 337
rect -1283 297 -1271 331
rect -703 297 -691 331
rect -1283 291 -691 297
rect -625 331 -33 337
rect -625 297 -613 331
rect -45 297 -33 331
rect -625 291 -33 297
rect 33 331 625 337
rect 33 297 45 331
rect 613 297 625 331
rect 33 291 625 297
rect 691 331 1283 337
rect 691 297 703 331
rect 1271 297 1283 331
rect 691 291 1283 297
rect -1339 238 -1293 250
rect -1339 -238 -1333 238
rect -1299 -238 -1293 238
rect -1339 -250 -1293 -238
rect -681 238 -635 250
rect -681 -238 -675 238
rect -641 -238 -635 238
rect -681 -250 -635 -238
rect -23 238 23 250
rect -23 -238 -17 238
rect 17 -238 23 238
rect -23 -250 23 -238
rect 635 238 681 250
rect 635 -238 641 238
rect 675 -238 681 238
rect 635 -250 681 -238
rect 1293 238 1339 250
rect 1293 -238 1299 238
rect 1333 -238 1339 238
rect 1293 -250 1339 -238
rect -1283 -297 -691 -291
rect -1283 -331 -1271 -297
rect -703 -331 -691 -297
rect -1283 -337 -691 -331
rect -625 -297 -33 -291
rect -625 -331 -613 -297
rect -45 -331 -33 -297
rect -625 -337 -33 -331
rect 33 -297 625 -291
rect 33 -331 45 -297
rect 613 -331 625 -297
rect 33 -337 625 -331
rect 691 -297 1283 -291
rect 691 -331 703 -297
rect 1271 -331 1283 -297
rect 691 -337 1283 -331
<< labels >>
rlabel poly -1287 250 -687 297 1 G
rlabel locali -1333 238 -1299 254 1 D
rlabel locali -675 238 -641 254 1 S
rlabel nsubdiffcont -1351 399 1351 433 1 B
<< properties >>
string FIXED_BBOX -1430 -416 1430 416
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 2.5 l 3.0 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
