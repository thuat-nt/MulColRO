magic
tech sky130A
magscale 1 2
timestamp 1695441144
<< nwell >>
rect -1812 -2219 1812 2219
<< pmoslvt >>
rect -1616 -2000 -1016 2000
rect -958 -2000 -358 2000
rect -300 -2000 300 2000
rect 358 -2000 958 2000
rect 1016 -2000 1616 2000
<< pdiff >>
rect -1674 1988 -1616 2000
rect -1674 -1988 -1662 1988
rect -1628 -1988 -1616 1988
rect -1674 -2000 -1616 -1988
rect -1016 1988 -958 2000
rect -1016 -1988 -1004 1988
rect -970 -1988 -958 1988
rect -1016 -2000 -958 -1988
rect -358 1988 -300 2000
rect -358 -1988 -346 1988
rect -312 -1988 -300 1988
rect -358 -2000 -300 -1988
rect 300 1988 358 2000
rect 300 -1988 312 1988
rect 346 -1988 358 1988
rect 300 -2000 358 -1988
rect 958 1988 1016 2000
rect 958 -1988 970 1988
rect 1004 -1988 1016 1988
rect 958 -2000 1016 -1988
rect 1616 1988 1674 2000
rect 1616 -1988 1628 1988
rect 1662 -1988 1674 1988
rect 1616 -2000 1674 -1988
<< pdiffc >>
rect -1662 -1988 -1628 1988
rect -1004 -1988 -970 1988
rect -346 -1988 -312 1988
rect 312 -1988 346 1988
rect 970 -1988 1004 1988
rect 1628 -1988 1662 1988
<< nsubdiff >>
rect -1776 2149 -1680 2183
rect 1680 2149 1776 2183
rect -1776 2087 -1742 2149
rect 1742 2087 1776 2149
rect -1776 -2149 -1742 -2087
rect 1742 -2149 1776 -2087
rect -1776 -2183 -1680 -2149
rect 1680 -2183 1776 -2149
<< nsubdiffcont >>
rect -1680 2149 1680 2183
rect -1776 -2087 -1742 2087
rect 1742 -2087 1776 2087
rect -1680 -2183 1680 -2149
<< poly >>
rect -1616 2081 -1016 2097
rect -1616 2047 -1600 2081
rect -1032 2047 -1016 2081
rect -1616 2000 -1016 2047
rect -958 2081 -358 2097
rect -958 2047 -942 2081
rect -374 2047 -358 2081
rect -958 2000 -358 2047
rect -300 2081 300 2097
rect -300 2047 -284 2081
rect 284 2047 300 2081
rect -300 2000 300 2047
rect 358 2081 958 2097
rect 358 2047 374 2081
rect 942 2047 958 2081
rect 358 2000 958 2047
rect 1016 2081 1616 2097
rect 1016 2047 1032 2081
rect 1600 2047 1616 2081
rect 1016 2000 1616 2047
rect -1616 -2047 -1016 -2000
rect -1616 -2081 -1600 -2047
rect -1032 -2081 -1016 -2047
rect -1616 -2097 -1016 -2081
rect -958 -2047 -358 -2000
rect -958 -2081 -942 -2047
rect -374 -2081 -358 -2047
rect -958 -2097 -358 -2081
rect -300 -2047 300 -2000
rect -300 -2081 -284 -2047
rect 284 -2081 300 -2047
rect -300 -2097 300 -2081
rect 358 -2047 958 -2000
rect 358 -2081 374 -2047
rect 942 -2081 958 -2047
rect 358 -2097 958 -2081
rect 1016 -2047 1616 -2000
rect 1016 -2081 1032 -2047
rect 1600 -2081 1616 -2047
rect 1016 -2097 1616 -2081
<< polycont >>
rect -1600 2047 -1032 2081
rect -942 2047 -374 2081
rect -284 2047 284 2081
rect 374 2047 942 2081
rect 1032 2047 1600 2081
rect -1600 -2081 -1032 -2047
rect -942 -2081 -374 -2047
rect -284 -2081 284 -2047
rect 374 -2081 942 -2047
rect 1032 -2081 1600 -2047
<< locali >>
rect -1776 2149 -1680 2183
rect 1680 2149 1776 2183
rect -1776 2087 -1742 2149
rect 1742 2087 1776 2149
rect -1616 2047 -1600 2081
rect -1032 2047 -1016 2081
rect -958 2047 -942 2081
rect -374 2047 -358 2081
rect -300 2047 -284 2081
rect 284 2047 300 2081
rect 358 2047 374 2081
rect 942 2047 958 2081
rect 1016 2047 1032 2081
rect 1600 2047 1616 2081
rect -1662 1988 -1628 2004
rect -1662 -2004 -1628 -1988
rect -1004 1988 -970 2004
rect -1004 -2004 -970 -1988
rect -346 1988 -312 2004
rect -346 -2004 -312 -1988
rect 312 1988 346 2004
rect 312 -2004 346 -1988
rect 970 1988 1004 2004
rect 970 -2004 1004 -1988
rect 1628 1988 1662 2004
rect 1628 -2004 1662 -1988
rect -1616 -2081 -1600 -2047
rect -1032 -2081 -1016 -2047
rect -958 -2081 -942 -2047
rect -374 -2081 -358 -2047
rect -300 -2081 -284 -2047
rect 284 -2081 300 -2047
rect 358 -2081 374 -2047
rect 942 -2081 958 -2047
rect 1016 -2081 1032 -2047
rect 1600 -2081 1616 -2047
rect -1776 -2149 -1742 -2087
rect 1742 -2149 1776 -2087
rect -1776 -2183 -1680 -2149
rect 1680 -2183 1776 -2149
<< viali >>
rect -1600 2047 -1032 2081
rect -942 2047 -374 2081
rect -284 2047 284 2081
rect 374 2047 942 2081
rect 1032 2047 1600 2081
rect -1662 -1988 -1628 1988
rect -1004 -1988 -970 1988
rect -346 -1988 -312 1988
rect 312 -1988 346 1988
rect 970 -1988 1004 1988
rect 1628 -1988 1662 1988
rect -1600 -2081 -1032 -2047
rect -942 -2081 -374 -2047
rect -284 -2081 284 -2047
rect 374 -2081 942 -2047
rect 1032 -2081 1600 -2047
<< metal1 >>
rect -1612 2081 -1020 2087
rect -1612 2047 -1600 2081
rect -1032 2047 -1020 2081
rect -1612 2041 -1020 2047
rect -954 2081 -362 2087
rect -954 2047 -942 2081
rect -374 2047 -362 2081
rect -954 2041 -362 2047
rect -296 2081 296 2087
rect -296 2047 -284 2081
rect 284 2047 296 2081
rect -296 2041 296 2047
rect 362 2081 954 2087
rect 362 2047 374 2081
rect 942 2047 954 2081
rect 362 2041 954 2047
rect 1020 2081 1612 2087
rect 1020 2047 1032 2081
rect 1600 2047 1612 2081
rect 1020 2041 1612 2047
rect -1668 1988 -1622 2000
rect -1668 -1988 -1662 1988
rect -1628 -1988 -1622 1988
rect -1668 -2000 -1622 -1988
rect -1010 1988 -964 2000
rect -1010 -1988 -1004 1988
rect -970 -1988 -964 1988
rect -1010 -2000 -964 -1988
rect -352 1988 -306 2000
rect -352 -1988 -346 1988
rect -312 -1988 -306 1988
rect -352 -2000 -306 -1988
rect 306 1988 352 2000
rect 306 -1988 312 1988
rect 346 -1988 352 1988
rect 306 -2000 352 -1988
rect 964 1988 1010 2000
rect 964 -1988 970 1988
rect 1004 -1988 1010 1988
rect 964 -2000 1010 -1988
rect 1622 1988 1668 2000
rect 1622 -1988 1628 1988
rect 1662 -1988 1668 1988
rect 1622 -2000 1668 -1988
rect -1612 -2047 -1020 -2041
rect -1612 -2081 -1600 -2047
rect -1032 -2081 -1020 -2047
rect -1612 -2087 -1020 -2081
rect -954 -2047 -362 -2041
rect -954 -2081 -942 -2047
rect -374 -2081 -362 -2047
rect -954 -2087 -362 -2081
rect -296 -2047 296 -2041
rect -296 -2081 -284 -2047
rect 284 -2081 296 -2047
rect -296 -2087 296 -2081
rect 362 -2047 954 -2041
rect 362 -2081 374 -2047
rect 942 -2081 954 -2047
rect 362 -2087 954 -2081
rect 1020 -2047 1612 -2041
rect 1020 -2081 1032 -2047
rect 1600 -2081 1612 -2047
rect 1020 -2087 1612 -2081
<< labels >>
rlabel locali -1004 1988 -970 2004 1 S
rlabel poly -1616 2000 -1016 2047 1 G
rlabel locali -1662 1988 -1628 2004 1 D
<< properties >>
string FIXED_BBOX -1759 -2166 1759 2166
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 20.0 l 3.0 m 1 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
