magic
tech sky130A
magscale 1 2
timestamp 1695461801
<< metal3 >>
rect -56 31 56 88
rect -56 -88 56 -31
<< rmetal3 >>
rect -56 -31 56 31
<< properties >>
string gencell sky130_fd_pr__res_generic_m3
string library sky130
string parameters w 0.56 l 0.31 m 1 nx 1 wmin 0.30 lmin 0.30 rho 0.047 val 26.017m dummy 0 dw 0.0 term 0.0 roverlap 0
<< end >>
