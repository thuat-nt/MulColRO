magic
tech sky130A
magscale 1 2
timestamp 1695698273
<< metal3 >>
rect -1100 30 1100 87
rect -1100 -87 1100 -30
<< rmetal3 >>
rect -1100 -30 1100 30
<< properties >>
string gencell sky130_fd_pr__res_generic_m3
string library sky130
string parameters w 11.0 l 0.30 m 1 nx 1 wmin 0.30 lmin 0.30 rho 0.047 val 1.068m dummy 0 dw 0.0 term 0.0 roverlap 0
<< end >>
