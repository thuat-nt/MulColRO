magic
tech sky130A
magscale 1 2
timestamp 1695455187
<< locali >>
rect 2 10670 3680 10764
rect 2 10298 2458 10670
rect 3162 10298 3680 10670
rect 2 10018 3680 10298
rect -22 8912 3738 10018
rect 5052 116 8620 644
rect 5052 -204 5758 116
rect 6200 -186 8620 116
rect 6200 -204 8634 -186
rect 5052 -268 8634 -204
rect 5130 -456 6902 -268
rect 8226 -284 8634 -268
rect 8276 -294 8634 -284
<< viali >>
rect 2458 10298 3162 10670
rect 5758 -204 6200 116
<< metal1 >>
rect -44 10670 8600 11418
rect -44 10298 2458 10670
rect 3162 10298 8600 10670
rect -44 10230 8600 10298
rect 214 4956 662 8866
rect 712 7938 840 8460
rect 712 7482 738 7938
rect 808 7482 840 7938
rect 712 7108 840 7482
rect 214 4508 316 4956
rect 528 4508 662 4956
rect 64 2148 172 2504
rect 64 1494 78 2148
rect 152 1494 172 2148
rect 64 1102 172 1494
rect 214 672 662 4508
rect 872 4948 1320 8850
rect 872 4500 992 4948
rect 1204 4500 1320 4948
rect 872 656 1320 4500
rect 1534 4956 1982 8866
rect 2022 7922 2150 8466
rect 2022 7466 2050 7922
rect 2120 7466 2150 7922
rect 2022 7114 2150 7466
rect 1534 4508 1638 4956
rect 1850 4508 1982 4956
rect 1372 2148 1480 2492
rect 1372 1494 1392 2148
rect 1466 1494 1480 2148
rect 1372 1090 1480 1494
rect 1534 672 1982 4508
rect 2204 4948 2652 8866
rect 2204 4500 2334 4948
rect 2546 4500 2652 4948
rect 2204 672 2652 4500
rect 2856 4948 3304 8866
rect 3344 7900 3472 8436
rect 3344 7444 3372 7900
rect 3442 7444 3472 7900
rect 4202 7920 4402 7948
rect 4202 7784 4238 7920
rect 4374 7784 4402 7920
rect 4202 7748 4402 7784
rect 3344 7084 3472 7444
rect 4802 5398 4940 10230
rect 2856 4500 2980 4948
rect 3192 4500 3304 4948
rect 5300 4928 5748 8890
rect 5782 7838 5918 8204
rect 5782 7380 5800 7838
rect 5892 7380 5918 7838
rect 5782 7100 5918 7380
rect 2692 2128 2800 2470
rect 2692 1474 2708 2128
rect 2782 1474 2800 2128
rect 2692 1068 2800 1474
rect 2856 672 3304 4500
rect 5300 4480 5412 4928
rect 5624 4480 5748 4928
rect 4228 3404 4428 3444
rect 4228 3282 4284 3404
rect 4402 3282 4428 3404
rect 4228 3244 4428 3282
rect 4238 1818 4438 1844
rect 4238 1664 4264 1818
rect 4418 1664 4438 1818
rect 4238 1644 4438 1664
rect 4804 238 4942 4464
rect 5132 2164 5240 2478
rect 5132 1510 5152 2164
rect 5226 1510 5240 2164
rect 5132 1076 5240 1510
rect 5300 696 5748 4480
rect 5952 4924 6400 8894
rect 5952 4476 6078 4924
rect 6290 4476 6400 4924
rect 5952 808 6400 4476
rect 6610 4928 7058 8890
rect 7102 7810 7238 8186
rect 7102 7352 7118 7810
rect 7210 7352 7238 7810
rect 7102 7082 7238 7352
rect 6610 4480 6726 4928
rect 6938 4480 7058 4928
rect 6442 2136 6550 2484
rect 6442 1482 6466 2136
rect 6540 1482 6550 2136
rect 6442 1082 6550 1482
rect 6610 696 7058 4480
rect 7274 4922 7722 8878
rect 7274 4474 7394 4922
rect 7606 4474 7722 4922
rect 7274 684 7722 4474
rect 7926 4910 8374 8884
rect 8410 7798 8546 8188
rect 8410 7340 8434 7798
rect 8526 7340 8546 7798
rect 8410 7084 8546 7340
rect 7926 4462 8038 4910
rect 8250 4462 8374 4910
rect 7764 2128 7872 2448
rect 7764 1474 7782 2128
rect 7856 1474 7872 2128
rect 7764 1046 7872 1474
rect 7926 690 8374 4462
rect -114 116 8274 238
rect -114 -204 5758 116
rect 6200 10 8274 116
rect 6200 -200 8530 10
rect 6200 -204 8284 -200
rect -114 -308 8284 -204
rect -114 -950 8530 -308
<< via1 >>
rect 738 7482 808 7938
rect 316 4508 528 4956
rect 78 1494 152 2148
rect 992 4500 1204 4948
rect 2050 7466 2120 7922
rect 1638 4508 1850 4956
rect 1392 1494 1466 2148
rect 2334 4500 2546 4948
rect 3372 7444 3442 7900
rect 4238 7784 4374 7920
rect 2980 4500 3192 4948
rect 5800 7380 5892 7838
rect 3636 4724 3754 4856
rect 2708 1474 2782 2128
rect 5412 4480 5624 4928
rect 4284 3282 4402 3404
rect 4264 1664 4418 1818
rect 5152 1510 5226 2164
rect 6078 4476 6290 4924
rect 7118 7352 7210 7810
rect 6726 4480 6938 4928
rect 6466 1482 6540 2136
rect 7394 4474 7606 4922
rect 8434 7340 8526 7798
rect 8038 4462 8250 4910
rect 7782 1474 7856 2128
<< metal2 >>
rect 42 8352 3478 8718
rect 5116 8352 8552 8740
rect 42 7938 8552 8352
rect 42 7482 738 7938
rect 808 7922 8552 7938
rect 808 7482 2050 7922
rect 42 7466 2050 7482
rect 2120 7920 8552 7922
rect 2120 7900 4238 7920
rect 2120 7466 3372 7900
rect 42 7444 3372 7466
rect 3442 7784 4238 7900
rect 4374 7838 8552 7920
rect 4374 7784 5800 7838
rect 3442 7444 5800 7784
rect 42 7380 5800 7444
rect 5892 7810 8552 7838
rect 5892 7380 7118 7810
rect 42 7352 7118 7380
rect 7210 7798 8552 7810
rect 7210 7352 8434 7798
rect 42 7340 8434 7352
rect 8526 7340 8552 7798
rect 42 7226 8552 7340
rect 42 6772 3478 7226
rect 5116 6794 8552 7226
rect 52 4956 3470 5178
rect 52 4508 316 4956
rect 528 4948 1638 4956
rect 528 4508 992 4948
rect 52 4500 992 4508
rect 1204 4508 1638 4948
rect 1850 4948 3470 4956
rect 1850 4508 2334 4948
rect 1204 4500 2334 4508
rect 2546 4500 2980 4948
rect 3192 4904 3470 4948
rect 5126 4928 8544 5168
rect 5126 4914 5412 4928
rect 3192 4856 3796 4904
rect 3192 4724 3636 4856
rect 3754 4724 3796 4856
rect 3192 4668 3796 4724
rect 4744 4684 5412 4914
rect 3192 4500 3470 4668
rect 52 4264 3470 4500
rect 5126 4480 5412 4684
rect 5624 4924 6726 4928
rect 5624 4480 6078 4924
rect 5126 4476 6078 4480
rect 6290 4480 6726 4924
rect 6938 4922 8544 4928
rect 6938 4480 7394 4922
rect 6290 4476 7394 4480
rect 5126 4474 7394 4476
rect 7606 4910 8544 4922
rect 7606 4474 8038 4910
rect 5126 4462 8038 4474
rect 8250 4462 8544 4910
rect 5126 4254 8544 4462
rect 5126 3474 5310 4254
rect 4218 3404 5310 3474
rect 4218 3282 4284 3404
rect 4402 3282 5310 3404
rect 4218 3220 5310 3282
rect 4218 3216 5270 3220
rect 34 2336 3470 2756
rect 5112 2336 8548 2746
rect 34 2164 8548 2336
rect 34 2148 5152 2164
rect 34 1494 78 2148
rect 152 1494 1392 2148
rect 1466 2128 5152 2148
rect 1466 1494 2708 2128
rect 34 1474 2708 1494
rect 2782 1818 5152 2128
rect 2782 1664 4264 1818
rect 4418 1664 5152 1818
rect 2782 1510 5152 1664
rect 5226 2136 8548 2164
rect 5226 1510 6466 2136
rect 2782 1482 6466 1510
rect 6540 2128 8548 2136
rect 6540 1482 7782 2128
rect 2782 1474 7782 1482
rect 7856 1474 8548 2128
rect 34 1210 8548 1474
rect 34 810 3470 1210
rect 5112 808 8548 1210
rect 5112 800 5802 808
rect 6520 800 8548 808
use not  x1
timestamp 1695395215
transform -1 0 5462 0 1 4624
box 476 -578 1868 990
use sky130_fd_pr__nfet_01v8_lvt_4833E6  XM1
timestamp 1695367880
transform 1 0 6830 0 1 4780
box -1812 -4210 1812 4210
use sky130_fd_pr__pfet_01v8_lvt_RMWXAE  XM10
timestamp 1695367880
transform 1 0 1759 0 1 4766
box -1812 -4219 1812 4219
<< labels >>
flabel metal1 4238 1644 4438 1844 0 FreeSans 256 0 0 0 in
port 2 nsew
flabel metal1 4202 7748 4402 7948 0 FreeSans 256 0 0 0 out
port 1 nsew
rlabel via1 4284 3282 4402 3404 1 toggle
port 6 nsew
rlabel metal1 -44 10230 8600 11418 1 VDD
port 4 nsew
rlabel space -114 -950 8530 238 1 GROUND
port 5 nsew
rlabel metal1 2416 -750 3238 -114 1 GROUND
<< end >>
