magic
tech sky130A
magscale 1 2
timestamp 1695698600
<< error_p >>
rect 161373 630858 161407 636816
rect 158627 630551 158661 630858
rect 158741 630647 158775 630681
rect 159399 630647 159433 630681
rect 160057 630647 160091 630681
rect 160715 630647 160749 630681
rect 161373 630647 161407 630681
rect 162031 630647 162085 630681
rect 158691 630613 158695 630647
rect 158707 630613 162085 630647
rect 158595 628741 158661 630551
rect 158737 630561 158741 630579
rect 158737 630545 158787 630561
rect 158798 630551 158816 630566
rect 158826 630551 158844 630564
rect 159339 630545 159386 630592
rect 159395 630561 159399 630579
rect 159395 630545 159445 630561
rect 159997 630551 160044 630592
rect 159988 630545 160044 630551
rect 160053 630561 160057 630579
rect 160053 630545 160103 630561
rect 160118 630551 160124 630554
rect 160146 630551 160152 630564
rect 160655 630545 160702 630592
rect 160711 630561 160715 630579
rect 160711 630545 160761 630561
rect 161313 630551 161360 630592
rect 161308 630545 161360 630551
rect 161369 630561 161373 630579
rect 161369 630545 161419 630561
rect 161971 630545 162018 630592
rect 158741 630511 159386 630545
rect 159399 630511 160044 630545
rect 160057 630511 160702 630545
rect 160715 630511 161360 630545
rect 161373 630511 162018 630545
rect 158741 630464 158787 630511
rect 158697 630452 158715 630464
rect 158741 630452 158775 630464
rect 158697 628840 158775 630452
rect 158798 629164 158816 630505
rect 158826 629136 158844 630505
rect 159399 630464 159445 630511
rect 159988 630505 160009 630511
rect 160016 630477 160037 630511
rect 160057 630464 160103 630511
rect 159356 630452 159387 630463
rect 159399 630452 159433 630464
rect 160014 630452 160045 630463
rect 160057 630452 160091 630464
rect 141358 625403 141614 625412
rect 141386 625375 141586 625384
rect 135890 625106 136456 625140
rect 135890 624818 135924 625106
rect 136261 625026 136272 625037
rect 135945 624964 136026 625011
rect 136085 624992 136272 625026
rect 136273 624964 136354 625011
rect 135992 624926 136026 624964
rect 136045 624926 136301 624932
rect 136320 624926 136354 624964
rect 136045 624912 136302 624926
rect 136261 624904 136272 624909
rect 136073 624898 136273 624904
rect 136073 624884 136274 624898
rect 136312 624884 136408 624898
rect 136085 624864 136272 624884
rect 136422 624870 136456 625106
rect 136284 624856 136456 624870
rect 136047 624826 136299 624829
rect 136422 624818 136456 624856
rect 135890 624795 136456 624818
rect 135890 624784 135924 624795
rect 136422 624784 136456 624795
rect 135890 624783 136456 624784
rect 135924 624769 136422 624783
rect 135890 624750 136456 624769
rect 136506 624732 137126 625154
rect 140980 624780 140996 624782
rect 140888 624671 141508 624780
rect 141620 624766 142062 624800
rect 141558 624739 142124 624766
rect 140888 624637 144758 624671
rect 140888 624601 141508 624637
rect 141558 624472 141592 624637
rect 141660 624603 141694 624606
rect 141988 624603 142022 624606
rect 142090 624472 142124 624637
rect 128884 621530 128918 624234
rect 129070 621550 137046 621564
rect 137198 621530 137232 624234
rect 158595 623879 158629 628741
rect 158697 628679 158743 628840
rect 159296 628787 159306 630186
rect 159324 628815 159334 630158
rect 159367 628840 159433 630452
rect 160025 628840 160091 630452
rect 160118 629152 160124 630505
rect 160146 629124 160152 630505
rect 160715 630464 160761 630511
rect 161308 630505 161325 630511
rect 161336 630477 161353 630511
rect 161373 630464 161419 630511
rect 160672 630452 160703 630463
rect 160715 630452 160749 630464
rect 161330 630452 161361 630463
rect 161373 630452 161407 630464
rect 159367 628828 159401 628840
rect 160025 628828 160059 628840
rect 159355 628815 159414 628828
rect 159324 628806 159414 628815
rect 159421 628806 159452 628815
rect 159355 628787 159414 628806
rect 159296 628781 159414 628787
rect 158803 628747 159414 628781
rect 159449 628781 159480 628787
rect 160013 628781 160072 628828
rect 160606 628787 160626 630192
rect 160634 628815 160654 630164
rect 160683 628840 160749 630452
rect 161341 628840 161407 630452
rect 161440 629130 161444 630505
rect 161468 629102 161472 630505
rect 161988 630452 162019 630463
rect 162031 630452 162065 630613
rect 160683 628828 160717 628840
rect 161341 628828 161375 628840
rect 160671 628815 160730 628828
rect 160634 628812 160730 628815
rect 160737 628812 160762 628815
rect 160671 628787 160730 628812
rect 160606 628784 160730 628787
rect 160765 628784 160790 628787
rect 160671 628781 160730 628784
rect 161329 628781 161388 628828
rect 161928 628787 161948 630162
rect 161956 628787 161976 630134
rect 161999 628840 162065 630452
rect 162113 630551 162131 630613
rect 162145 630551 162179 630858
rect 163698 630556 163732 630858
rect 163812 630652 163846 630686
rect 164470 630652 164504 630686
rect 165128 630652 165162 630686
rect 165786 630652 165820 630686
rect 166444 630652 166478 630686
rect 167102 630652 167156 630686
rect 163762 630618 163766 630652
rect 163778 630618 167156 630652
rect 161999 628828 162033 628840
rect 161987 628781 162045 628828
rect 159449 628778 160072 628781
rect 159461 628747 160072 628778
rect 160119 628747 160730 628781
rect 160777 628747 161388 628781
rect 161435 628747 162045 628781
rect 159355 628731 159401 628747
rect 160013 628731 160059 628747
rect 160671 628731 160717 628747
rect 161329 628731 161375 628747
rect 161987 628731 162033 628747
rect 162113 628741 162179 630551
rect 163666 628764 163732 630556
rect 163808 630566 163812 630584
rect 163808 630550 163858 630566
rect 164410 630550 164448 630588
rect 164466 630566 164470 630584
rect 164466 630550 164516 630566
rect 165068 630556 165106 630588
rect 165058 630550 165106 630556
rect 165124 630566 165128 630584
rect 165124 630550 165174 630566
rect 165726 630550 165764 630588
rect 165782 630566 165786 630584
rect 165782 630550 165832 630566
rect 166384 630550 166422 630588
rect 166440 630566 166444 630584
rect 166440 630550 166490 630566
rect 167042 630550 167080 630588
rect 163812 630516 164448 630550
rect 164470 630546 165106 630550
rect 164470 630516 165108 630546
rect 163812 630478 163858 630516
rect 164470 630478 164516 630516
rect 165058 630510 165080 630516
rect 165086 630482 165108 630516
rect 165128 630516 165764 630550
rect 165786 630516 166422 630550
rect 166444 630516 167080 630550
rect 165128 630478 165174 630516
rect 165786 630478 165832 630516
rect 166380 630510 166396 630516
rect 166408 630482 166424 630510
rect 166444 630478 166490 630516
rect 163768 630466 163786 630478
rect 163812 630466 163846 630478
rect 164427 630466 164458 630477
rect 164470 630466 164504 630478
rect 165085 630466 165116 630477
rect 165128 630466 165162 630478
rect 165743 630466 165774 630477
rect 165786 630466 165820 630478
rect 166401 630466 166432 630477
rect 166444 630466 166478 630478
rect 163768 628854 163846 630466
rect 161341 628679 161375 628731
rect 158697 628645 162045 628679
rect 158709 623975 158743 624009
rect 159367 623975 159401 624009
rect 160025 623975 160059 624009
rect 160683 623975 160717 624009
rect 161341 623975 161375 628645
rect 161999 623975 162033 624009
rect 158677 623941 162067 623975
rect 140782 621530 140816 623860
rect 149096 621530 149130 623860
rect 158581 622377 158629 623879
rect 158709 623889 158743 623941
rect 159367 623920 159401 623941
rect 160025 623920 160059 623941
rect 160683 623920 160717 623941
rect 161341 623920 161375 623941
rect 161999 623920 162033 623941
rect 159325 623889 159401 623920
rect 159983 623889 160059 623920
rect 160641 623889 160717 623920
rect 161299 623889 161375 623920
rect 158709 623792 158755 623889
rect 159325 623873 159413 623889
rect 159983 623873 160071 623889
rect 160641 623873 160729 623889
rect 161299 623873 161387 623889
rect 161957 623873 162033 623920
rect 162113 623879 162147 628741
rect 163666 626922 163700 628764
rect 163768 628702 163814 628854
rect 164366 628810 164392 629930
rect 164394 628810 164420 629902
rect 164438 628854 164504 630466
rect 165096 628854 165162 630466
rect 164438 628842 164472 628854
rect 165096 628842 165130 628854
rect 164426 628804 164476 628842
rect 164530 628810 164548 628826
rect 165084 628804 165134 628842
rect 165686 628810 165702 629912
rect 165714 628810 165730 629884
rect 165754 628854 165820 630466
rect 166412 628854 166478 630466
rect 166510 629108 166516 630510
rect 166538 629080 166544 630510
rect 167059 630466 167090 630477
rect 167102 630466 167136 630618
rect 165754 628842 165788 628854
rect 166412 628842 166446 628854
rect 165742 628804 165792 628842
rect 166400 628804 166450 628842
rect 166994 628810 167018 629914
rect 167022 628810 167046 629886
rect 167070 628854 167136 630466
rect 167184 630556 167202 630618
rect 167216 630556 167250 630858
rect 167070 628842 167104 628854
rect 167058 628804 167108 628842
rect 163874 628770 164476 628804
rect 164532 628770 165134 628804
rect 165190 628770 165792 628804
rect 165848 628770 166450 628804
rect 166506 628770 167108 628804
rect 164426 628754 164472 628770
rect 165084 628754 165130 628770
rect 165742 628754 165788 628770
rect 166400 628754 166446 628770
rect 167058 628754 167104 628770
rect 167184 628764 167250 630556
rect 164438 628702 164472 628754
rect 163768 628668 167116 628702
rect 164438 626922 164472 628668
rect 166406 626922 166428 627112
rect 167184 626922 167218 628764
rect 163666 626894 167218 626922
rect 163360 626452 163362 626500
rect 163332 626424 163362 626444
rect 163666 623884 163700 626894
rect 164438 626866 164472 626894
rect 166406 626866 166428 626894
rect 163738 626838 167156 626866
rect 163780 623980 163814 624014
rect 164438 623980 164472 626838
rect 166406 626444 166428 626838
rect 165130 624182 165136 625256
rect 165130 624014 165162 624182
rect 165096 623980 165162 624014
rect 165186 623980 165190 624210
rect 165754 623980 165788 624014
rect 166348 623980 166374 624174
rect 166406 624146 166430 625256
rect 166376 624014 166430 624146
rect 166376 623980 166446 624014
rect 167070 623980 167104 624014
rect 163748 623946 167138 623980
rect 158757 623839 159413 623873
rect 159415 623839 160071 623873
rect 160073 623839 160729 623873
rect 160731 623839 161387 623873
rect 161389 623839 162033 623873
rect 159333 623833 159337 623839
rect 159361 623805 159365 623839
rect 159367 623792 159413 623839
rect 160025 623792 160071 623839
rect 160649 623833 160653 623839
rect 160677 623805 160681 623839
rect 160683 623792 160729 623839
rect 161341 623792 161387 623839
rect 161965 623833 161969 623839
rect 161993 623805 161997 623839
rect 158709 623780 158743 623792
rect 159342 623780 159355 623791
rect 159367 623780 159401 623792
rect 160000 623780 160013 623791
rect 160025 623780 160059 623792
rect 160658 623780 160671 623791
rect 160683 623780 160717 623792
rect 161316 623780 161329 623791
rect 161341 623780 161375 623792
rect 161974 623780 161987 623791
rect 161999 623780 162033 623839
rect 158695 622476 158743 623780
rect 159353 622476 159401 623780
rect 160011 622476 160059 623780
rect 125686 621496 152286 621530
rect 128884 621428 128918 621496
rect 128986 621428 129020 621496
rect 129466 621428 129504 621466
rect 130224 621428 130262 621466
rect 130982 621428 131020 621466
rect 131740 621428 131778 621466
rect 132498 621428 132536 621466
rect 133256 621428 133294 621466
rect 134014 621428 134052 621466
rect 134772 621428 134810 621466
rect 135530 621428 135568 621466
rect 136288 621428 136326 621466
rect 137046 621428 137058 621466
rect 128884 621394 129504 621428
rect 129556 621394 130262 621428
rect 130314 621394 131020 621428
rect 131072 621394 131778 621428
rect 131830 621394 132536 621428
rect 132588 621394 133294 621428
rect 133346 621394 134052 621428
rect 134104 621394 134810 621428
rect 134862 621394 135568 621428
rect 135620 621394 136326 621428
rect 136378 621394 137058 621428
rect 127220 616796 127254 621344
rect 128884 620812 128918 621394
rect 128986 620954 129020 621394
rect 137098 621378 137130 621466
rect 137136 621394 137168 621428
rect 129058 621356 129059 621357
rect 137057 621356 137058 621357
rect 137098 621356 137142 621378
rect 129057 621355 129058 621356
rect 137058 621355 137059 621356
rect 129483 621344 129528 621355
rect 130241 621344 130286 621355
rect 130999 621344 131044 621355
rect 131757 621344 131802 621355
rect 132515 621344 132560 621355
rect 133273 621344 133318 621355
rect 134031 621344 134076 621355
rect 134789 621344 134834 621355
rect 135547 621344 135592 621355
rect 136305 621344 136350 621355
rect 129482 620938 129483 620939
rect 129481 620937 129482 620938
rect 129494 620926 129528 621344
rect 129539 620938 129540 620939
rect 130240 620938 130241 620939
rect 129540 620937 129541 620938
rect 130239 620937 130240 620938
rect 130252 620926 130286 621344
rect 130297 620938 130298 620939
rect 130998 620938 130999 620939
rect 130298 620937 130299 620938
rect 130997 620937 130998 620938
rect 131010 620926 131044 621344
rect 131055 620938 131056 620939
rect 131756 620938 131757 620939
rect 131056 620937 131057 620938
rect 131755 620937 131756 620938
rect 131768 620926 131802 621344
rect 131813 620938 131814 620939
rect 132514 620938 132515 620939
rect 131814 620937 131815 620938
rect 132513 620937 132514 620938
rect 132526 620926 132560 621344
rect 132571 620938 132572 620939
rect 133272 620938 133273 620939
rect 132572 620937 132573 620938
rect 133271 620937 133272 620938
rect 133284 620926 133318 621344
rect 133329 620938 133330 620939
rect 134030 620938 134031 620939
rect 133330 620937 133331 620938
rect 134029 620937 134030 620938
rect 134042 620926 134076 621344
rect 134087 620938 134088 620939
rect 134788 620938 134789 620939
rect 134088 620937 134089 620938
rect 134787 620937 134788 620938
rect 134800 620926 134834 621344
rect 134845 620938 134846 620939
rect 135546 620938 135547 620939
rect 134846 620937 134847 620938
rect 135545 620937 135546 620938
rect 135558 620926 135592 621344
rect 135603 620938 135604 620939
rect 136304 620938 136305 620939
rect 135604 620937 135605 620938
rect 136303 620937 136304 620938
rect 136316 620926 136350 621344
rect 137062 620954 137142 621356
rect 136361 620938 136362 620939
rect 137062 620938 137120 620954
rect 136362 620937 136363 620938
rect 137046 620926 137057 620937
rect 129070 620892 137062 620926
rect 129494 620812 129528 620892
rect 130252 620812 130286 620892
rect 131010 620812 131044 620892
rect 131768 620812 131802 620892
rect 132526 620812 132560 620892
rect 133284 620812 133318 620892
rect 134042 620812 134076 620892
rect 134800 620812 134834 620892
rect 135558 620812 135592 620892
rect 136316 620812 136350 620892
rect 137074 620858 137096 620938
rect 137074 620854 137084 620858
rect 137074 620812 137108 620846
rect 137198 620812 137232 621496
rect 140782 621428 140816 621496
rect 140868 621466 140894 621486
rect 139410 621394 140852 621428
rect 128884 620778 137232 620812
rect 132574 620362 132600 620524
rect 132602 620362 132628 620524
rect 132378 619900 133016 620362
rect 133284 620308 133318 620342
rect 133412 620308 133438 620486
rect 133440 620308 133466 620486
rect 133066 620274 133614 620308
rect 133066 619992 133100 620274
rect 133284 620194 133318 620274
rect 133412 620205 133438 620274
rect 133412 620200 133439 620205
rect 133440 620200 133466 620274
rect 133428 620194 133439 620200
rect 133130 620150 133202 620188
rect 133252 620160 133439 620194
rect 133168 620116 133202 620150
rect 133271 620148 133272 620149
rect 133272 620147 133273 620148
rect 133272 620118 133273 620119
rect 133271 620117 133272 620118
rect 133284 620106 133318 620160
rect 133440 620150 133512 620188
rect 133330 620148 133331 620149
rect 133329 620147 133330 620148
rect 133329 620118 133330 620119
rect 133330 620117 133331 620118
rect 133428 620106 133439 620117
rect 133478 620116 133512 620150
rect 133252 620072 133439 620106
rect 133284 619992 133318 620072
rect 133412 619992 133430 620066
rect 133440 619992 133458 620066
rect 133580 619992 133614 620274
rect 133066 619958 133614 619992
rect 132580 619750 132600 619900
rect 132608 619778 132628 619900
rect 133412 619876 133430 619958
rect 133440 619904 133458 619958
rect 133412 619778 133432 619876
rect 133440 619750 133460 619904
rect 129706 619295 130028 619326
rect 132752 619295 133074 619314
rect 128853 616574 137291 619295
rect 140106 616796 140140 621344
rect 140782 620438 140816 621394
rect 140868 621378 140918 621466
rect 141594 621428 141632 621466
rect 142352 621428 142390 621466
rect 143110 621428 143148 621466
rect 143868 621428 143906 621466
rect 144626 621428 144664 621466
rect 145384 621428 145422 621466
rect 146142 621428 146180 621466
rect 146900 621428 146938 621466
rect 147658 621428 147696 621466
rect 148416 621428 148454 621466
rect 148994 621428 149028 621496
rect 149096 621428 149130 621496
rect 140926 621394 141632 621428
rect 141684 621394 142390 621428
rect 142442 621394 143148 621428
rect 143200 621394 143906 621428
rect 143958 621394 144664 621428
rect 144716 621394 145422 621428
rect 145474 621394 146180 621428
rect 146232 621394 146938 621428
rect 146990 621394 147696 621428
rect 147748 621394 148454 621428
rect 148506 621394 149130 621428
rect 140868 621356 140932 621378
rect 140956 621356 140957 621357
rect 148955 621356 148956 621357
rect 140853 621341 140932 621356
rect 140955 621355 140956 621356
rect 148956 621355 148957 621356
rect 141611 621344 141656 621355
rect 142369 621344 142414 621355
rect 143127 621344 143172 621355
rect 143885 621344 143930 621355
rect 144643 621344 144688 621355
rect 145401 621344 145446 621355
rect 146159 621344 146204 621355
rect 146917 621344 146962 621355
rect 147675 621344 147720 621355
rect 148433 621344 148478 621355
rect 140868 621238 140932 621341
rect 140868 621222 140910 621238
rect 141610 621222 141611 621223
rect 141609 621221 141610 621222
rect 141622 621210 141656 621344
rect 141667 621222 141668 621223
rect 142368 621222 142369 621223
rect 141668 621221 141669 621222
rect 142367 621221 142368 621222
rect 142380 621210 142414 621344
rect 142425 621222 142426 621223
rect 143126 621222 143127 621223
rect 142426 621221 142427 621222
rect 143125 621221 143126 621222
rect 143138 621210 143172 621344
rect 143183 621222 143184 621223
rect 143884 621222 143885 621223
rect 143184 621221 143185 621222
rect 143883 621221 143884 621222
rect 143896 621210 143930 621344
rect 143941 621222 143942 621223
rect 144642 621222 144643 621223
rect 143942 621221 143943 621222
rect 144641 621221 144642 621222
rect 144654 621210 144688 621344
rect 144699 621222 144700 621223
rect 145400 621222 145401 621223
rect 144700 621221 144701 621222
rect 145399 621221 145400 621222
rect 145412 621210 145446 621344
rect 145457 621222 145458 621223
rect 146158 621222 146159 621223
rect 145458 621221 145459 621222
rect 146157 621221 146158 621222
rect 146170 621210 146204 621344
rect 146215 621222 146216 621223
rect 146916 621222 146917 621223
rect 146216 621221 146217 621222
rect 146915 621221 146916 621222
rect 146928 621210 146962 621344
rect 146973 621222 146974 621223
rect 147674 621222 147675 621223
rect 146974 621221 146975 621222
rect 147673 621221 147674 621222
rect 147686 621210 147720 621344
rect 147731 621222 147732 621223
rect 148432 621222 148433 621223
rect 147732 621221 147733 621222
rect 148431 621221 148432 621222
rect 148444 621210 148478 621344
rect 148994 621238 149028 621394
rect 148489 621222 148490 621223
rect 148490 621221 148491 621222
rect 148944 621210 148955 621221
rect 140860 621182 140918 621186
rect 140850 621148 140918 621182
rect 140968 621176 148955 621210
rect 141609 621164 141610 621165
rect 141610 621163 141611 621164
rect 140868 620580 140932 621148
rect 140868 620564 140910 620580
rect 141622 620574 141656 621176
rect 141668 621164 141669 621165
rect 142367 621164 142368 621165
rect 141667 621163 141668 621164
rect 142368 621163 142369 621164
rect 141686 620574 142340 620576
rect 141580 620552 142340 620574
rect 142368 620564 142369 620565
rect 142367 620563 142368 620564
rect 142380 620552 142414 621176
rect 142426 621164 142427 621165
rect 143125 621164 143126 621165
rect 142425 621163 142426 621164
rect 143126 621163 143127 621164
rect 142425 620564 142426 620565
rect 143126 620564 143127 620565
rect 142426 620563 142427 620564
rect 143125 620563 143126 620564
rect 143138 620552 143172 621176
rect 143184 621164 143185 621165
rect 143883 621164 143884 621165
rect 143183 621163 143184 621164
rect 143884 621163 143885 621164
rect 143183 620564 143184 620565
rect 143884 620564 143885 620565
rect 143184 620563 143185 620564
rect 143883 620563 143884 620564
rect 143896 620552 143930 621176
rect 144578 621170 144648 621176
rect 143942 621164 143943 621165
rect 144641 621164 144642 621165
rect 143941 621163 143942 621164
rect 144642 621163 144643 621164
rect 144606 621142 144648 621150
rect 144578 620612 144600 620650
rect 144606 620584 144628 620650
rect 143941 620564 143942 620565
rect 144642 620564 144643 620565
rect 143942 620563 143943 620564
rect 144641 620563 144642 620564
rect 144654 620552 144688 621176
rect 144694 621170 144758 621176
rect 144700 621164 144701 621165
rect 145399 621164 145400 621165
rect 144699 621163 144700 621164
rect 145400 621163 145401 621164
rect 144694 621142 144730 621150
rect 144699 620564 144700 620565
rect 145400 620564 145401 620565
rect 144700 620563 144701 620564
rect 145399 620563 145400 620564
rect 145412 620552 145446 621176
rect 145458 621164 145459 621165
rect 146157 621164 146158 621165
rect 145457 621163 145458 621164
rect 146158 621163 146159 621164
rect 145457 620564 145458 620565
rect 146158 620564 146159 620565
rect 145458 620563 145459 620564
rect 146157 620563 146158 620564
rect 146170 620552 146204 621176
rect 146216 621164 146217 621165
rect 146915 621164 146916 621165
rect 146215 621163 146216 621164
rect 146916 621163 146917 621164
rect 146215 620564 146216 620565
rect 146916 620564 146917 620565
rect 146216 620563 146217 620564
rect 146915 620563 146916 620564
rect 146928 620552 146962 621176
rect 146974 621164 146975 621165
rect 147673 621164 147674 621165
rect 146973 621163 146974 621164
rect 147674 621163 147675 621164
rect 147602 621132 147680 621156
rect 147630 621104 147680 621128
rect 146973 620564 146974 620565
rect 147674 620564 147675 620565
rect 146974 620563 146975 620564
rect 147673 620563 147674 620564
rect 147686 620552 147720 621176
rect 147732 621164 147733 621165
rect 148431 621164 148432 621165
rect 147731 621163 147732 621164
rect 148432 621163 148433 621164
rect 147726 621132 147782 621156
rect 147726 621104 147754 621128
rect 147731 620564 147732 620565
rect 148432 620564 148433 620565
rect 147732 620563 147733 620564
rect 148431 620563 148432 620564
rect 148444 620552 148478 621176
rect 148490 621164 148491 621165
rect 148489 621163 148490 621164
rect 148956 621148 149028 621186
rect 148994 620580 149028 621148
rect 148489 620564 148490 620565
rect 148490 620563 148491 620564
rect 148944 620552 148955 620563
rect 140968 620518 148955 620552
rect 141580 620502 142340 620518
rect 140844 620438 140864 620472
rect 141580 620438 141700 620502
rect 142380 620438 142414 620518
rect 143138 620438 143172 620518
rect 143896 620438 143930 620518
rect 144654 620438 144688 620518
rect 145412 620438 145446 620518
rect 146170 620438 146204 620518
rect 146928 620438 146962 620518
rect 147686 620438 147720 620518
rect 148444 620438 148478 620518
rect 149096 620438 149130 621394
rect 140782 620404 149130 620438
rect 144654 619934 144688 619968
rect 144400 619900 144948 619934
rect 144400 619618 144434 619900
rect 144464 619776 144536 619814
rect 144502 619742 144536 619776
rect 144546 619664 144548 619854
rect 144574 619780 144576 619826
rect 144654 619820 144688 619900
rect 144762 619820 144773 619831
rect 144586 619786 144773 619820
rect 144641 619774 144642 619775
rect 144642 619773 144643 619774
rect 144606 619760 144648 619766
rect 144642 619744 144643 619745
rect 144641 619743 144642 619744
rect 144574 619692 144576 619738
rect 144578 619732 144648 619738
rect 144654 619732 144688 619786
rect 144774 619776 144846 619814
rect 144700 619774 144701 619775
rect 144699 619773 144700 619774
rect 144694 619760 144730 619766
rect 144699 619744 144700 619745
rect 144700 619743 144701 619744
rect 144694 619732 144758 619738
rect 144762 619732 144773 619743
rect 144812 619742 144846 619776
rect 144586 619698 144773 619732
rect 144654 619618 144688 619698
rect 144914 619618 144948 619900
rect 144400 619584 144948 619618
rect 144998 619526 145636 619988
rect 144900 618921 145222 619332
rect 140723 616574 149161 618921
rect 150718 616796 150752 621344
rect 151586 616752 151594 621388
rect 151614 616752 151650 621388
rect 158581 615705 158615 622377
rect 158695 622315 158729 622476
rect 159353 622464 159387 622476
rect 160011 622464 160045 622476
rect 158731 622349 158735 622451
rect 158759 622417 158763 622423
rect 159339 622417 159387 622464
rect 159997 622417 160045 622464
rect 158755 622383 158763 622417
rect 158771 622383 159387 622417
rect 159413 622383 159421 622417
rect 159429 622383 160045 622417
rect 158759 622377 158763 622383
rect 159341 622367 159387 622383
rect 159999 622367 160045 622383
rect 159353 622315 159387 622367
rect 160011 622315 160045 622367
rect 160047 622349 160051 622451
rect 160592 622423 160594 623520
rect 160620 622423 160622 623492
rect 160669 622476 160717 623780
rect 161327 622476 161375 623780
rect 160669 622464 160703 622476
rect 161327 622464 161361 622476
rect 160075 622417 160079 622423
rect 160655 622417 160703 622464
rect 161313 622417 161361 622464
rect 160071 622383 160079 622417
rect 160087 622383 160703 622417
rect 160729 622383 160737 622417
rect 160745 622383 161361 622417
rect 160075 622377 160079 622383
rect 160592 622370 160594 622377
rect 160620 622342 160622 622377
rect 160657 622367 160703 622383
rect 161315 622367 161361 622383
rect 160669 622315 160703 622367
rect 161327 622315 161361 622367
rect 161363 622349 161367 622451
rect 161914 622423 161916 623490
rect 161942 622423 161944 623462
rect 161985 622476 162033 623780
rect 161985 622464 162019 622476
rect 161391 622417 161395 622423
rect 161971 622417 162019 622464
rect 161387 622383 161395 622417
rect 161403 622383 162019 622417
rect 161391 622377 161395 622383
rect 161914 622370 161916 622377
rect 161942 622342 161944 622377
rect 161973 622367 162019 622383
rect 161985 622315 162019 622367
rect 162099 622377 162147 623879
rect 163652 622400 163700 623884
rect 163780 623894 163814 623946
rect 164396 623912 164434 623916
rect 163780 623806 163826 623894
rect 164396 623878 164436 623912
rect 163828 623844 164436 623878
rect 164404 623838 164408 623844
rect 164432 623810 164436 623844
rect 164438 623894 164472 623946
rect 164438 623806 164484 623894
rect 165054 623878 165092 623916
rect 164486 623844 165092 623878
rect 165096 623884 165162 623946
rect 165186 623884 165190 623946
rect 165096 623838 165142 623884
rect 165712 623878 165750 623916
rect 165144 623844 165750 623878
rect 165754 623894 165788 623946
rect 166348 623916 166374 623946
rect 166376 623916 166446 623946
rect 166348 623894 166446 623916
rect 167028 623912 167066 623916
rect 163780 623794 163814 623806
rect 164413 623794 164426 623805
rect 164438 623794 164472 623806
rect 165071 623794 165084 623805
rect 165096 623794 165162 623838
rect 163766 622490 163814 623794
rect 158683 622281 162031 622315
rect 162099 615705 162133 622377
rect 163652 615728 163686 622400
rect 163766 622338 163800 622490
rect 163802 622372 163806 622474
rect 164352 622446 164360 623258
rect 164380 622446 164388 623230
rect 164424 622490 164472 623794
rect 165082 622780 165162 623794
rect 164424 622478 164458 622490
rect 165082 622478 165136 622780
rect 165186 622752 165190 623838
rect 165754 623806 165800 623894
rect 166348 623884 166458 623894
rect 166370 623878 166408 623884
rect 165802 623844 166408 623878
rect 166412 623838 166458 623884
rect 167028 623878 167068 623912
rect 166460 623844 167068 623878
rect 167036 623838 167040 623844
rect 165729 623794 165742 623805
rect 165754 623794 165788 623806
rect 165740 622490 165788 623794
rect 166348 622716 166374 623838
rect 166376 623806 166458 623838
rect 167064 623810 167068 623844
rect 166376 622744 166446 623806
rect 167045 623794 167058 623805
rect 167070 623794 167104 623946
rect 167184 623884 167218 626894
rect 167836 625530 175812 625564
rect 168418 624948 169522 624968
rect 166364 622670 166374 622716
rect 166392 622670 166446 622744
rect 166980 622670 166986 623242
rect 167008 622670 167014 623214
rect 166398 622532 166446 622670
rect 165740 622478 165774 622490
rect 163830 622440 163834 622446
rect 164410 622440 164458 622478
rect 165068 622446 165122 622478
rect 165068 622440 165116 622446
rect 163826 622406 163834 622440
rect 163842 622406 164458 622440
rect 164484 622406 164492 622440
rect 164500 622406 165116 622440
rect 163830 622400 163834 622406
rect 164352 622394 164360 622400
rect 164380 622366 164388 622400
rect 164412 622390 164458 622406
rect 165070 622400 165116 622406
rect 165118 622400 165122 622446
rect 165146 622440 165150 622446
rect 165726 622440 165774 622478
rect 166364 622446 166374 622532
rect 166392 622490 166446 622532
rect 166392 622478 166432 622490
rect 166384 622440 166432 622478
rect 165142 622406 165150 622440
rect 165158 622406 165774 622440
rect 165800 622406 165808 622440
rect 165816 622406 166432 622440
rect 165146 622400 165150 622406
rect 165070 622390 165122 622400
rect 165728 622390 165774 622406
rect 164424 622338 164458 622390
rect 165082 622344 165122 622390
rect 165082 622338 165116 622344
rect 165740 622338 165774 622390
rect 166364 622338 166374 622400
rect 166386 622390 166432 622406
rect 166392 622338 166432 622390
rect 166434 622372 166438 622474
rect 166980 622446 166986 622532
rect 167008 622446 167014 622532
rect 167056 622490 167104 623794
rect 167056 622478 167090 622490
rect 166462 622440 166466 622446
rect 167042 622440 167090 622478
rect 166458 622406 166466 622440
rect 166474 622406 167090 622440
rect 166462 622400 166466 622406
rect 166980 622388 166986 622400
rect 167008 622366 167014 622400
rect 167044 622390 167090 622406
rect 167056 622338 167090 622390
rect 167170 622400 167218 623884
rect 167614 623870 170925 624011
rect 167497 623839 170925 623870
rect 167614 623836 170925 623839
rect 167417 623458 167440 623820
rect 167463 623805 170925 623836
rect 167445 623458 167468 623792
rect 167614 622818 170925 623805
rect 172408 623946 175943 623980
rect 172408 623590 172442 623946
rect 173152 623878 173190 623916
rect 173810 623878 173848 623916
rect 174468 623878 174506 623916
rect 175126 623878 175164 623916
rect 175784 623878 175822 623916
rect 172584 623844 173190 623878
rect 173242 623844 173848 623878
rect 173900 623844 174506 623878
rect 174558 623844 175164 623878
rect 175216 623844 175822 623878
rect 175862 623834 175880 623844
rect 172511 623794 172556 623805
rect 173169 623794 173214 623805
rect 173827 623794 173872 623805
rect 174485 623794 174530 623805
rect 175143 623794 175188 623805
rect 172522 623590 172556 623794
rect 172567 623602 172568 623603
rect 173168 623602 173169 623603
rect 172568 623601 172569 623602
rect 173167 623601 173168 623602
rect 173180 623590 173214 623794
rect 173225 623602 173226 623603
rect 173826 623602 173827 623603
rect 173226 623601 173227 623602
rect 173825 623601 173826 623602
rect 173838 623590 173872 623794
rect 173883 623602 173884 623603
rect 174484 623602 174485 623603
rect 173884 623601 173885 623602
rect 174483 623601 174484 623602
rect 174496 623590 174530 623794
rect 174541 623602 174542 623603
rect 175142 623602 175143 623603
rect 174542 623601 174543 623602
rect 175141 623601 175142 623602
rect 175154 623590 175188 623794
rect 175778 623682 175796 623834
rect 175856 623832 175880 623834
rect 175828 623806 175846 623810
rect 175856 623806 175884 623832
rect 175806 623805 175884 623806
rect 175801 623794 175884 623805
rect 175806 623654 175884 623794
rect 175812 623618 175884 623654
rect 175812 623606 175880 623618
rect 175199 623602 175200 623603
rect 175800 623602 175801 623603
rect 175200 623601 175201 623602
rect 175799 623601 175800 623602
rect 175812 623590 175858 623606
rect 175862 623602 175880 623606
rect 175892 623602 175896 623946
rect 175926 623618 175943 623946
rect 172408 623587 175858 623590
rect 172408 623578 175852 623587
rect 172408 623568 175846 623578
rect 175926 623575 175930 623618
rect 172408 623566 175852 623568
rect 172408 623556 175858 623566
rect 172408 622932 172442 623556
rect 172522 622932 172556 623556
rect 172568 623544 172569 623545
rect 173167 623544 173168 623545
rect 172567 623543 172568 623544
rect 173168 623543 173169 623544
rect 172567 622944 172568 622945
rect 173168 622944 173169 622945
rect 172568 622943 172569 622944
rect 173167 622943 173168 622944
rect 173180 622932 173214 623556
rect 173226 623544 173227 623545
rect 173825 623544 173826 623545
rect 173225 623543 173226 623544
rect 173826 623543 173827 623544
rect 173225 622944 173226 622945
rect 173826 622944 173827 622945
rect 173226 622943 173227 622944
rect 173825 622943 173826 622944
rect 173838 622932 173872 623556
rect 173884 623544 173885 623545
rect 174483 623544 174484 623545
rect 173883 623543 173884 623544
rect 174484 623543 174485 623544
rect 173883 622944 173884 622945
rect 174484 622944 174485 622945
rect 173884 622943 173885 622944
rect 174483 622943 174484 622944
rect 174496 622932 174530 623556
rect 174542 623544 174543 623545
rect 175141 623544 175142 623545
rect 174541 623543 174542 623544
rect 175142 623543 175143 623544
rect 174541 622944 174542 622945
rect 175142 622944 175143 622945
rect 174542 622943 174543 622944
rect 175141 622943 175142 622944
rect 175154 622932 175188 623556
rect 175200 623544 175201 623545
rect 175799 623544 175800 623545
rect 175199 623543 175200 623544
rect 175800 623543 175801 623544
rect 175812 623540 175858 623556
rect 175862 623540 175880 623544
rect 175812 623528 175880 623540
rect 175812 623478 175884 623528
rect 175199 622944 175200 622945
rect 175800 622944 175801 622945
rect 175200 622943 175201 622944
rect 175799 622943 175800 622944
rect 175812 622932 175858 623478
rect 175862 622960 175884 623478
rect 175862 622944 175880 622960
rect 175892 622944 175896 623544
rect 175926 622960 175943 623575
rect 172408 622929 175858 622932
rect 172408 622898 175846 622929
rect 175926 622910 175930 622960
rect 172408 622818 172442 622898
rect 172522 622818 172556 622898
rect 173180 622818 173214 622898
rect 173838 622818 173872 622898
rect 174496 622818 174530 622898
rect 175154 622818 175188 622898
rect 175812 622818 175846 622898
rect 167614 622784 175858 622818
rect 175926 622784 175936 622852
rect 175964 622818 175998 624034
rect 197393 623583 197427 629947
rect 199475 626148 199521 628208
rect 199524 626148 199549 628208
rect 197507 623679 197541 623713
rect 198165 623679 198199 623713
rect 198823 623679 198857 623713
rect 199475 623679 199521 624960
rect 199524 623679 199549 624960
rect 200139 623679 200173 629848
rect 200754 628178 200770 628514
rect 200911 623975 200945 629947
rect 203236 624011 203270 629862
rect 205379 624016 206052 627223
rect 211884 626508 213348 626514
rect 211440 625723 212220 625734
rect 211478 625685 212182 625696
rect 211946 625132 213298 625148
rect 208964 625065 209022 625078
rect 212700 625065 212792 625078
rect 208998 625031 209022 625044
rect 212700 625031 212758 625044
rect 202428 623975 203835 624011
rect 205379 623980 208906 624016
rect 200247 623941 203835 623975
rect 200247 623679 200281 623941
rect 200376 623873 200843 623920
rect 200423 623839 200843 623873
rect 200785 623792 200843 623839
rect 200350 623780 200406 623791
rect 200361 623679 200406 623780
rect 200797 623713 200842 623792
rect 200797 623679 200851 623713
rect 200911 623679 200945 623941
rect 201648 623848 201661 623879
rect 201615 623833 201661 623848
rect 202385 623848 202408 623879
rect 202428 623848 203835 623941
rect 202385 623833 203835 623848
rect 202428 623720 203835 623833
rect 197457 623645 197461 623679
rect 197473 623645 200945 623679
rect 167614 622748 170925 622784
rect 163754 622304 167102 622338
rect 164424 615818 164458 622304
rect 166364 621936 166374 622304
rect 166392 621936 166430 622304
rect 165806 621430 166398 621444
rect 166432 621430 166586 621444
rect 165840 621396 166398 621410
rect 166432 621396 166586 621410
rect 166364 617976 166374 620748
rect 166392 617976 166430 620748
rect 165124 617050 165148 617510
rect 165130 616108 165148 617050
rect 165082 615818 165122 615830
rect 165076 615806 165122 615818
rect 166364 615778 166374 616072
rect 166392 615830 166430 616072
rect 166524 616016 166526 617530
rect 166392 615818 166432 615830
rect 166392 615806 166438 615818
rect 167170 615728 167204 622400
rect 167413 622328 167414 622414
rect 167451 622290 167452 622452
rect 167620 622410 168042 622748
rect 168109 621265 168143 621299
rect 168767 621265 168801 621299
rect 169425 621265 169459 621299
rect 170083 621265 170117 621299
rect 170741 621265 170775 621299
rect 170855 621265 170889 622748
rect 170890 622368 170925 622622
rect 171144 621906 171179 622368
rect 171600 622196 171702 622208
rect 172408 621301 172442 622784
rect 172484 622556 172498 622642
rect 172522 622518 172536 622680
rect 197361 621773 197427 623583
rect 197503 623593 197507 623611
rect 197503 623577 197553 623593
rect 197564 623583 197582 623598
rect 197592 623583 197610 623596
rect 198105 623577 198152 623624
rect 198161 623593 198165 623611
rect 198161 623577 198211 623593
rect 198763 623583 198810 623624
rect 198754 623577 198810 623583
rect 198819 623593 198823 623611
rect 198819 623577 198869 623593
rect 198884 623583 198890 623586
rect 198912 623583 198918 623596
rect 199421 623577 199468 623624
rect 199475 623593 199521 623645
rect 199524 623593 199549 623645
rect 199475 623583 199549 623593
rect 199477 623577 199527 623583
rect 200079 623577 200126 623624
rect 200139 623611 200173 623645
rect 200135 623593 200173 623611
rect 200135 623577 200185 623593
rect 200247 623577 200281 623645
rect 200361 623642 200406 623645
rect 200797 623642 200842 623645
rect 200361 623624 200395 623642
rect 200361 623577 200408 623624
rect 200737 623577 200784 623624
rect 197507 623543 198152 623577
rect 198165 623543 198810 623577
rect 198823 623543 199468 623577
rect 199481 623543 200126 623577
rect 200139 623543 200784 623577
rect 197507 623496 197553 623543
rect 197463 623484 197481 623496
rect 197507 623484 197541 623496
rect 197463 621860 197541 623484
rect 197564 622196 197582 623537
rect 197592 622168 197610 623537
rect 198165 623496 198211 623543
rect 198754 623537 198775 623543
rect 198782 623509 198803 623543
rect 198823 623496 198869 623543
rect 199481 623537 199527 623543
rect 198122 623484 198153 623495
rect 198165 623484 198199 623496
rect 198780 623484 198811 623495
rect 198823 623484 198857 623496
rect 198062 621860 198072 623218
rect 198090 621860 198100 623190
rect 198133 621860 198199 623484
rect 198791 621860 198857 623484
rect 198884 622184 198890 623537
rect 198912 622156 198918 623537
rect 199475 623496 199549 623537
rect 199468 623495 199521 623496
rect 199438 623484 199521 623495
rect 199344 621860 199392 623252
rect 199449 623196 199521 623484
rect 199524 623196 199549 623496
rect 200139 623496 200185 623543
rect 200096 623484 200127 623495
rect 200139 623484 200173 623496
rect 199400 621860 199420 623196
rect 199449 621860 199515 623196
rect 200107 621872 200173 623484
rect 200107 621860 200141 621872
rect 197463 621856 199828 621860
rect 197463 621846 197509 621856
rect 197522 621846 199828 621856
rect 197463 621822 199828 621846
rect 197361 621370 197395 621773
rect 197463 621711 197509 621822
rect 197522 621813 199828 621822
rect 200095 621813 200154 621860
rect 200247 621813 200281 623543
rect 200361 621860 200395 623543
rect 200797 623495 200831 623642
rect 200754 623484 200831 623495
rect 200765 621872 200831 623484
rect 200765 621860 200810 621872
rect 200361 621813 200408 621860
rect 200753 621813 200812 621860
rect 197569 621779 198180 621813
rect 198215 621810 198838 621813
rect 198227 621779 198838 621810
rect 198885 621779 199496 621813
rect 199543 621779 200154 621813
rect 200185 621779 200812 621813
rect 198121 621763 198167 621779
rect 198779 621763 198825 621779
rect 199437 621763 199489 621779
rect 200095 621763 200141 621779
rect 199468 621711 199489 621763
rect 200107 621711 200141 621763
rect 200247 621711 200281 621779
rect 200361 621711 200395 621779
rect 200753 621763 200799 621779
rect 200765 621711 200799 621763
rect 200879 621711 200945 623645
rect 202396 623684 203835 623720
rect 205318 623946 208906 623980
rect 203894 623684 203928 623718
rect 204552 623684 204586 623718
rect 205210 623684 205244 623718
rect 205318 623684 205352 623946
rect 205379 623684 208906 623946
rect 202396 623669 208906 623684
rect 209003 623941 212555 623975
rect 209003 623783 209037 623941
rect 209747 623873 209794 623920
rect 210405 623873 210452 623920
rect 211063 623873 211110 623920
rect 211721 623873 211768 623920
rect 212379 623873 212426 623920
rect 209179 623839 209794 623873
rect 209837 623839 210452 623873
rect 210495 623839 211110 623873
rect 211153 623839 211768 623873
rect 211811 623839 212426 623873
rect 212324 623833 212391 623839
rect 212324 623805 212419 623826
rect 209163 623792 209763 623795
rect 209821 623792 210421 623795
rect 210479 623792 211079 623795
rect 211137 623792 211737 623795
rect 211795 623792 212395 623795
rect 212521 623783 212555 623941
rect 216294 623884 216310 623904
rect 209003 623749 212555 623783
rect 209003 623669 209037 623749
rect 209117 623669 209151 623749
rect 209775 623669 209809 623749
rect 210433 623669 210467 623749
rect 211091 623669 211125 623749
rect 211749 623669 211783 623749
rect 212407 623669 212441 623749
rect 212521 623669 212555 623749
rect 202396 623650 213685 623669
rect 202396 623620 203835 623650
rect 202396 623578 203872 623620
rect 203882 623598 203902 623644
rect 203882 623588 203940 623598
rect 203890 623582 203940 623588
rect 204492 623582 204530 623620
rect 204548 623598 204552 623616
rect 204548 623582 204598 623598
rect 205150 623582 205188 623620
rect 205206 623598 205210 623616
rect 205248 623598 205250 623650
rect 205206 623582 205256 623598
rect 205304 623588 205306 623614
rect 205318 623582 205352 623650
rect 205379 623635 213685 623650
rect 205379 623599 208906 623635
rect 205432 623582 205470 623599
rect 205808 623582 205846 623599
rect 202396 623548 203874 623578
rect 202396 623542 203846 623548
rect 200976 622134 200982 623486
rect 202396 622998 203835 623542
rect 203852 623514 203874 623548
rect 203894 623548 204530 623582
rect 204552 623548 205188 623582
rect 205210 623548 205846 623582
rect 203852 623509 203866 623514
rect 203894 623510 203940 623548
rect 204552 623510 204598 623548
rect 205210 623542 205256 623548
rect 205318 623542 205352 623548
rect 205210 623510 205282 623542
rect 203851 623498 203882 623509
rect 203894 623498 203928 623510
rect 204509 623498 204540 623509
rect 204552 623498 204586 623510
rect 205167 623498 205198 623509
rect 205210 623498 205244 623510
rect 202378 622140 203835 622998
rect 203852 622176 203928 623498
rect 197463 621677 200945 621711
rect 202396 621836 203835 622140
rect 203856 621886 203928 622176
rect 204520 622118 204586 623498
rect 205178 622118 205244 623498
rect 205248 622366 205282 623510
rect 205304 622366 205352 623542
rect 205318 622228 205352 622366
rect 205248 622140 205282 622228
rect 205248 622118 205250 622140
rect 204520 621886 204597 622118
rect 205178 621886 205255 622118
rect 205304 622084 205352 622228
rect 203856 621874 203896 621886
rect 204520 621874 204554 621886
rect 205178 621874 205250 621886
rect 205304 621874 205306 622084
rect 205318 621874 205352 622084
rect 205432 622118 205466 623548
rect 205868 623509 205902 623599
rect 205825 623498 205902 623509
rect 205432 622116 205477 622118
rect 205836 622116 205902 623498
rect 205950 622116 206016 623599
rect 206052 623230 206068 623232
rect 206046 622366 206068 623230
rect 206090 623134 206124 623599
rect 206090 623052 206190 623134
rect 206046 622126 206068 622228
rect 206090 622116 206124 623052
rect 206400 622440 206862 623078
rect 206454 622356 206804 622390
rect 206182 622228 206216 622240
rect 206182 622200 206216 622212
rect 206454 622116 206488 622356
rect 206770 622328 206804 622356
rect 206646 622288 206684 622326
rect 206736 622294 206804 622328
rect 206612 622254 206684 622288
rect 206664 622234 206724 622244
rect 206770 622234 206816 622294
rect 206664 622228 206742 622234
rect 206770 622228 206874 622234
rect 206664 622215 206696 622216
rect 206557 622204 206602 622215
rect 206645 622206 206696 622215
rect 206770 622206 206816 622228
rect 206645 622204 206742 622206
rect 206568 622116 206602 622204
rect 206656 622200 206742 622204
rect 206770 622200 206874 622206
rect 206656 622116 206690 622200
rect 206770 622150 206816 622200
rect 206748 622116 206816 622150
rect 207406 622116 207440 622150
rect 208064 622116 208098 622150
rect 208722 622116 208756 622150
rect 208836 622116 208870 623599
rect 209003 622972 209037 623635
rect 209704 623376 209718 623514
rect 209704 623116 209712 623376
rect 209732 623348 209746 623486
rect 209732 623116 209740 623348
rect 209117 622972 209130 622974
rect 208878 622202 208904 622940
rect 209003 622550 209640 622972
rect 209752 622964 209775 622992
rect 209752 622958 209828 622964
rect 209854 622958 209860 623018
rect 209882 622958 209888 623018
rect 209690 622924 210256 622958
rect 209690 622602 209724 622924
rect 209758 622808 209828 622924
rect 209854 622878 209860 622924
rect 209752 622782 209828 622808
rect 209752 622744 209843 622782
rect 209845 622776 209860 622878
rect 209882 622850 209888 622924
rect 209873 622844 209888 622850
rect 210061 622844 210072 622855
rect 209873 622810 210072 622844
rect 209873 622804 209888 622810
rect 210073 622782 210154 622829
rect 209845 622744 209860 622750
rect 210120 622744 210154 622782
rect 209752 622718 209828 622744
rect 209758 622636 209828 622718
rect 209752 622602 209828 622636
rect 209844 622602 209860 622744
rect 209873 622716 209888 622722
rect 210061 622716 210072 622727
rect 209872 622682 210072 622716
rect 209872 622602 209888 622682
rect 210222 622602 210256 622924
rect 209690 622568 210256 622602
rect 209003 622152 209037 622550
rect 209083 622202 209096 622550
rect 209117 622168 209130 622550
rect 209758 622508 209828 622568
rect 209704 622220 209730 622420
rect 209732 622192 209758 622448
rect 209844 622156 209860 622568
rect 209872 622184 209888 622568
rect 212521 622152 212555 623635
rect 208967 622116 212591 622152
rect 205432 622082 212591 622116
rect 205432 622054 205477 622082
rect 205404 622020 205477 622054
rect 205432 621874 205500 622020
rect 205836 622002 205902 622082
rect 205950 622002 206016 622082
rect 206090 622002 206124 622082
rect 206454 622002 206488 622082
rect 206568 622012 206602 622082
rect 206614 622012 206644 622014
rect 206656 622012 206690 622082
rect 206578 622006 206680 622012
rect 206574 622002 206684 622006
rect 206748 622002 206816 622082
rect 207406 622002 207440 622082
rect 208064 622002 208098 622082
rect 208722 622002 208756 622082
rect 208836 622002 208870 622082
rect 205502 621940 205574 621978
rect 205624 621968 208870 622002
rect 203850 621836 203900 621874
rect 204376 621836 204558 621874
rect 204576 621842 205218 621874
rect 204576 621836 205216 621842
rect 205234 621836 205500 621874
rect 205540 621836 205574 621940
rect 205836 621886 205902 621968
rect 205836 621870 205881 621886
rect 205836 621836 205874 621870
rect 202396 621802 203900 621836
rect 203956 621802 204558 621836
rect 204614 621802 205216 621836
rect 205260 621802 205874 621836
rect 202396 621734 203835 621802
rect 203850 621786 203896 621802
rect 204508 621786 204554 621802
rect 205166 621796 205212 621802
rect 205260 621796 205274 621802
rect 205166 621786 205218 621796
rect 205178 621740 205218 621786
rect 205178 621734 205212 621740
rect 205318 621734 205352 621802
rect 205432 621734 205500 621802
rect 205540 621738 205574 621802
rect 205836 621738 205870 621802
rect 205540 621734 205612 621738
rect 205836 621734 205881 621738
rect 205950 621734 206016 621968
rect 206077 621956 206078 621957
rect 206078 621955 206079 621956
rect 202396 621700 206016 621734
rect 206090 621882 206124 621968
rect 206136 621956 206137 621957
rect 206135 621955 206136 621956
rect 206090 621810 206135 621882
rect 206454 621876 206488 621968
rect 206596 621956 206684 621968
rect 206735 621956 206736 621957
rect 206612 621944 206684 621956
rect 206736 621955 206737 621956
rect 206748 621938 206816 621968
rect 207393 621956 207394 621957
rect 207394 621955 207395 621956
rect 206748 621876 206804 621938
rect 206454 621842 206804 621876
rect 206090 621724 206162 621810
rect 199468 621370 199489 621677
rect 196176 621336 199632 621370
rect 172372 621265 175996 621301
rect 167655 621231 175996 621265
rect 167655 617747 167689 621231
rect 168109 621230 168143 621231
rect 168109 621157 168149 621230
rect 168168 621157 168177 621202
rect 168109 621151 168143 621157
rect 168767 621151 168801 621231
rect 169425 621151 169459 621231
rect 170083 621151 170117 621231
rect 170741 621151 170775 621231
rect 170855 621151 170889 621231
rect 167710 621089 167791 621136
rect 167850 621117 170889 621151
rect 168109 621111 168143 621117
rect 168096 621105 168097 621106
rect 168097 621104 168098 621105
rect 167757 620521 167791 621089
rect 168109 621046 168149 621111
rect 168155 621105 168156 621106
rect 168154 621104 168155 621105
rect 168168 621074 168177 621111
rect 168754 621105 168755 621106
rect 168755 621104 168756 621105
rect 168097 620505 168098 620506
rect 168096 620504 168097 620505
rect 168109 620493 168143 621046
rect 168154 620505 168155 620506
rect 168755 620505 168756 620506
rect 168155 620504 168156 620505
rect 168754 620504 168755 620505
rect 168767 620493 168801 621117
rect 168813 621105 168814 621106
rect 169412 621105 169413 621106
rect 168812 621104 168813 621105
rect 169413 621104 169414 621105
rect 168812 620505 168813 620506
rect 169413 620505 169414 620506
rect 168813 620504 168814 620505
rect 169412 620504 169413 620505
rect 169425 620493 169459 621117
rect 169471 621105 169472 621106
rect 170070 621105 170071 621106
rect 169470 621104 169471 621105
rect 170071 621104 170072 621105
rect 169470 620505 169471 620506
rect 170071 620505 170072 620506
rect 169471 620504 169472 620505
rect 170070 620504 170071 620505
rect 170083 620493 170117 621117
rect 170129 621105 170130 621106
rect 170728 621105 170729 621106
rect 170128 621104 170129 621105
rect 170729 621104 170730 621105
rect 170128 620505 170129 620506
rect 170729 620505 170730 620506
rect 170129 620504 170130 620505
rect 170728 620504 170729 620505
rect 170741 620493 170775 621117
rect 170855 620493 170889 621117
rect 172372 620493 176014 621231
rect 189214 621206 189218 621211
rect 189144 621178 189190 621183
rect 189144 621171 189212 621178
rect 189150 621168 189212 621171
rect 167710 620431 167791 620478
rect 167850 620459 176014 620493
rect 168096 620447 168097 620448
rect 168097 620446 168098 620447
rect 167757 619863 167791 620431
rect 168097 619847 168098 619848
rect 168096 619846 168097 619847
rect 168109 619835 168143 620459
rect 168155 620447 168156 620448
rect 168754 620447 168755 620448
rect 168154 620446 168155 620447
rect 168755 620446 168756 620447
rect 168767 619850 168801 620459
rect 168813 620447 168814 620448
rect 169412 620447 169413 620448
rect 168812 620446 168813 620447
rect 169413 620446 169414 620447
rect 168992 619850 169204 619982
rect 168154 619847 168155 619848
rect 168155 619846 168156 619847
rect 168682 619835 169204 619850
rect 169413 619847 169414 619848
rect 169412 619846 169413 619847
rect 169425 619835 169459 620459
rect 169471 620447 169472 620448
rect 170070 620447 170071 620448
rect 169470 620446 169471 620447
rect 170071 620446 170072 620447
rect 169470 619847 169471 619848
rect 170071 619847 170072 619848
rect 169471 619846 169472 619847
rect 170070 619846 170071 619847
rect 170083 619835 170117 620459
rect 170129 620447 170130 620448
rect 170728 620447 170729 620448
rect 170128 620446 170129 620447
rect 170729 620446 170730 620447
rect 170128 619847 170129 619848
rect 170729 619847 170730 619848
rect 170129 619846 170130 619847
rect 170728 619846 170729 619847
rect 170741 619835 170775 620459
rect 170855 619835 170889 620459
rect 171566 620416 171956 620450
rect 170920 619934 171176 619940
rect 171566 619918 171600 620416
rect 171780 620348 171827 620395
rect 171742 620314 171827 620348
rect 171669 620255 171714 620266
rect 171797 620255 171842 620266
rect 171680 620079 171714 620255
rect 171808 620079 171842 620255
rect 171780 620020 171827 620067
rect 171742 619986 171827 620020
rect 171922 619918 171956 620416
rect 172076 619934 172332 619952
rect 170948 619906 171148 619912
rect 171566 619884 171956 619918
rect 172104 619906 172304 619924
rect 167710 619773 167791 619820
rect 167850 619801 170889 619835
rect 168096 619789 168097 619790
rect 168097 619788 168098 619789
rect 167757 619205 167791 619773
rect 168097 619189 168098 619190
rect 168096 619188 168097 619189
rect 168109 619177 168143 619801
rect 168155 619789 168156 619790
rect 168154 619788 168155 619789
rect 168682 619780 169204 619801
rect 169412 619789 169413 619790
rect 169413 619788 169414 619789
rect 168154 619189 168155 619190
rect 168755 619189 168756 619190
rect 168155 619188 168156 619189
rect 168754 619188 168755 619189
rect 168767 619177 168801 619780
rect 168992 619534 169204 619780
rect 168812 619189 168813 619190
rect 169413 619189 169414 619190
rect 168813 619188 168814 619189
rect 169412 619188 169413 619189
rect 169425 619177 169459 619801
rect 169471 619789 169472 619790
rect 170070 619789 170071 619790
rect 169470 619788 169471 619789
rect 170071 619788 170072 619789
rect 169470 619189 169471 619190
rect 170071 619189 170072 619190
rect 169471 619188 169472 619189
rect 170070 619188 170071 619189
rect 170083 619177 170117 619801
rect 170129 619789 170130 619790
rect 170728 619789 170729 619790
rect 170128 619788 170129 619789
rect 170729 619788 170730 619789
rect 170128 619189 170129 619190
rect 170729 619189 170730 619190
rect 170129 619188 170130 619189
rect 170728 619188 170729 619189
rect 170741 619177 170775 619801
rect 170855 619177 170889 619801
rect 171148 619720 171408 619740
rect 171148 619692 171408 619712
rect 171552 619214 171974 619834
rect 172104 619724 172304 619740
rect 172076 619696 172332 619712
rect 172372 619177 176014 620459
rect 186992 619757 187428 619780
rect 187026 619723 187394 619746
rect 187899 619658 187933 621125
rect 189158 620986 189212 621168
rect 189158 620698 189190 620986
rect 189150 620695 189190 620698
rect 189144 620683 189190 620695
rect 189214 620958 189240 621206
rect 190460 621180 190506 621183
rect 190442 621171 190506 621180
rect 196888 621182 196892 621187
rect 190442 621168 190500 621171
rect 190442 620994 190458 621168
rect 196888 620996 196916 621182
rect 189214 620655 189218 620958
rect 190460 620695 190500 620698
rect 190460 620683 190506 620695
rect 189212 620602 189780 620636
rect 191984 620336 192208 620356
rect 194176 620340 194396 620360
rect 192004 620184 192005 620336
rect 192188 620184 192208 620336
rect 194196 620184 194197 620340
rect 194376 620184 194396 620340
rect 196888 620144 196892 620996
rect 167710 619115 167791 619162
rect 167850 619143 176014 619177
rect 168096 619131 168097 619132
rect 168097 619130 168098 619131
rect 167757 618547 167791 619115
rect 168097 618531 168098 618532
rect 168096 618530 168097 618531
rect 168109 618519 168143 619143
rect 168155 619131 168156 619132
rect 168754 619131 168755 619132
rect 168154 619130 168155 619131
rect 168755 619130 168756 619131
rect 168154 618531 168155 618532
rect 168755 618531 168756 618532
rect 168155 618530 168156 618531
rect 168754 618530 168755 618531
rect 168767 618519 168801 619143
rect 168813 619131 168814 619132
rect 169412 619131 169413 619132
rect 168812 619130 168813 619131
rect 169413 619130 169414 619131
rect 168812 618531 168813 618532
rect 169413 618531 169414 618532
rect 168813 618530 168814 618531
rect 169412 618530 169413 618531
rect 169425 618519 169459 619143
rect 169471 619131 169472 619132
rect 170070 619131 170071 619132
rect 169470 619130 169471 619131
rect 170071 619130 170072 619131
rect 169470 618531 169471 618532
rect 170071 618531 170072 618532
rect 169471 618530 169472 618531
rect 170070 618530 170071 618531
rect 170083 618519 170117 619143
rect 170129 619131 170130 619132
rect 170728 619131 170729 619132
rect 170128 619130 170129 619131
rect 170729 619130 170730 619131
rect 170128 618531 170129 618532
rect 170729 618531 170730 618532
rect 170129 618530 170130 618531
rect 170728 618530 170729 618531
rect 170741 618519 170775 619143
rect 170855 618519 170889 619143
rect 172116 619072 172158 619078
rect 172296 619072 172324 619078
rect 172088 619044 172158 619050
rect 172296 619044 172352 619050
rect 167710 618457 167791 618504
rect 167850 618485 170889 618519
rect 168096 618473 168097 618474
rect 168097 618472 168098 618473
rect 167757 617889 167791 618457
rect 168097 617873 168098 617874
rect 168096 617872 168097 617873
rect 168109 617861 168143 618485
rect 168155 618473 168156 618474
rect 168754 618473 168755 618474
rect 168154 618472 168155 618473
rect 168755 618472 168756 618473
rect 168154 617873 168155 617874
rect 168755 617873 168756 617874
rect 168155 617872 168156 617873
rect 168754 617872 168755 617873
rect 168767 617861 168801 618485
rect 168813 618473 168814 618474
rect 169412 618473 169413 618474
rect 168812 618472 168813 618473
rect 169413 618472 169414 618473
rect 168812 617873 168813 617874
rect 169413 617873 169414 617874
rect 168813 617872 168814 617873
rect 169412 617872 169413 617873
rect 169425 617861 169459 618485
rect 169471 618473 169472 618474
rect 170070 618473 170071 618474
rect 169470 618472 169471 618473
rect 170071 618472 170072 618473
rect 169470 617873 169471 617874
rect 170071 617873 170072 617874
rect 169471 617872 169472 617873
rect 170070 617872 170071 617873
rect 170083 617861 170117 618485
rect 170129 618473 170130 618474
rect 170728 618473 170729 618474
rect 170128 618472 170129 618473
rect 170729 618472 170730 618473
rect 170128 617873 170129 617874
rect 170729 617873 170730 617874
rect 170129 617872 170130 617873
rect 170728 617872 170729 617873
rect 170741 617861 170775 618485
rect 170855 617861 170889 618485
rect 171554 618479 171810 618498
rect 171582 618451 171782 618470
rect 167850 617827 170889 617861
rect 168109 617747 168143 617827
rect 168767 617747 168801 617827
rect 169425 617747 169459 617827
rect 170083 617747 170117 617827
rect 170741 617747 170775 617827
rect 170855 617747 170889 617827
rect 172372 617747 176014 619143
rect 187356 619624 189496 619658
rect 187356 619133 187390 619624
rect 187797 619556 187831 619624
rect 187899 619556 187933 619624
rect 187532 619522 187933 619556
rect 187749 619475 187750 619476
rect 187750 619474 187751 619475
rect 187459 619463 187504 619474
rect 187470 619133 187504 619463
rect 187797 619161 187831 619522
rect 187515 619145 187516 619146
rect 187516 619144 187517 619145
rect 187738 619133 187749 619144
rect 187356 619099 187749 619133
rect 180124 618435 180380 618444
rect 180152 618407 180352 618416
rect 187356 618326 187390 619099
rect 187470 618487 187504 619099
rect 187516 619087 187517 619088
rect 187515 619086 187516 619087
rect 187750 619071 187831 619118
rect 187515 618487 187516 618488
rect 187516 618486 187517 618487
rect 187534 618486 187536 618509
rect 187797 618503 187831 619071
rect 187534 618475 187564 618481
rect 187738 618475 187749 618486
rect 187432 618462 187750 618475
rect 187432 618449 187754 618462
rect 187482 618441 187754 618449
rect 187492 618435 187750 618441
rect 187516 618429 187750 618435
rect 187520 618428 187572 618429
rect 187899 618428 187933 619522
rect 190674 619266 190698 619476
rect 188828 618750 188852 618758
rect 188828 618498 188854 618750
rect 188828 618486 188852 618498
rect 187516 618407 187933 618428
rect 187532 618394 187933 618407
rect 187797 618326 187831 618394
rect 187899 618326 187933 618394
rect 167655 617713 175996 617747
rect 170855 617398 170889 617713
rect 172372 617677 175996 617713
rect 167614 617362 170925 617398
rect 172408 617362 172442 617677
rect 174526 617412 174530 617574
rect 174564 617450 174568 617536
rect 172522 617362 172556 617396
rect 173180 617362 173214 617396
rect 173838 617362 173872 617396
rect 174496 617362 174530 617396
rect 175154 617362 175188 617396
rect 175812 617362 175846 617396
rect 167614 617328 175858 617362
rect 175926 617328 175936 617396
rect 167614 616358 170925 617328
rect 172408 617248 172442 617328
rect 172522 617248 172556 617328
rect 173180 617248 173214 617328
rect 173838 617248 173872 617328
rect 174496 617248 174530 617328
rect 175154 617248 175188 617328
rect 175812 617248 175846 617328
rect 175930 617266 175960 617300
rect 172408 617226 175846 617248
rect 175926 617233 175930 617236
rect 172408 617224 175852 617226
rect 172408 617214 175858 617224
rect 171694 616844 172142 617006
rect 171618 616794 172142 616844
rect 171618 616690 171772 616794
rect 167606 615738 170925 616358
rect 140998 615297 141618 615682
rect 141668 615634 142234 615668
rect 141668 615502 141702 615634
rect 141823 615564 141860 615588
rect 142040 615565 142079 615588
rect 142039 615564 142079 615565
rect 142039 615560 142050 615564
rect 141723 615502 141804 615539
rect 141851 615536 141860 615560
rect 142039 615554 142051 615560
rect 141863 615539 142051 615554
rect 141863 615536 142132 615539
rect 141863 615520 142050 615536
rect 142051 615502 142132 615536
rect 142200 615502 142234 615634
rect 167614 615573 170925 615738
rect 172408 616590 172442 617214
rect 172522 616590 172556 617214
rect 172568 617202 172569 617203
rect 173167 617202 173168 617203
rect 172567 617201 172568 617202
rect 173168 617201 173169 617202
rect 172567 616602 172568 616603
rect 173168 616602 173169 616603
rect 172568 616601 172569 616602
rect 173167 616601 173168 616602
rect 173180 616590 173214 617214
rect 173226 617202 173227 617203
rect 173825 617202 173826 617203
rect 173225 617201 173226 617202
rect 173826 617201 173827 617202
rect 173225 616602 173226 616603
rect 173826 616602 173827 616603
rect 173226 616601 173227 616602
rect 173825 616601 173826 616602
rect 173838 616590 173872 617214
rect 173884 617202 173885 617203
rect 174483 617202 174484 617203
rect 173883 617201 173884 617202
rect 174484 617201 174485 617202
rect 173883 616602 173884 616603
rect 174484 616602 174485 616603
rect 173884 616601 173885 616602
rect 174483 616601 174484 616602
rect 174496 616590 174530 617214
rect 174542 617202 174543 617203
rect 175141 617202 175142 617203
rect 174541 617201 174542 617202
rect 175142 617201 175143 617202
rect 175136 616603 175142 616624
rect 174541 616602 174542 616603
rect 175136 616602 175143 616603
rect 174542 616601 174543 616602
rect 175136 616590 175142 616602
rect 175154 616590 175188 617214
rect 175200 617202 175201 617203
rect 175799 617202 175800 617203
rect 175199 617201 175200 617202
rect 175800 617201 175801 617202
rect 175812 617198 175858 617214
rect 175862 617198 175880 617202
rect 175812 617186 175880 617198
rect 175812 617130 175884 617186
rect 175812 616682 175858 617130
rect 175862 616682 175884 617130
rect 175812 616618 175884 616682
rect 175812 616606 175880 616618
rect 175199 616602 175200 616603
rect 175800 616602 175801 616603
rect 175200 616601 175201 616602
rect 175799 616601 175800 616602
rect 175812 616590 175858 616606
rect 175862 616602 175880 616606
rect 175892 616602 175896 617202
rect 175926 616618 175943 617233
rect 172408 616587 175858 616590
rect 172408 616578 175852 616587
rect 172408 616568 175846 616578
rect 175926 616575 175930 616618
rect 172408 616566 175852 616568
rect 172408 616556 175858 616566
rect 172408 615932 172442 616556
rect 172522 615932 172556 616556
rect 172568 616544 172569 616545
rect 173167 616544 173168 616545
rect 172567 616543 172568 616544
rect 173168 616543 173169 616544
rect 172567 615944 172568 615945
rect 173168 615944 173169 615945
rect 172568 615943 172569 615944
rect 173167 615943 173168 615944
rect 173180 615932 173214 616556
rect 173226 616544 173227 616545
rect 173825 616544 173826 616545
rect 173225 616543 173226 616544
rect 173826 616543 173827 616544
rect 173225 615944 173226 615945
rect 173826 615944 173827 615945
rect 173226 615943 173227 615944
rect 173825 615943 173826 615944
rect 173838 615932 173872 616556
rect 173884 616544 173885 616545
rect 174483 616544 174484 616545
rect 173883 616543 173884 616544
rect 174484 616543 174485 616544
rect 173883 615944 173884 615945
rect 174484 615944 174485 615945
rect 173884 615943 173885 615944
rect 174483 615943 174484 615944
rect 174496 615932 174530 616556
rect 174542 616544 174543 616545
rect 175136 616544 175142 616556
rect 174541 616543 174542 616544
rect 175136 616543 175143 616544
rect 175136 616538 175142 616543
rect 174541 615944 174542 615945
rect 175142 615944 175143 615945
rect 174542 615943 174543 615944
rect 175141 615943 175142 615944
rect 175154 615932 175188 616556
rect 175200 616544 175201 616545
rect 175799 616544 175800 616545
rect 175199 616543 175200 616544
rect 175800 616543 175801 616544
rect 175812 616540 175858 616556
rect 175862 616540 175880 616544
rect 175812 616528 175880 616540
rect 175812 616478 175884 616528
rect 175812 616030 175858 616478
rect 175862 616030 175884 616478
rect 175812 615960 175884 616030
rect 175812 615948 175880 615960
rect 175199 615944 175200 615945
rect 175800 615944 175801 615945
rect 175200 615943 175201 615944
rect 175799 615943 175800 615944
rect 175812 615932 175858 615948
rect 175862 615944 175880 615948
rect 175892 615944 175896 616544
rect 175926 615960 175943 616575
rect 172408 615929 175858 615932
rect 172408 615920 175852 615929
rect 172408 615910 175846 615920
rect 175926 615917 175930 615960
rect 172408 615908 175852 615910
rect 172408 615898 175858 615908
rect 172408 615666 172442 615898
rect 172522 615818 172556 615898
rect 172568 615886 172569 615887
rect 173167 615886 173168 615887
rect 172567 615885 172568 615886
rect 173168 615885 173169 615886
rect 173180 615818 173214 615898
rect 173226 615886 173227 615887
rect 173825 615886 173826 615887
rect 173225 615885 173226 615886
rect 173826 615885 173827 615886
rect 173306 615834 173754 615842
rect 173838 615818 173872 615898
rect 173884 615886 173885 615887
rect 174483 615886 174484 615887
rect 173883 615885 173884 615886
rect 174484 615885 174485 615886
rect 174496 615818 174530 615898
rect 174542 615886 174543 615887
rect 175141 615886 175142 615887
rect 174541 615885 174542 615886
rect 175142 615885 175143 615886
rect 175154 615818 175188 615898
rect 175200 615886 175201 615887
rect 175799 615886 175800 615887
rect 175199 615885 175200 615886
rect 175800 615885 175801 615886
rect 175812 615882 175858 615898
rect 175862 615882 175880 615886
rect 175812 615870 175880 615882
rect 175812 615818 175884 615870
rect 175824 615814 175884 615818
rect 173278 615806 173782 615814
rect 175824 615806 175858 615814
rect 173152 615768 173190 615806
rect 173810 615768 173848 615806
rect 174468 615768 174506 615806
rect 175126 615768 175164 615806
rect 175784 615768 175822 615806
rect 175828 615802 175846 615806
rect 175862 615780 175884 615814
rect 175862 615768 175880 615780
rect 172584 615734 173190 615768
rect 173242 615734 173848 615768
rect 173900 615734 174506 615768
rect 174558 615734 175164 615768
rect 175216 615734 175822 615768
rect 175892 615670 175896 615886
rect 175926 615666 175943 615917
rect 172408 615632 175943 615666
rect 175964 615632 175998 617328
rect 176570 616974 176604 618300
rect 187356 618292 189496 618326
rect 187899 618108 187933 618292
rect 179746 617812 179762 617814
rect 179654 617703 180274 617812
rect 180386 617798 180828 617832
rect 180324 617771 180890 617798
rect 179654 617669 185078 617703
rect 179654 617633 180274 617669
rect 180324 617504 180358 617669
rect 180426 617635 180460 617638
rect 180754 617635 180788 617638
rect 180856 617504 180890 617669
rect 187344 617633 187969 618108
rect 176684 616974 176708 617008
rect 180166 616988 180200 617128
rect 180342 617088 185078 617122
rect 180246 617060 180348 617078
rect 180274 617032 180320 617050
rect 180280 616988 180314 617022
rect 185338 616988 185372 617022
rect 185452 616988 185486 617128
rect 187380 616988 187414 617633
rect 188724 617612 188744 617894
rect 187494 616988 187528 617022
rect 176476 616940 176770 616974
rect 179644 616954 187896 616988
rect 176570 616906 176604 616940
rect 176570 616838 176628 616906
rect 176702 616878 176718 616912
rect 176570 616578 176604 616838
rect 176622 616603 176638 616779
rect 176646 616603 176656 616779
rect 176672 616591 176722 616845
rect 176570 616510 176628 616578
rect 176684 616565 176694 616591
rect 176570 616442 176604 616510
rect 176684 616442 176708 616476
rect 176736 616442 176770 616940
rect 176476 616408 176770 616442
rect 176570 616358 176604 616408
rect 176534 615994 176784 616358
rect 176714 615808 176748 615820
rect 176492 615774 176748 615808
rect 179548 615766 179582 616892
rect 180166 616874 180200 616954
rect 180280 616874 180314 616954
rect 185338 616874 185372 616954
rect 185452 616874 185486 616954
rect 180166 616840 185486 616874
rect 180166 616110 180200 616840
rect 180280 616262 180314 616840
rect 180326 616828 180327 616829
rect 185325 616828 185326 616829
rect 180325 616827 180326 616828
rect 185326 616827 185327 616828
rect 180280 616246 180314 616250
rect 181350 616246 181390 616254
rect 181406 616246 181418 616282
rect 185338 616262 185372 616840
rect 185338 616246 185372 616250
rect 180308 616220 185344 616246
rect 180304 616216 185348 616220
rect 180246 616212 185406 616216
rect 180304 616182 185348 616212
rect 180326 616178 185348 616182
rect 180326 616170 185326 616178
rect 181350 616146 181390 616170
rect 181406 616156 181418 616170
rect 185452 616110 185486 616840
rect 187380 616758 187414 616954
rect 187482 616898 187540 616940
rect 187494 616894 187528 616898
rect 187522 616886 187710 616894
rect 187522 616880 187722 616886
rect 187460 616874 187722 616880
rect 187456 616872 187722 616874
rect 187460 616860 187722 616872
rect 187518 616850 187722 616860
rect 187518 616840 187832 616850
rect 187540 616828 187832 616840
rect 187556 616826 187832 616828
rect 187760 616758 187794 616812
rect 187862 616758 187896 616954
rect 187380 616724 188204 616758
rect 187760 616264 187794 616724
rect 187862 616264 187896 616724
rect 190646 616518 190648 617906
rect 190622 616312 190648 616518
rect 190646 616306 190648 616312
rect 190972 617038 196892 619780
rect 197361 617038 197395 621336
rect 199468 621332 199489 621336
rect 197475 621299 197522 621315
rect 197463 621234 197522 621299
rect 198133 621284 198180 621315
rect 198791 621284 198838 621315
rect 199449 621284 199496 621315
rect 198121 621268 198180 621284
rect 198779 621268 198838 621284
rect 199437 621268 199496 621284
rect 197572 621234 198180 621268
rect 198230 621234 198838 621268
rect 198888 621234 199496 621268
rect 197463 621225 197498 621234
rect 198121 621225 198156 621234
rect 198779 621225 198814 621234
rect 199437 621225 199472 621234
rect 197463 621187 197509 621225
rect 197414 617146 197440 617262
rect 197442 617187 197468 617234
rect 197475 617187 197509 621187
rect 197510 621186 197543 621191
rect 198121 621187 198167 621225
rect 197510 618822 197544 621186
rect 197510 617199 197555 618822
rect 197564 617190 197568 617402
rect 197592 617187 197596 617430
rect 198133 617187 198167 621187
rect 198168 621186 198201 621191
rect 198779 621187 198825 621225
rect 198168 618822 198202 621186
rect 198791 620144 198825 621187
rect 198757 619476 198768 620144
rect 198785 619476 198825 620144
rect 198168 617199 198213 618822
rect 198791 618288 198825 619476
rect 198757 617222 198768 618288
rect 198785 617222 198825 618288
rect 198791 617187 198825 617222
rect 198826 621186 198859 621191
rect 199437 621187 199483 621225
rect 198826 618822 198860 621186
rect 199387 619476 199418 620144
rect 199443 619476 199446 620144
rect 198826 617199 198871 618822
rect 198884 617192 198894 617400
rect 198912 617187 198922 617428
rect 199387 617187 199418 618288
rect 199443 617187 199446 618288
rect 199449 617187 199483 621187
rect 199484 621186 199517 621191
rect 199484 618822 199518 621186
rect 199484 617199 199529 618822
rect 197442 617146 197522 617187
rect 197463 617106 197522 617146
rect 197525 617140 198180 617187
rect 198183 617140 198838 617187
rect 198841 617140 199496 617187
rect 197463 617090 197498 617106
rect 197463 617075 197478 617090
rect 197532 617072 197550 617140
rect 197560 617106 198180 617140
rect 198230 617106 198838 617140
rect 197560 617100 197578 617106
rect 198121 617090 198156 617106
rect 198779 617090 198814 617106
rect 198848 617072 198858 617140
rect 198876 617100 198886 617140
rect 198888 617106 199496 617140
rect 199437 617090 199489 617106
rect 199468 617038 199489 617090
rect 199598 617038 199632 621336
rect 190972 617007 199632 617038
rect 200107 617007 200141 621677
rect 200247 617007 200281 621677
rect 200361 618822 200395 621677
rect 200580 619534 200582 619690
rect 200765 618822 200799 621677
rect 200361 617007 200406 618822
rect 200765 617007 200810 618822
rect 200879 617007 200913 621677
rect 201652 620154 201711 620188
rect 202297 620164 202312 620246
rect 201590 620120 201980 620154
rect 202335 620126 202350 620284
rect 200916 619476 200926 619672
rect 201590 619622 201624 620120
rect 201677 619959 201711 620120
rect 201804 620052 201851 620099
rect 201766 620018 201851 620052
rect 201723 619959 201738 619970
rect 201821 619959 201866 619970
rect 201677 619783 201738 619959
rect 201832 619783 201866 619959
rect 201677 619656 201711 619783
rect 201804 619724 201851 619771
rect 201766 619690 201851 619724
rect 201652 619622 201711 619656
rect 201946 619622 201980 620120
rect 200972 619476 200982 619616
rect 201590 619588 201980 619622
rect 201576 618918 201998 619538
rect 202301 619476 202328 619628
rect 202329 619476 202375 619684
rect 201578 617946 201584 618202
rect 201606 617974 201612 618174
rect 190972 617004 200913 617007
rect 190972 616664 196892 617004
rect 197361 616911 197395 617004
rect 197443 616973 200913 617004
rect 190972 616444 196902 616664
rect 187682 616250 188074 616264
rect 187618 616238 188074 616250
rect 187682 616222 188074 616238
rect 188748 616228 189294 616264
rect 189844 616234 190170 616264
rect 190506 616234 190836 616264
rect 187590 616216 188074 616222
rect 187590 616210 187722 616216
rect 187862 616208 187896 616216
rect 187682 616160 188130 616208
rect 188720 616200 189322 616208
rect 189816 616206 190170 616208
rect 190506 616206 190864 616208
rect 180166 616076 185486 616110
rect 176642 615732 186894 615766
rect 179548 615652 179582 615732
rect 186860 615676 186894 615732
rect 179619 615656 179722 615664
rect 179612 615652 179722 615656
rect 186708 615652 186719 615663
rect 186720 615656 186894 615676
rect 179514 615618 186719 615652
rect 141668 615481 142324 615502
rect 141634 615447 142324 615481
rect 152664 615458 154304 615478
rect 141668 615435 142324 615447
rect 141670 615428 142324 615435
rect 141847 615413 142055 615426
rect 141851 615401 142051 615413
rect 141668 615374 141702 615401
rect 141847 615392 142055 615401
rect 141851 615380 142051 615392
rect 142200 615374 142234 615401
rect 141813 615366 142089 615367
rect 141702 615333 142200 615366
rect 141702 615299 142200 615312
rect 129524 614809 129558 614843
rect 132582 614809 132616 614843
rect 135640 614809 135674 614843
rect 135754 614809 135788 615054
rect 127997 614775 136267 614809
rect 127997 614196 128031 614775
rect 129524 614695 129558 614775
rect 132582 614695 132616 614775
rect 135640 614695 135674 614775
rect 135754 614695 135788 614775
rect 128052 614633 128133 614680
rect 128192 614661 135788 614695
rect 129511 614649 129512 614650
rect 129512 614648 129513 614649
rect 128099 614196 128133 614633
rect 129180 614620 129236 614634
rect 129524 614196 129558 614661
rect 129570 614649 129571 614650
rect 132569 614649 132570 614650
rect 129569 614648 129570 614649
rect 132570 614648 132571 614649
rect 129754 614620 129810 614634
rect 132582 614196 132616 614661
rect 132628 614649 132629 614650
rect 135627 614649 135628 614650
rect 132627 614648 132628 614649
rect 135628 614648 135629 614649
rect 135640 614196 135674 614661
rect 135754 614196 135788 614661
rect 125438 614132 141752 614196
rect 127997 614116 128031 614132
rect 128099 614116 128133 614132
rect 129524 614116 129558 614132
rect 132582 614116 132616 614132
rect 135332 614130 135388 614132
rect 135640 614116 135674 614132
rect 135754 614116 135788 614132
rect 125438 614052 141832 614116
rect 127997 611291 128031 614052
rect 129512 614049 129513 614050
rect 129511 614048 129512 614049
rect 129524 614037 129558 614052
rect 129569 614049 129570 614050
rect 132570 614049 132571 614050
rect 129570 614048 129571 614049
rect 132569 614048 132570 614049
rect 132582 614037 132616 614052
rect 132627 614049 132628 614050
rect 135628 614049 135629 614050
rect 132628 614048 132629 614049
rect 135627 614048 135628 614049
rect 135640 614037 135674 614052
rect 135754 614037 135788 614052
rect 128052 613975 128133 614022
rect 128192 614003 135788 614037
rect 129511 613991 129512 613992
rect 129512 613990 129513 613991
rect 128099 613407 128133 613975
rect 129524 613784 129558 614003
rect 129570 613991 129571 613992
rect 132569 613991 132570 613992
rect 129569 613990 129570 613991
rect 132570 613990 132571 613991
rect 129180 613472 129236 613476
rect 129180 613416 129236 613420
rect 129410 613400 129618 613784
rect 129754 613472 129810 613476
rect 129754 613416 129810 613420
rect 128908 613396 129618 613400
rect 128908 613379 129562 613396
rect 129569 613391 129570 613392
rect 132570 613391 132571 613392
rect 129570 613390 129571 613391
rect 132569 613390 132570 613391
rect 132582 613379 132616 614003
rect 132628 613991 132629 613992
rect 135627 613991 135628 613992
rect 132627 613990 132628 613991
rect 135628 613990 135629 613991
rect 135332 613952 135388 613976
rect 135332 613896 135388 613920
rect 132627 613391 132628 613392
rect 135628 613391 135629 613392
rect 132628 613390 132629 613391
rect 135627 613390 135628 613391
rect 135640 613379 135674 614003
rect 135754 613379 135788 614003
rect 144760 613778 145208 613858
rect 144758 613646 145208 613778
rect 144758 613550 144878 613646
rect 128052 613317 128133 613364
rect 128192 613345 135788 613379
rect 128908 613326 129562 613345
rect 129570 613333 129571 613334
rect 132569 613333 132570 613334
rect 129569 613332 129570 613333
rect 132570 613332 132571 613333
rect 128099 612749 128133 613317
rect 129180 613312 129236 613314
rect 129180 613256 129236 613258
rect 129362 612746 129518 612755
rect 129512 612733 129513 612734
rect 129511 612732 129512 612733
rect 129334 612721 129518 612727
rect 129524 612721 129558 613326
rect 129754 613312 129810 613314
rect 129754 613256 129810 613258
rect 129564 612746 129658 612755
rect 129569 612733 129570 612734
rect 132570 612733 132571 612734
rect 129570 612732 129571 612733
rect 132569 612732 132570 612733
rect 129564 612721 129686 612727
rect 132582 612721 132616 613345
rect 132628 613333 132629 613334
rect 135627 613333 135628 613334
rect 132627 613332 132628 613333
rect 135628 613332 135629 613333
rect 135332 612810 135388 612826
rect 135534 612780 135634 612798
rect 135332 612754 135388 612770
rect 135506 612752 135634 612770
rect 132627 612733 132628 612734
rect 135628 612733 135629 612734
rect 132628 612732 132629 612733
rect 135627 612732 135628 612733
rect 135640 612721 135674 613345
rect 135754 612798 135788 613345
rect 135680 612780 135788 612798
rect 135754 612770 135788 612780
rect 135680 612752 135788 612770
rect 135754 612721 135788 612752
rect 128052 612659 128133 612706
rect 128192 612687 135788 612721
rect 129511 612675 129512 612676
rect 129512 612674 129513 612675
rect 128099 612091 128133 612659
rect 129180 612140 129236 612156
rect 129180 612084 129236 612100
rect 129512 612075 129513 612076
rect 129511 612074 129512 612075
rect 129524 612063 129558 612687
rect 129570 612675 129571 612676
rect 132569 612675 132570 612676
rect 129569 612674 129570 612675
rect 132570 612674 132571 612675
rect 129754 612140 129810 612156
rect 129754 612084 129810 612100
rect 129569 612075 129570 612076
rect 132570 612075 132571 612076
rect 129570 612074 129571 612075
rect 132569 612074 132570 612075
rect 132582 612063 132616 612687
rect 132628 612675 132629 612676
rect 135627 612675 135628 612676
rect 132627 612674 132628 612675
rect 135628 612674 135629 612675
rect 135332 612642 135388 612644
rect 135332 612586 135388 612588
rect 132627 612075 132628 612076
rect 135628 612075 135629 612076
rect 132628 612074 132629 612075
rect 135627 612074 135628 612075
rect 135640 612063 135674 612687
rect 135754 612063 135788 612687
rect 128052 612001 128133 612048
rect 128192 612029 135788 612063
rect 129511 612017 129512 612018
rect 129512 612016 129513 612017
rect 128099 611433 128133 612001
rect 129512 611417 129513 611418
rect 129511 611416 129512 611417
rect 129524 611405 129558 612029
rect 129570 612017 129571 612018
rect 132569 612017 132570 612018
rect 129569 612016 129570 612017
rect 132570 612016 132571 612017
rect 129569 611417 129570 611418
rect 132570 611417 132571 611418
rect 129570 611416 129571 611417
rect 132569 611416 132570 611417
rect 132582 611405 132616 612029
rect 132628 612017 132629 612018
rect 135627 612017 135628 612018
rect 132627 612016 132628 612017
rect 135628 612016 135629 612017
rect 135332 611488 135388 611504
rect 135332 611432 135388 611448
rect 132627 611417 132628 611418
rect 135628 611417 135629 611418
rect 132628 611416 132629 611417
rect 135627 611416 135628 611417
rect 135640 611405 135674 612029
rect 135754 611405 135788 612029
rect 149206 611544 149240 614762
rect 152684 614116 152685 615458
rect 154284 614116 154304 615458
rect 167768 615320 167792 615336
rect 167746 615290 167792 615320
rect 167718 615262 167820 615264
rect 179548 615194 179582 615618
rect 179634 615606 179722 615618
rect 179650 615586 179684 615606
rect 186720 615590 186792 615628
rect 186758 615570 186792 615590
rect 186720 615558 186808 615570
rect 179612 615496 179684 615534
rect 179734 615524 186808 615558
rect 186720 615512 186808 615524
rect 179650 615206 179684 615496
rect 186758 615222 186792 615512
rect 179634 615198 179722 615206
rect 179612 615194 179722 615198
rect 186708 615194 186719 615205
rect 179514 615160 186719 615194
rect 179548 615080 179582 615160
rect 179619 615148 179722 615160
rect 186860 615080 186894 615656
rect 176642 615046 186894 615080
rect 152684 613846 154284 613866
rect 152684 613769 152685 613846
rect 154284 613769 154304 613846
rect 152684 613768 154304 613769
rect 179548 613532 179582 615046
rect 187862 613532 187896 616160
rect 190972 615860 196892 616444
rect 190972 615844 196932 615860
rect 190972 615596 196892 615844
rect 196932 615780 196948 615844
rect 197180 615780 197184 615860
rect 190972 615493 196893 615596
rect 196931 615532 196932 615533
rect 196932 615531 196933 615532
rect 196946 615493 196973 615536
rect 190972 615492 196892 615493
rect 190972 615172 197116 615492
rect 197347 615409 197395 616911
rect 197475 616921 197509 616973
rect 198133 616952 198167 616973
rect 198791 616952 198825 616973
rect 199449 616952 199489 616973
rect 200107 616952 200141 616973
rect 198091 616921 198167 616952
rect 198749 616921 198825 616952
rect 199407 616921 199489 616952
rect 200065 616921 200141 616952
rect 197475 616824 197521 616921
rect 198091 616905 198179 616921
rect 198749 616905 198837 616921
rect 199407 616905 199495 616921
rect 200065 616905 200153 616921
rect 200247 616905 200281 616973
rect 200361 616970 200406 616973
rect 200765 616970 200810 616973
rect 200361 616952 200395 616970
rect 200765 616952 200799 616970
rect 200361 616905 200408 616952
rect 200723 616905 200799 616952
rect 197523 616871 198179 616905
rect 198181 616871 198837 616905
rect 198839 616871 199495 616905
rect 199497 616871 200153 616905
rect 200155 616871 200799 616905
rect 198099 616865 198103 616871
rect 198127 616837 198131 616871
rect 198133 616824 198179 616871
rect 198791 616824 198837 616871
rect 199415 616865 199419 616871
rect 199443 616837 199447 616871
rect 199449 616824 199495 616871
rect 200107 616824 200153 616871
rect 197475 616812 197509 616824
rect 198108 616812 198121 616823
rect 198133 616812 198167 616824
rect 198766 616812 198779 616823
rect 198791 616812 198825 616824
rect 199424 616812 199437 616823
rect 199449 616812 199489 616824
rect 200082 616812 200095 616823
rect 200107 616812 200141 616824
rect 197461 615508 197509 616812
rect 198119 615508 198167 616812
rect 198777 615508 198825 616812
rect 197461 615436 197495 615508
rect 198119 615496 198153 615508
rect 198777 615496 198811 615508
rect 197497 615436 197501 615483
rect 197525 615449 197529 615455
rect 198105 615449 198153 615496
rect 198763 615449 198811 615496
rect 190972 615171 196892 615172
rect 190972 615064 196893 615171
rect 196932 615132 196933 615133
rect 196931 615131 196932 615132
rect 196946 615124 196973 615171
rect 190972 613860 196892 615064
rect 183764 612558 184402 612801
rect 180862 612432 181050 612458
rect 180834 612404 181022 612430
rect 179284 612357 179299 612397
rect 187433 611917 187467 612415
rect 179525 611883 187795 611917
rect 179284 611699 179299 611745
rect 128192 611371 135788 611405
rect 129524 611291 129558 611371
rect 132582 611291 132616 611371
rect 135640 611291 135674 611371
rect 135754 611291 135788 611371
rect 148716 611510 150968 611544
rect 148716 611454 148750 611510
rect 149104 611466 149138 611510
rect 148716 611430 149054 611454
rect 149206 611430 149240 611510
rect 148716 611420 149240 611430
rect 148716 611340 148750 611420
rect 148902 611396 149240 611420
rect 148818 611368 148852 611374
rect 149206 611340 149240 611396
rect 144758 611306 149240 611340
rect 127997 611257 136267 611291
rect 135754 610698 135788 611257
rect 143502 610682 143758 610708
rect 143530 610654 143730 610680
rect 131602 610172 132222 610594
rect 132582 610580 132616 610614
rect 132272 610546 132838 610580
rect 132272 610224 132306 610546
rect 132327 610444 132408 610451
rect 132327 610404 132416 610444
rect 132374 610366 132416 610404
rect 132394 610324 132416 610366
rect 132422 610296 132444 610472
rect 132582 610466 132616 610546
rect 132643 610466 132654 610477
rect 132467 610432 132654 610466
rect 132569 610420 132570 610421
rect 132570 610419 132571 610420
rect 132570 610350 132571 610351
rect 132569 610349 132570 610350
rect 132582 610338 132616 610432
rect 132628 610420 132629 610421
rect 132627 610419 132628 610420
rect 132655 610404 132736 610451
rect 132702 610366 132736 610404
rect 132627 610350 132628 610351
rect 132628 610349 132629 610350
rect 132643 610338 132654 610349
rect 132467 610304 132654 610338
rect 132582 610224 132616 610304
rect 132804 610224 132838 610546
rect 144474 610450 144828 610872
rect 148716 610698 148750 611306
rect 179525 611178 179559 611883
rect 185570 611837 186026 611865
rect 179680 611832 180862 611837
rect 181062 611832 186026 611837
rect 187378 611832 187384 611837
rect 179708 611804 180862 611809
rect 181062 611804 186026 611809
rect 186386 611803 186842 611824
rect 187284 611809 187396 611815
rect 187284 611804 187412 611809
rect 187284 611803 187396 611804
rect 179720 611800 187396 611803
rect 179580 611751 179661 611788
rect 179720 611773 187381 611800
rect 179704 611769 187381 611773
rect 179708 611763 180862 611769
rect 181062 611763 185626 611769
rect 186386 611756 186842 611769
rect 187284 611757 187381 611769
rect 186000 611754 186842 611756
rect 179580 611745 179708 611751
rect 179580 611739 180862 611745
rect 181062 611739 185626 611745
rect 186000 611739 186456 611754
rect 187272 611739 187283 611750
rect 179580 611735 187288 611739
rect 179580 611714 187283 611735
rect 187284 611714 187365 611724
rect 179580 611705 187365 611714
rect 179586 611699 180862 611705
rect 181062 611699 185626 611705
rect 179611 611693 179708 611699
rect 179614 611671 179621 611686
rect 179627 611207 179661 611693
rect 186000 611686 186456 611705
rect 186978 611699 187365 611705
rect 187284 611686 187365 611699
rect 179667 611671 180862 611686
rect 181062 611671 185626 611686
rect 186978 611677 187365 611686
rect 186978 611671 187312 611677
rect 183442 611502 183890 611574
rect 183018 611362 183890 611502
rect 183018 611290 183466 611362
rect 179627 611178 180010 611207
rect 179525 611174 180010 611178
rect 181412 611174 187325 611179
rect 179284 611041 179299 611087
rect 132272 610190 132838 610224
rect 138832 610114 138888 610126
rect 139280 610114 139336 610126
rect 140524 610114 140580 610126
rect 138832 610058 138888 610070
rect 139280 610058 139336 610070
rect 140524 610058 140580 610070
rect 144758 609787 144792 610450
rect 148680 609787 149271 609823
rect 140869 609776 144717 609787
rect 127984 608920 135824 609774
rect 140869 609764 144706 609776
rect 140869 609753 144717 609764
rect 144758 609753 149271 609787
rect 140869 609468 140903 609753
rect 144609 609673 144721 609685
rect 141064 609670 144721 609673
rect 140924 609611 141005 609658
rect 141064 609639 144706 609670
rect 144609 609627 144706 609639
rect 138832 609454 138888 609468
rect 139280 609454 139336 609468
rect 140524 609454 140580 609468
rect 140869 609454 140958 609468
rect 138832 609398 138888 609412
rect 139280 609398 139336 609412
rect 140524 609398 140580 609412
rect 140869 609406 140903 609454
rect 140971 609419 141005 609611
rect 144656 609434 144690 609627
rect 140835 609372 140903 609406
rect 140924 609418 141005 609419
rect 140924 609406 141052 609418
rect 144597 609406 144608 609417
rect 140924 609372 144608 609406
rect 126528 608886 135824 608920
rect 127984 608748 135824 608886
rect 138832 608794 138888 608810
rect 139280 608794 139336 608810
rect 140524 608794 140580 608810
rect 140869 608754 140903 609372
rect 140955 609360 141052 609372
rect 140971 609043 141005 609360
rect 144609 609344 144690 609391
rect 144656 609028 144690 609344
rect 144609 609027 144690 609028
rect 144609 609015 144706 609027
rect 140924 608953 141005 609000
rect 141064 608981 144706 609015
rect 144609 608969 144706 608981
rect 140971 608761 141005 608953
rect 144656 608776 144690 608969
rect 140924 608760 141005 608761
rect 140924 608754 141052 608760
rect 138832 608738 138888 608754
rect 139280 608738 139336 608754
rect 140524 608738 140580 608754
rect 140869 608748 141052 608754
rect 144597 608748 144608 608759
rect 140835 608738 144608 608748
rect 140835 608714 140903 608738
rect 140924 608714 144608 608738
rect 140869 608634 140903 608714
rect 140940 608702 141052 608714
rect 144758 608634 144792 609753
rect 138522 608600 144792 608634
rect 140869 608206 140903 608600
rect 127984 606150 135860 608200
rect 138522 608172 144792 608206
rect 140869 608092 140903 608172
rect 140835 608058 140903 608092
rect 140924 608092 141052 608104
rect 144597 608092 144608 608103
rect 140924 608058 144608 608092
rect 140869 608056 140903 608058
rect 140955 608056 141052 608058
rect 138832 608052 138888 608056
rect 139280 608052 139336 608056
rect 140524 608052 140580 608056
rect 140869 608052 141052 608056
rect 138832 607996 138888 608000
rect 139280 607996 139336 608000
rect 140524 607996 140580 608000
rect 140869 607496 140903 608052
rect 140955 608046 141052 608052
rect 140971 607727 141005 608046
rect 144609 608030 144690 608077
rect 144656 607712 144690 608030
rect 144609 607711 144690 607712
rect 144609 607699 144706 607711
rect 140924 607637 141005 607684
rect 141064 607665 144706 607699
rect 144609 607653 144706 607665
rect 138832 607494 138888 607496
rect 139280 607494 139336 607496
rect 140524 607494 140580 607496
rect 140869 607494 140942 607496
rect 140869 607440 140903 607494
rect 140971 607447 141005 607637
rect 144656 607462 144690 607653
rect 140924 607446 141005 607447
rect 140924 607440 141052 607446
rect 138832 607438 138888 607440
rect 139280 607438 139336 607440
rect 140524 607438 140580 607440
rect 140869 607438 141052 607440
rect 140869 607434 140903 607438
rect 140835 607400 140903 607434
rect 140924 607434 141052 607438
rect 144597 607434 144608 607445
rect 140924 607400 144608 607434
rect 139280 606830 139336 606838
rect 140524 606830 140580 606838
rect 140869 606782 140903 607400
rect 140955 607388 141052 607400
rect 140971 607069 141005 607388
rect 144609 607372 144690 607419
rect 144656 607054 144690 607372
rect 144609 607053 144690 607054
rect 144609 607041 144706 607053
rect 140924 606979 141005 607026
rect 141064 607007 144706 607041
rect 144609 606995 144706 607007
rect 140971 606789 141005 606979
rect 144656 606804 144690 606995
rect 140924 606788 141005 606789
rect 140924 606782 141052 606788
rect 138832 606774 138888 606782
rect 139280 606774 139336 606782
rect 140524 606774 140580 606782
rect 140869 606776 141052 606782
rect 144597 606776 144608 606787
rect 140835 606774 144608 606776
rect 140835 606742 140903 606774
rect 140924 606742 144608 606774
rect 140869 606688 140903 606742
rect 140955 606730 141052 606742
rect 138832 606680 138888 606688
rect 139280 606680 139336 606688
rect 140524 606680 140580 606688
rect 140869 606680 140958 606688
rect 140869 606269 140903 606680
rect 140971 606411 141005 606730
rect 144609 606714 144690 606761
rect 144656 606396 144690 606714
rect 144609 606395 144690 606396
rect 144609 606383 144706 606395
rect 141064 606352 144706 606383
rect 141064 606349 144721 606352
rect 144609 606337 144721 606349
rect 144758 606269 144792 608172
rect 148680 606269 149271 609753
rect 150928 609414 150962 610698
rect 179284 610383 179299 610429
rect 179525 609858 179559 611174
rect 179621 611161 179667 611174
rect 179708 611146 180010 611151
rect 180416 611145 181070 611164
rect 187331 611158 187365 611677
rect 187284 611157 187365 611158
rect 187284 611151 187381 611157
rect 181412 611146 187381 611151
rect 185570 611145 187034 611146
rect 187284 611145 187381 611146
rect 179580 611093 179661 611130
rect 179720 611115 187381 611145
rect 179704 611111 187381 611115
rect 180416 611102 181070 611111
rect 181412 611105 187381 611111
rect 179580 611081 179708 611093
rect 180012 611090 181070 611102
rect 187284 611099 187381 611105
rect 180012 611081 180666 611090
rect 187272 611087 187283 611092
rect 181412 611081 187284 611087
rect 179580 611077 187288 611081
rect 179580 611066 187284 611077
rect 179580 611047 187365 611066
rect 179611 611035 179708 611047
rect 179627 610515 179661 611035
rect 180012 611028 180666 611047
rect 181010 611041 187365 611047
rect 187284 611034 187365 611041
rect 181010 611019 187365 611034
rect 181010 611013 187312 611019
rect 181010 610985 181468 611013
rect 183442 610856 183890 610928
rect 183026 610716 183890 610856
rect 183026 610698 183474 610716
rect 185576 610521 186056 610549
rect 179680 610512 186056 610521
rect 179708 610487 186056 610493
rect 186408 610487 186864 610502
rect 187331 610500 187365 611019
rect 187284 610499 187365 610500
rect 187284 610487 187381 610499
rect 187433 610487 187467 611883
rect 197347 610698 197381 615409
rect 197461 615347 197501 615436
rect 197521 615436 197529 615449
rect 197537 615436 198153 615449
rect 197521 615415 198153 615436
rect 198179 615415 198187 615449
rect 198195 615415 198811 615449
rect 197525 615409 197578 615415
rect 197520 615381 197578 615408
rect 198107 615399 198153 615415
rect 198765 615399 198811 615415
rect 197520 615347 197529 615381
rect 198119 615347 198153 615399
rect 198777 615347 198811 615399
rect 198813 615381 198817 615483
rect 199358 615455 199360 616552
rect 199435 616524 199489 616812
rect 199386 615455 199388 616524
rect 199435 615496 199514 616524
rect 199421 615455 199514 615496
rect 199524 615455 199542 616552
rect 200093 615508 200141 616812
rect 200247 615643 200281 616871
rect 200361 615804 200395 616871
rect 200765 616823 200799 616871
rect 200740 616812 200799 616823
rect 200751 615792 200799 616812
rect 200751 615745 200811 615792
rect 200423 615711 200811 615745
rect 200680 615643 200682 615698
rect 200708 615643 200738 615698
rect 200751 615680 200811 615711
rect 200751 615643 200799 615680
rect 200865 615643 200913 616973
rect 201580 616574 201584 617574
rect 201656 616548 201730 617174
rect 201642 616394 201796 616548
rect 201560 616318 201584 616374
rect 201580 616060 201584 616318
rect 202301 615764 202320 618288
rect 202329 615792 202375 618288
rect 202396 617048 203835 621700
rect 205178 620542 205212 621700
rect 204440 619848 204902 620486
rect 205112 620460 205212 620542
rect 204530 619798 204554 619848
rect 204564 619798 204588 619848
rect 204498 619764 204848 619798
rect 204498 619290 204554 619764
rect 204564 619290 204588 619764
rect 204618 619696 204728 619734
rect 204656 619662 204728 619696
rect 204601 619612 204657 619623
rect 204689 619612 204745 619623
rect 204612 619436 204657 619612
rect 204700 619436 204745 619612
rect 204618 619386 204728 619424
rect 204656 619352 204728 619386
rect 204498 619284 204532 619290
rect 204814 619284 204848 619764
rect 204498 619250 204848 619284
rect 205140 619132 205176 619218
rect 204530 618944 204554 619072
rect 204564 618944 204588 619072
rect 202382 617012 203835 617048
rect 203862 617012 203896 617046
rect 204520 617012 204554 617046
rect 205178 617012 205212 620460
rect 205248 620066 205250 620144
rect 205304 620010 205306 620144
rect 205248 617012 205250 617178
rect 205304 617012 205306 617234
rect 205318 617012 205352 621700
rect 205432 618660 205500 621700
rect 205540 621372 205612 621700
rect 205836 621355 205881 621700
rect 205950 621355 205984 621700
rect 206090 621664 206135 621724
rect 206748 621664 206793 621842
rect 206078 621356 206079 621357
rect 206077 621355 206078 621356
rect 205613 621344 206030 621355
rect 206090 621344 206124 621664
rect 206135 621356 206136 621357
rect 206736 621356 206737 621357
rect 206136 621355 206137 621356
rect 206735 621355 206736 621356
rect 206748 621344 206782 621664
rect 206793 621356 206794 621357
rect 207394 621356 207395 621357
rect 206794 621355 206795 621356
rect 207393 621355 207394 621356
rect 207406 621344 207440 621968
rect 207452 621956 207453 621957
rect 208051 621956 208052 621957
rect 207451 621955 207452 621956
rect 208052 621955 208053 621956
rect 207451 621356 207452 621357
rect 208052 621356 208053 621357
rect 207452 621355 207453 621356
rect 208051 621355 208052 621356
rect 208064 621344 208098 621968
rect 208110 621956 208111 621957
rect 208709 621956 208710 621957
rect 208109 621955 208110 621956
rect 208710 621955 208711 621956
rect 208109 621356 208110 621357
rect 208710 621356 208711 621357
rect 208110 621355 208111 621356
rect 208709 621355 208710 621356
rect 208722 621344 208756 621968
rect 208836 621344 208870 621968
rect 205502 621282 205612 621320
rect 205624 621310 208870 621344
rect 205540 620826 205612 621282
rect 205540 620714 205574 620826
rect 205836 620800 205881 621310
rect 205836 620686 205870 620800
rect 205950 620686 205984 621310
rect 206077 621298 206078 621299
rect 206078 621297 206079 621298
rect 206012 620770 206068 620784
rect 206012 620714 206068 620728
rect 206078 620698 206079 620699
rect 206077 620697 206078 620698
rect 206090 620686 206124 621310
rect 206136 621298 206137 621299
rect 206735 621298 206736 621299
rect 206135 621297 206136 621298
rect 206736 621297 206737 621298
rect 206135 620698 206136 620699
rect 206736 620698 206737 620699
rect 206136 620697 206137 620698
rect 206735 620697 206736 620698
rect 206748 620686 206782 621310
rect 206794 621298 206795 621299
rect 207393 621298 207394 621299
rect 206793 621297 206794 621298
rect 207394 621297 207395 621298
rect 206793 620698 206794 620699
rect 207394 620698 207395 620699
rect 206794 620697 206795 620698
rect 207393 620697 207394 620698
rect 207406 620686 207440 621310
rect 207452 621298 207453 621299
rect 208051 621298 208052 621299
rect 207451 621297 207452 621298
rect 208052 621297 208053 621298
rect 207451 620698 207452 620699
rect 208052 620698 208053 620699
rect 207452 620697 207453 620698
rect 208051 620697 208052 620698
rect 208064 620686 208098 621310
rect 208110 621298 208111 621299
rect 208709 621298 208710 621299
rect 208109 621297 208110 621298
rect 208710 621297 208711 621298
rect 208109 620698 208110 620699
rect 208710 620698 208711 620699
rect 208110 620697 208111 620698
rect 208709 620697 208710 620698
rect 208722 620686 208756 621310
rect 208836 620686 208870 621310
rect 205502 620624 205574 620662
rect 205624 620652 208870 620686
rect 205540 620056 205574 620624
rect 205836 620028 205870 620652
rect 205950 620028 205984 620652
rect 206077 620640 206078 620641
rect 206078 620639 206079 620640
rect 206078 620040 206079 620041
rect 206077 620039 206078 620040
rect 206090 620028 206124 620652
rect 206136 620640 206137 620641
rect 206735 620640 206736 620641
rect 206135 620639 206136 620640
rect 206736 620639 206737 620640
rect 206135 620040 206136 620041
rect 206736 620040 206737 620041
rect 206136 620039 206137 620040
rect 206735 620039 206736 620040
rect 206748 620028 206782 620652
rect 206794 620640 206795 620641
rect 207393 620640 207394 620641
rect 206793 620639 206794 620640
rect 207394 620639 207395 620640
rect 206793 620040 206794 620041
rect 207394 620040 207395 620041
rect 206794 620039 206795 620040
rect 207393 620039 207394 620040
rect 207406 620028 207440 620652
rect 207452 620640 207453 620641
rect 208051 620640 208052 620641
rect 207451 620639 207452 620640
rect 208052 620639 208053 620640
rect 207451 620040 207452 620041
rect 208052 620040 208053 620041
rect 207452 620039 207453 620040
rect 208051 620039 208052 620040
rect 208064 620028 208098 620652
rect 208110 620640 208111 620641
rect 208709 620640 208710 620641
rect 208109 620639 208110 620640
rect 208710 620639 208711 620640
rect 208109 620040 208110 620041
rect 208710 620040 208711 620041
rect 208110 620039 208111 620040
rect 208709 620039 208710 620040
rect 208722 620028 208756 620652
rect 208836 620028 208870 620652
rect 205502 619966 205574 620004
rect 205624 619994 208870 620028
rect 205540 619398 205574 619966
rect 205836 619370 205870 619994
rect 205950 619370 205984 619994
rect 206077 619982 206078 619983
rect 206078 619981 206079 619982
rect 206012 619448 206076 619462
rect 206012 619392 206068 619406
rect 206078 619382 206079 619383
rect 206077 619381 206078 619382
rect 206090 619370 206124 619994
rect 206136 619982 206137 619983
rect 206735 619982 206736 619983
rect 206135 619981 206136 619982
rect 206736 619981 206737 619982
rect 206135 619382 206136 619383
rect 206736 619382 206737 619383
rect 206136 619381 206137 619382
rect 206735 619381 206736 619382
rect 206748 619370 206782 619994
rect 206794 619982 206795 619983
rect 207393 619982 207394 619983
rect 206793 619981 206794 619982
rect 207394 619981 207395 619982
rect 206793 619382 206794 619383
rect 207394 619382 207395 619383
rect 206794 619381 206795 619382
rect 207393 619381 207394 619382
rect 207406 619370 207440 619994
rect 207452 619982 207453 619983
rect 208051 619982 208052 619983
rect 207451 619981 207452 619982
rect 208052 619981 208053 619982
rect 207451 619382 207452 619383
rect 208052 619382 208053 619383
rect 207452 619381 207453 619382
rect 208051 619381 208052 619382
rect 208064 619370 208098 619994
rect 208110 619982 208111 619983
rect 208709 619982 208710 619983
rect 208109 619981 208110 619982
rect 208710 619981 208711 619982
rect 208109 619382 208110 619383
rect 208710 619382 208711 619383
rect 208110 619381 208111 619382
rect 208709 619381 208710 619382
rect 208722 619370 208756 619994
rect 208836 619370 208870 619994
rect 205502 619308 205574 619346
rect 205624 619336 208870 619370
rect 205540 618740 205574 619308
rect 205836 618712 205870 619336
rect 205950 618712 205984 619336
rect 206077 619324 206078 619325
rect 206078 619323 206079 619324
rect 206012 619298 206076 619300
rect 206012 619242 206068 619244
rect 206090 618822 206124 619336
rect 206136 619324 206137 619325
rect 206735 619324 206736 619325
rect 206135 619323 206136 619324
rect 206736 619323 206737 619324
rect 206748 618822 206782 619336
rect 206794 619324 206795 619325
rect 207393 619324 207394 619325
rect 206793 619323 206794 619324
rect 207394 619323 207395 619324
rect 207406 618822 207440 619336
rect 207452 619324 207453 619325
rect 208051 619324 208052 619325
rect 207451 619323 207452 619324
rect 208052 619323 208053 619324
rect 208064 618822 208098 619336
rect 208110 619324 208111 619325
rect 208709 619324 208710 619325
rect 208109 619323 208110 619324
rect 208710 619323 208711 619324
rect 208722 618822 208756 619336
rect 206090 618725 206135 618822
rect 206748 618725 206793 618822
rect 207406 618725 207451 618822
rect 208064 618725 208109 618822
rect 206078 618724 206079 618725
rect 206090 618724 206136 618725
rect 206736 618724 206737 618725
rect 206748 618724 206794 618725
rect 207394 618724 207395 618725
rect 207406 618724 207452 618725
rect 208052 618724 208053 618725
rect 208064 618724 208110 618725
rect 208710 618724 208711 618725
rect 208722 618724 208767 618822
rect 206077 618723 206078 618724
rect 206090 618712 206124 618724
rect 206136 618723 206137 618724
rect 206735 618723 206736 618724
rect 206136 618712 206736 618723
rect 206748 618712 206782 618724
rect 206794 618723 206795 618724
rect 207393 618723 207394 618724
rect 206794 618712 207394 618723
rect 207406 618712 207440 618724
rect 207452 618723 207453 618724
rect 208051 618723 208052 618724
rect 207452 618712 208052 618723
rect 208064 618712 208098 618724
rect 208110 618723 208111 618724
rect 208709 618723 208710 618724
rect 208110 618712 208710 618723
rect 208722 618712 208756 618724
rect 208836 618712 208870 619336
rect 208967 620052 212591 622082
rect 213200 620652 213616 620674
rect 213234 620618 213650 620640
rect 208967 619960 212642 620052
rect 208967 619952 212591 619960
rect 208967 619940 212614 619952
rect 208967 619934 212842 619940
rect 208967 619932 213018 619934
rect 208967 618712 212591 619932
rect 212614 619906 212814 619912
rect 212614 619904 213046 619906
rect 213196 619848 213658 620486
rect 213254 619764 213604 619798
rect 213254 619284 213288 619764
rect 213446 619696 213484 619734
rect 213412 619662 213484 619696
rect 213357 619612 213402 619623
rect 213445 619612 213490 619623
rect 213368 619436 213402 619612
rect 213456 619436 213490 619612
rect 213446 619404 213484 619424
rect 213412 619382 213484 619404
rect 213396 619370 213484 619382
rect 213396 619336 213462 619370
rect 213570 619284 213604 619764
rect 213254 619250 213604 619284
rect 205624 618678 212591 618712
rect 205432 618598 205477 618660
rect 205836 618598 205870 618678
rect 205950 618598 205984 618678
rect 206090 618598 206124 618678
rect 206748 618598 206782 618678
rect 207406 618598 207440 618678
rect 208064 618598 208098 618678
rect 208722 618598 208756 618678
rect 208836 618598 208870 618678
rect 208967 618598 212591 618678
rect 205432 618564 212591 618598
rect 205432 618550 205477 618564
rect 205432 618510 205466 618550
rect 205432 618454 205477 618510
rect 205432 618368 205548 618454
rect 205432 618229 205477 618368
rect 205836 618229 205870 618564
rect 205950 618229 205984 618564
rect 206054 618292 206068 618492
rect 206752 618352 206782 618514
rect 206790 618390 206820 618476
rect 205998 618236 206012 618292
rect 208722 618229 208756 618564
rect 208836 618229 208870 618564
rect 208967 618528 212591 618564
rect 205397 618193 208906 618229
rect 209003 618193 209037 618528
rect 209117 618193 209151 618528
rect 209775 618193 209809 618227
rect 210433 618193 210467 618227
rect 211057 618193 211060 618288
rect 211085 618193 211088 618288
rect 211091 618193 211125 618227
rect 211749 618193 211783 618227
rect 212407 618193 212441 618227
rect 212521 618193 212555 618528
rect 205397 618159 213703 618193
rect 205397 617012 208906 618159
rect 202382 617007 208906 617012
rect 209003 618079 209037 618159
rect 209117 618079 209151 618159
rect 209163 618079 209763 618090
rect 209775 618079 209809 618159
rect 210433 618079 210467 618159
rect 211057 618085 211060 618159
rect 211085 618085 211088 618159
rect 211091 618079 211125 618159
rect 211749 618079 211783 618159
rect 212407 618079 212441 618159
rect 212521 618079 212555 618159
rect 209003 618045 212555 618079
rect 209003 617421 209037 618045
rect 209117 618033 209151 618045
rect 209163 618033 209164 618034
rect 209762 618033 209763 618034
rect 209775 618033 209809 618045
rect 209821 618033 209822 618034
rect 210420 618033 210421 618034
rect 209117 618032 209163 618033
rect 209763 618032 209764 618033
rect 209775 618032 209821 618033
rect 210421 618032 210422 618033
rect 209117 617434 209162 618032
rect 209775 617434 209820 618032
rect 209117 617433 209163 617434
rect 209763 617433 209764 617434
rect 209775 617433 209821 617434
rect 210421 617433 210422 617434
rect 209117 617421 209151 617433
rect 209163 617432 209164 617433
rect 209762 617432 209763 617433
rect 209163 617421 209763 617432
rect 209775 617421 209809 617433
rect 209821 617432 209822 617433
rect 210420 617432 210421 617433
rect 209821 617421 209858 617432
rect 210433 617421 210467 618045
rect 210479 618033 210480 618034
rect 210478 618032 210479 618033
rect 211057 617962 211060 618039
rect 211078 618033 211079 618034
rect 211079 618032 211080 618033
rect 211085 617962 211088 618039
rect 210478 617433 210479 617434
rect 210479 617432 210480 617433
rect 211057 617427 211060 617514
rect 211079 617433 211080 617434
rect 211078 617432 211079 617433
rect 211085 617427 211088 617514
rect 211091 617421 211125 618045
rect 211137 618033 211138 618034
rect 211736 618033 211737 618034
rect 211136 618032 211137 618033
rect 211737 618032 211738 618033
rect 211684 617514 211743 617524
rect 211712 617486 211743 617496
rect 211136 617433 211137 617434
rect 211737 617433 211738 617434
rect 211137 617432 211138 617433
rect 211736 617432 211737 617433
rect 211749 617421 211783 618045
rect 211795 618033 211796 618034
rect 212394 618033 212395 618034
rect 211794 618032 211795 618033
rect 212395 618032 212396 618033
rect 211789 617514 211848 617524
rect 211789 617486 211820 617496
rect 211794 617433 211795 617434
rect 212395 617433 212396 617434
rect 211795 617432 211796 617433
rect 212394 617432 212395 617433
rect 212407 617421 212441 618045
rect 212521 617421 212555 618045
rect 209003 617387 212555 617421
rect 209003 617007 209037 617387
rect 209117 617375 209151 617387
rect 209163 617375 209164 617376
rect 209762 617375 209763 617376
rect 209775 617375 209809 617387
rect 209821 617375 209822 617376
rect 210420 617375 210421 617376
rect 209117 617374 209163 617375
rect 209763 617374 209764 617375
rect 209775 617374 209821 617375
rect 210421 617374 210422 617375
rect 209117 617007 209162 617374
rect 202382 616978 209655 617007
rect 202382 616948 203835 616978
rect 202382 616876 203858 616948
rect 203862 616926 203896 616978
rect 201615 615736 201661 615751
rect 201648 615705 201661 615736
rect 202382 615643 203835 616876
rect 203862 616838 203908 616926
rect 204478 616910 204516 616948
rect 203910 616876 204516 616910
rect 204520 616926 204554 616978
rect 204520 616838 204566 616926
rect 205136 616910 205174 616948
rect 204568 616876 205174 616910
rect 205178 616926 205212 616978
rect 205178 616838 205224 616926
rect 205234 616916 205250 616978
rect 205304 616942 205306 616978
rect 205290 616916 205306 616942
rect 205318 616910 205352 616978
rect 205397 616974 209655 616978
rect 205397 616973 209680 616974
rect 205397 616910 208906 616973
rect 205226 616876 208906 616910
rect 209003 616905 209037 616973
rect 209117 616952 209162 616973
rect 209117 616905 209164 616952
rect 209290 616940 209680 616973
rect 209290 616905 209324 616940
rect 209479 616919 209526 616940
rect 209479 616905 209551 616919
rect 203837 616826 203850 616837
rect 203862 616826 203896 616838
rect 204495 616826 204508 616837
rect 204520 616826 204554 616838
rect 205153 616826 205166 616837
rect 205178 616826 205212 616838
rect 200247 615609 203835 615643
rect 200093 615496 200127 615508
rect 198841 615449 198845 615455
rect 199421 615449 199469 615455
rect 200079 615449 200127 615496
rect 200680 615455 200682 615609
rect 200708 615496 200738 615609
rect 200751 615508 200799 615609
rect 200751 615496 200785 615508
rect 200708 615455 200785 615496
rect 200737 615449 200785 615455
rect 198837 615415 198845 615449
rect 198853 615415 199469 615449
rect 199495 615415 199503 615449
rect 199511 615415 200127 615449
rect 200153 615415 200161 615449
rect 200169 615415 200785 615449
rect 198841 615409 198845 615415
rect 199423 615409 199469 615415
rect 199358 615402 199360 615409
rect 199386 615374 199388 615409
rect 199423 615399 199514 615409
rect 199435 615347 199514 615399
rect 199524 615347 199542 615409
rect 200081 615399 200127 615415
rect 200680 615402 200682 615409
rect 200093 615347 200127 615399
rect 200708 615347 200738 615409
rect 200739 615399 200785 615415
rect 200751 615347 200785 615399
rect 200865 615409 200913 615609
rect 202382 615573 203835 615609
rect 202418 615432 202466 615573
rect 202532 615522 202580 615573
rect 197449 615313 200797 615347
rect 197492 615180 197501 615313
rect 197520 615208 197529 615313
rect 199468 615172 199514 615313
rect 199468 614968 199475 615172
rect 199524 615144 199542 615313
rect 200708 615264 200724 615313
rect 179580 610435 179661 610472
rect 179708 610457 187381 610487
rect 179704 610453 187381 610457
rect 187399 610453 187501 610487
rect 179708 610447 185632 610453
rect 186388 610444 186864 610453
rect 179580 610429 179708 610435
rect 185984 610432 186864 610444
rect 187284 610441 187381 610453
rect 179580 610423 185632 610429
rect 185984 610423 186440 610432
rect 187272 610423 187283 610434
rect 179580 610419 187288 610423
rect 179580 610392 187283 610419
rect 187284 610392 187365 610408
rect 179580 610389 187365 610392
rect 179586 610383 185632 610389
rect 179611 610377 179708 610383
rect 179614 610355 179621 610364
rect 179627 609891 179661 610377
rect 185984 610374 186440 610389
rect 186984 610383 187365 610389
rect 187284 610373 187365 610383
rect 187284 610364 187371 610373
rect 187433 610364 187467 610453
rect 179667 610355 185632 610364
rect 186984 610348 187467 610364
rect 199468 610360 199475 613780
rect 200865 610698 200899 615409
rect 202418 610748 202452 615432
rect 202532 615370 202566 615522
rect 202636 615478 202652 615573
rect 202664 615478 202680 615573
rect 203118 615478 203126 615573
rect 203146 615478 203154 615573
rect 203190 615522 203238 615573
rect 203848 615522 203896 616826
rect 204506 615522 204554 616826
rect 205164 615522 205212 616826
rect 205234 615776 205250 616870
rect 205290 615734 205306 616870
rect 205318 615666 205352 616876
rect 205397 616852 208906 616876
rect 208911 616871 209551 616905
rect 205397 616769 208917 616852
rect 205397 616763 208906 616769
rect 209003 616763 209037 616871
rect 209117 616763 209151 616871
rect 209290 616763 209324 616871
rect 209466 616838 209551 616871
rect 209507 616823 209541 616828
rect 209496 616812 209541 616823
rect 209507 616795 209541 616812
rect 209507 616790 209552 616795
rect 209393 616779 209438 616790
rect 209404 616763 209438 616779
rect 209507 616763 209566 616790
rect 209621 616763 209680 616940
rect 209775 616970 209820 617374
rect 209763 616775 209764 616776
rect 209762 616774 209763 616775
rect 209775 616763 209809 616970
rect 209820 616775 209821 616776
rect 210421 616775 210422 616776
rect 209821 616774 209822 616775
rect 210420 616774 210421 616775
rect 210433 616763 210467 617387
rect 210479 617375 210480 617376
rect 210478 617374 210479 617375
rect 211057 617304 211060 617381
rect 211078 617375 211079 617376
rect 211079 617374 211080 617375
rect 211085 617304 211088 617381
rect 210478 616775 210479 616776
rect 210479 616774 210480 616775
rect 211057 616769 211060 616856
rect 211079 616775 211080 616776
rect 211078 616774 211079 616775
rect 211085 616769 211088 616856
rect 211091 616763 211125 617387
rect 211137 617375 211138 617376
rect 211736 617375 211737 617376
rect 211136 617374 211137 617375
rect 211737 617374 211738 617375
rect 211749 617048 211783 617387
rect 211795 617375 211796 617376
rect 212394 617375 212395 617376
rect 211794 617374 211795 617375
rect 212395 617374 212396 617375
rect 212324 617336 212401 617360
rect 212407 617048 212441 617387
rect 212521 617360 212555 617387
rect 212447 617336 212576 617360
rect 212521 617048 212555 617336
rect 211138 617012 213835 617048
rect 214074 617012 214108 623884
rect 216294 623268 216310 623838
rect 214916 622368 214938 623230
rect 214916 622126 214938 622230
rect 216294 622052 216314 623268
rect 216294 618276 216310 622052
rect 214188 617012 214222 617046
rect 211138 616978 214726 617012
rect 211136 616775 211137 616776
rect 211138 616775 213835 616978
rect 213942 616842 213962 616944
rect 213970 616870 213990 616916
rect 211137 616774 213835 616775
rect 211138 616763 213835 616774
rect 205397 616729 213835 616763
rect 205397 616723 208906 616729
rect 205397 616642 208917 616723
rect 205397 616200 208906 616642
rect 205397 616194 208976 616200
rect 205397 616105 208906 616194
rect 208922 616138 208976 616144
rect 209003 616105 209037 616729
rect 209117 616105 209151 616729
rect 209290 616442 209324 616729
rect 209404 616603 209438 616729
rect 209507 616603 209566 616729
rect 209507 616591 209552 616603
rect 209504 616587 209552 616591
rect 209504 616544 209551 616587
rect 209466 616538 209551 616544
rect 209621 616538 209680 616729
rect 209762 616717 209763 616718
rect 209763 616716 209764 616717
rect 209775 616538 209809 616729
rect 209821 616717 209822 616718
rect 210420 616717 210421 616718
rect 209820 616716 209821 616717
rect 210421 616716 210422 616717
rect 209358 616442 209809 616538
rect 209290 616408 209809 616442
rect 209358 616358 209809 616408
rect 209272 616326 209809 616358
rect 209272 616105 209694 616326
rect 209763 616117 209764 616118
rect 209762 616116 209763 616117
rect 209775 616105 209809 616326
rect 209820 616117 209821 616118
rect 209821 616116 209822 616117
rect 209892 616111 209894 616194
rect 210392 616116 210427 616139
rect 210364 616105 210427 616111
rect 210433 616105 210467 616729
rect 210479 616717 210480 616718
rect 210478 616716 210479 616717
rect 211057 616642 211060 616723
rect 211078 616717 211079 616718
rect 211079 616716 211080 616717
rect 211085 616642 211088 616723
rect 210473 616116 210500 616139
rect 211057 616111 211060 616194
rect 211079 616117 211080 616118
rect 211078 616116 211079 616117
rect 211085 616111 211088 616194
rect 210473 616105 210528 616111
rect 211091 616105 211125 616729
rect 211138 616718 213835 616729
rect 211137 616717 213835 616718
rect 211136 616716 211137 616717
rect 211136 616117 211137 616118
rect 211138 616117 213835 616717
rect 211137 616116 213835 616117
rect 211138 616105 213835 616116
rect 205397 616071 213835 616105
rect 205397 615666 208906 616071
rect 205318 615632 208906 615666
rect 205397 615596 208906 615632
rect 209003 615643 209037 616071
rect 209117 615814 209151 616071
rect 209272 615842 209694 616071
rect 209762 616059 209763 616060
rect 209763 616058 209764 616059
rect 209775 615842 209809 616071
rect 209821 616059 209822 616060
rect 209820 616058 209821 616059
rect 209892 615972 209894 616065
rect 210420 616059 210421 616060
rect 210421 616058 210422 616059
rect 209117 615804 209162 615814
rect 209272 615804 209809 615842
rect 210433 615804 210467 616071
rect 210479 616059 210480 616060
rect 210478 616058 210479 616059
rect 211057 615972 211060 616065
rect 211078 616059 211079 616060
rect 211079 616058 211080 616059
rect 211085 615972 211088 616065
rect 211091 615804 211125 616071
rect 211138 616060 213835 616071
rect 211137 616059 213835 616060
rect 211136 616058 211137 616059
rect 209272 615792 209798 615804
rect 209132 615745 209798 615792
rect 210405 615745 210452 615792
rect 211063 615745 211110 615792
rect 209179 615711 209798 615745
rect 209837 615711 210452 615745
rect 210495 615711 211110 615745
rect 209350 615643 209798 615711
rect 211138 615643 213835 616059
rect 209003 615609 213835 615643
rect 214074 615666 214108 616978
rect 214176 616876 214588 616948
rect 214176 616838 214234 616876
rect 214188 615818 214233 616838
rect 214567 616826 214623 616837
rect 214578 615806 214623 616826
rect 214212 615768 214624 615806
rect 214250 615734 214624 615768
rect 214566 615718 214624 615734
rect 214609 615703 214624 615718
rect 214692 615666 214726 616978
rect 216266 615774 216268 618220
rect 216294 615774 216324 618276
rect 215110 615734 215476 615756
rect 215148 615666 215520 615718
rect 216266 615682 216268 615728
rect 216294 615710 216324 615728
rect 214074 615632 217530 615666
rect 203190 615510 203224 615522
rect 203848 615510 203882 615522
rect 204506 615510 204540 615522
rect 205164 615510 205198 615522
rect 205397 615510 206020 615596
rect 203176 615472 203224 615510
rect 203834 615472 203888 615510
rect 202592 615438 202600 615472
rect 202608 615438 203224 615472
rect 203250 615438 203258 615472
rect 203266 615438 203888 615472
rect 202636 615370 202652 615432
rect 202664 615370 202680 615432
rect 203118 615426 203126 615432
rect 203146 615398 203154 615432
rect 203178 615422 203224 615438
rect 203836 615422 203888 615438
rect 203190 615370 203224 615422
rect 203844 615370 203888 615422
rect 203900 615370 203916 615510
rect 204492 615472 204540 615510
rect 205150 615472 205198 615510
rect 203924 615438 204540 615472
rect 204566 615438 204574 615472
rect 204582 615438 205198 615472
rect 204494 615422 204540 615438
rect 205152 615422 205198 615438
rect 204506 615370 204540 615422
rect 205164 615370 205198 615422
rect 205200 615404 205206 615506
rect 205316 615484 206020 615510
rect 205228 615472 205274 615478
rect 205316 615472 206036 615484
rect 205224 615468 206036 615472
rect 205224 615447 206020 615468
rect 206103 615447 206137 615596
rect 206217 615484 206262 615596
rect 206386 615484 206808 615596
rect 206217 615468 206334 615484
rect 206386 615468 206832 615484
rect 206217 615460 206262 615468
rect 206217 615459 206263 615460
rect 206217 615447 206251 615459
rect 206263 615458 206264 615459
rect 206386 615458 206808 615468
rect 206875 615460 206920 615596
rect 206960 615468 206992 615484
rect 207533 615460 207578 615596
rect 208191 615460 208236 615596
rect 208849 615460 208894 615596
rect 209492 615502 209562 615609
rect 206863 615459 206864 615460
rect 206875 615459 206921 615460
rect 207521 615459 207522 615460
rect 207533 615459 207579 615460
rect 208179 615459 208180 615460
rect 208191 615459 208237 615460
rect 208837 615459 208838 615460
rect 208849 615459 208895 615460
rect 209495 615459 209496 615460
rect 206862 615458 206863 615459
rect 206263 615447 206863 615458
rect 206875 615447 206909 615459
rect 206921 615458 206922 615459
rect 207520 615458 207521 615459
rect 206921 615447 207521 615458
rect 207533 615447 207567 615459
rect 207579 615458 207580 615459
rect 208178 615458 208179 615459
rect 207579 615447 208179 615458
rect 208191 615447 208225 615459
rect 208237 615458 208238 615459
rect 208836 615458 208837 615459
rect 208237 615447 208837 615458
rect 208849 615447 208883 615459
rect 208895 615458 208896 615459
rect 209494 615458 209495 615459
rect 209507 615447 209541 615502
rect 209621 615447 209655 615609
rect 205224 615438 209655 615447
rect 205228 615432 205262 615438
rect 205397 615413 209655 615438
rect 205397 615370 206020 615413
rect 202520 615336 206020 615370
rect 202636 615264 202652 615336
rect 202664 615264 202680 615336
rect 202636 612882 202652 613780
rect 202664 612882 202680 613780
rect 202636 612482 202652 612682
rect 202664 612482 202680 612682
rect 202636 611130 202652 612282
rect 202664 611102 202680 612282
rect 186984 610327 187365 610348
rect 183450 610160 183898 610232
rect 183018 610020 183898 610160
rect 183018 609948 183466 610020
rect 179627 609858 180032 609891
rect 179525 609842 180032 609858
rect 179284 609725 179299 609771
rect 150584 608710 150962 609414
rect 179284 609073 179299 609113
rect 179525 608993 179559 609842
rect 179708 609829 180032 609835
rect 180436 609829 181090 609848
rect 181434 609842 187325 609863
rect 187331 609842 187365 610327
rect 187371 609842 187384 609863
rect 187284 609841 187365 609842
rect 187284 609835 187381 609841
rect 181434 609829 187412 609835
rect 187433 609829 187467 610348
rect 179708 609814 187501 609829
rect 179580 609777 179661 609814
rect 179720 609799 187381 609814
rect 179704 609795 187381 609799
rect 187399 609795 187501 609814
rect 180436 609786 181090 609795
rect 181434 609789 187381 609795
rect 179580 609765 179708 609777
rect 179992 609774 181090 609786
rect 187284 609783 187381 609789
rect 179992 609765 180646 609774
rect 187272 609771 187283 609776
rect 181434 609765 187284 609771
rect 179580 609761 187288 609765
rect 179580 609758 187283 609761
rect 179580 609750 187284 609758
rect 179580 609731 187365 609750
rect 179611 609719 179708 609731
rect 179627 609199 179661 609719
rect 179992 609712 180646 609731
rect 185994 609730 187365 609731
rect 180988 609725 187365 609730
rect 187284 609703 187365 609725
rect 180988 609697 187312 609702
rect 180988 609669 181490 609697
rect 183442 609514 183890 609586
rect 183018 609374 183890 609514
rect 183018 609302 183466 609374
rect 179680 609190 180262 609205
rect 180462 609190 186050 609205
rect 187331 609184 187365 609703
rect 187284 609183 187365 609184
rect 179708 609171 180262 609177
rect 180462 609171 186050 609177
rect 187284 609171 187381 609183
rect 187433 609171 187467 609795
rect 197522 609172 197536 610360
rect 179580 609119 179661 609156
rect 179708 609141 187381 609171
rect 179704 609137 187381 609141
rect 187399 609137 187501 609171
rect 179708 609131 180270 609137
rect 179580 609113 179708 609119
rect 180262 609118 180270 609131
rect 180456 609131 185602 609137
rect 180456 609118 180462 609131
rect 186424 609120 186430 609134
rect 187284 609125 187381 609137
rect 179580 609107 180270 609113
rect 180456 609107 185602 609113
rect 187272 609107 187283 609118
rect 179580 609103 187288 609107
rect 179580 609073 187283 609103
rect 179596 609072 179708 609073
rect 179586 609067 180270 609072
rect 180456 609067 185602 609072
rect 186954 609067 187284 609072
rect 179596 609061 179708 609067
rect 187433 609044 187467 609137
rect 179614 609039 179621 609044
rect 179667 609039 180270 609044
rect 180456 609039 185602 609044
rect 186954 609038 187467 609044
rect 186954 609011 187340 609038
rect 187433 608993 187467 609038
rect 179197 608959 187467 608993
rect 150928 608400 150962 608710
rect 179525 608461 179559 608959
rect 199468 608839 199475 609172
rect 199435 608836 199475 608839
rect 200751 608836 200785 610698
rect 202290 610430 202306 610604
rect 202318 610456 202334 610576
rect 202382 610450 202498 610748
rect 202548 610656 203096 610690
rect 202548 610628 202582 610656
rect 202514 610594 202582 610628
rect 202316 610446 202498 610450
rect 202382 610286 202498 610446
rect 202548 610436 202600 610594
rect 202910 610576 202921 610587
rect 202612 610532 202684 610570
rect 202734 610542 202921 610576
rect 202922 610532 202994 610570
rect 202650 610498 202684 610532
rect 202910 610488 202921 610499
rect 202960 610498 202994 610532
rect 202734 610454 202921 610488
rect 202548 610374 202582 610436
rect 203062 610374 203096 610656
rect 202548 610340 203096 610374
rect 202516 610148 202590 610222
rect 202464 610076 202590 610148
rect 203190 610098 203224 615336
rect 203844 615264 203888 615336
rect 203900 615264 203916 615336
rect 205397 615300 206020 615336
rect 205397 614789 206006 615300
rect 206103 614827 206137 615413
rect 206179 615360 206180 615413
rect 206217 615401 206251 615413
rect 206263 615401 206264 615402
rect 206862 615401 206863 615402
rect 206875 615401 206909 615413
rect 206921 615401 206922 615402
rect 207520 615401 207521 615402
rect 207533 615401 207567 615413
rect 207579 615401 207580 615402
rect 208178 615401 208179 615402
rect 208191 615401 208225 615413
rect 208237 615401 208238 615402
rect 208836 615401 208837 615402
rect 208849 615401 208883 615413
rect 208895 615401 208896 615402
rect 209494 615401 209495 615402
rect 206217 615400 206263 615401
rect 206863 615400 206864 615401
rect 206875 615400 206921 615401
rect 207521 615400 207522 615401
rect 207533 615400 207579 615401
rect 208179 615400 208180 615401
rect 208191 615400 208237 615401
rect 208837 615400 208838 615401
rect 208849 615400 208895 615401
rect 209495 615400 209496 615401
rect 206217 614827 206262 615400
rect 206022 614822 206464 614827
rect 206103 614789 206137 614822
rect 206217 614802 206262 614822
rect 206875 614802 206920 615400
rect 207533 614802 207578 615400
rect 208191 614802 208236 615400
rect 208772 614826 208794 614851
rect 208849 614802 208894 615400
rect 206217 614801 206263 614802
rect 206863 614801 206864 614802
rect 206875 614801 206921 614802
rect 207521 614801 207522 614802
rect 207533 614801 207579 614802
rect 208179 614801 208180 614802
rect 208191 614801 208237 614802
rect 208837 614801 208838 614802
rect 208849 614801 208895 614802
rect 206217 614789 206251 614801
rect 206263 614800 206264 614801
rect 206862 614800 206863 614801
rect 206263 614789 206863 614800
rect 206875 614789 206909 614801
rect 206921 614800 206922 614801
rect 207520 614800 207521 614801
rect 206921 614789 207521 614800
rect 207533 614789 207567 614801
rect 207579 614800 207580 614801
rect 208178 614800 208179 614801
rect 207579 614789 208179 614800
rect 208191 614789 208225 614801
rect 208237 614800 208238 614801
rect 208836 614800 208837 614801
rect 208237 614789 208837 614800
rect 208849 614795 208889 614801
rect 208895 614800 208896 614801
rect 208849 614789 208883 614795
rect 208895 614789 208898 614800
rect 208906 614795 208917 614872
rect 209495 614801 209496 614802
rect 209494 614800 209495 614801
rect 209507 614789 209541 615413
rect 209621 614789 209655 615413
rect 205397 614784 209655 614789
rect 205397 614675 206006 614784
rect 206103 614755 209655 614784
rect 206103 614675 206137 614755
rect 206217 614675 206251 614755
rect 206875 614675 206909 614755
rect 207533 614675 207567 614755
rect 208191 614675 208225 614755
rect 208772 614749 208883 614755
rect 208843 614675 208889 614749
rect 208906 614675 208917 614749
rect 209507 614675 209541 614755
rect 209621 614675 209655 614755
rect 211138 614675 213835 615609
rect 205397 614641 213835 614675
rect 205397 614605 206006 614641
rect 203750 610360 203764 610598
rect 203844 610542 203888 613780
rect 203900 610542 203916 613780
rect 205822 613122 205856 613156
rect 205936 613122 205970 614605
rect 205998 614570 206046 614578
rect 205998 614536 206012 614544
rect 206103 613158 206137 614641
rect 208843 614020 208889 614641
rect 208906 614076 208917 614641
rect 208862 613442 208883 613980
rect 209621 613978 209655 614641
rect 211138 614605 213835 614641
rect 208862 613372 208889 613442
rect 208862 613234 208883 613372
rect 208862 613178 208889 613234
rect 208896 613206 208917 613946
rect 209038 613556 209658 613978
rect 209708 613574 209709 613964
rect 210042 613538 210310 613772
rect 209520 613198 209547 613454
rect 209548 613226 209575 613426
rect 210458 613312 210464 613414
rect 210492 613346 210498 613380
rect 208862 613174 208883 613178
rect 206067 613122 209691 613158
rect 205456 613088 209691 613122
rect 205128 610360 205144 610506
rect 205234 610360 205236 610382
rect 201628 609772 201782 609876
rect 201520 609472 202016 609772
rect 202516 609568 202590 610076
rect 203128 610012 203224 610098
rect 200834 609268 202476 609288
rect 200834 609212 202476 609232
rect 203190 608850 203224 610012
rect 204532 609934 204540 609984
rect 204522 609508 204540 609934
rect 204566 609900 204574 609950
rect 204556 609542 204574 609900
rect 205456 609604 205490 613088
rect 205822 613008 205856 613088
rect 205936 613008 205970 613088
rect 205520 612946 205592 612984
rect 205642 612974 205970 613008
rect 205809 612962 205810 612963
rect 205810 612961 205811 612962
rect 205558 612378 205592 612946
rect 205810 612362 205811 612363
rect 205809 612361 205810 612362
rect 205822 612350 205856 612974
rect 205936 612350 205970 612974
rect 205520 612288 205592 612326
rect 205642 612316 205970 612350
rect 205809 612304 205810 612305
rect 205810 612303 205811 612304
rect 205558 611720 205592 612288
rect 205810 611704 205811 611705
rect 205809 611703 205810 611704
rect 205822 611692 205856 612316
rect 205936 611692 205970 612316
rect 205520 611630 205592 611668
rect 205642 611658 205970 611692
rect 205809 611646 205810 611647
rect 205810 611645 205811 611646
rect 205558 611062 205592 611630
rect 205810 611046 205811 611047
rect 205809 611045 205810 611046
rect 205822 611034 205856 611658
rect 205936 611034 205970 611658
rect 205520 610972 205592 611010
rect 205642 611000 205970 611034
rect 205809 610988 205810 610989
rect 205810 610987 205811 610988
rect 205558 610404 205592 610972
rect 205822 610468 205856 611000
rect 205936 610468 205970 611000
rect 206067 612972 209691 613088
rect 210296 613122 210758 613158
rect 211174 613122 211208 614605
rect 211288 613122 211322 613156
rect 211946 613122 211980 613156
rect 212604 613122 212638 613156
rect 213262 613122 213296 613156
rect 210296 613088 213804 613122
rect 206067 612968 209942 612972
rect 206067 610468 209691 612968
rect 209714 612940 209914 612944
rect 210296 612880 210758 613088
rect 211174 613008 211208 613088
rect 211288 613008 211322 613088
rect 211946 613008 211980 613088
rect 212604 613008 212638 613088
rect 213262 613008 213296 613088
rect 213618 613008 213629 613019
rect 210842 612968 211098 612984
rect 211174 612974 213629 613008
rect 210870 612940 211070 612956
rect 210354 612796 210704 612830
rect 210354 612316 210388 612796
rect 210546 612728 210584 612766
rect 210512 612694 210584 612728
rect 210457 612644 210502 612655
rect 210545 612644 210590 612655
rect 210468 612468 210502 612644
rect 210556 612468 210590 612644
rect 210546 612454 210584 612456
rect 210468 612428 210590 612454
rect 210546 612426 210584 612428
rect 210496 612400 210584 612426
rect 210512 612384 210584 612400
rect 210496 612368 210562 612384
rect 210468 612340 210590 612356
rect 210608 612316 210642 612350
rect 210670 612316 210704 612796
rect 210354 612282 210704 612316
rect 211174 612350 211208 612974
rect 211288 612350 211322 612974
rect 211334 612962 211335 612963
rect 211933 612962 211934 612963
rect 211333 612961 211334 612962
rect 211934 612961 211935 612962
rect 211333 612362 211334 612363
rect 211934 612362 211935 612363
rect 211334 612361 211335 612362
rect 211933 612361 211934 612362
rect 211946 612350 211980 612974
rect 211992 612962 211993 612963
rect 212591 612962 212592 612963
rect 211991 612961 211992 612962
rect 212592 612961 212593 612962
rect 211991 612362 211992 612363
rect 212592 612362 212593 612363
rect 211992 612361 211993 612362
rect 212591 612361 212592 612362
rect 212604 612350 212638 612974
rect 212650 612962 212651 612963
rect 213249 612962 213250 612963
rect 212649 612961 212650 612962
rect 213250 612961 213251 612962
rect 212649 612362 212650 612363
rect 213250 612362 213251 612363
rect 212650 612361 212651 612362
rect 213249 612361 213250 612362
rect 213262 612350 213296 612974
rect 213308 612962 213309 612963
rect 213307 612961 213308 612962
rect 213630 612946 213702 612984
rect 213668 612378 213702 612946
rect 213307 612362 213308 612363
rect 213308 612361 213309 612362
rect 213618 612350 213629 612361
rect 211174 612316 213629 612350
rect 205822 610454 209691 610468
rect 205810 610388 205811 610389
rect 205809 610387 205810 610388
rect 205822 610382 205862 610454
rect 205822 610376 205856 610382
rect 205936 610376 205970 610454
rect 205520 610314 205592 610352
rect 205642 610342 205970 610376
rect 205809 610330 205810 610331
rect 205810 610329 205811 610330
rect 205558 609746 205592 610314
rect 205810 609730 205811 609731
rect 205809 609729 205810 609730
rect 205822 609718 205856 610342
rect 205936 609718 205970 610342
rect 205642 609684 205970 609718
rect 205822 609604 205856 609684
rect 205936 609604 205970 609684
rect 206067 609604 209691 610454
rect 211174 611692 211208 612316
rect 211288 611692 211322 612316
rect 211334 612304 211335 612305
rect 211933 612304 211934 612305
rect 211333 612303 211334 612304
rect 211934 612303 211935 612304
rect 211333 611704 211334 611705
rect 211934 611704 211935 611705
rect 211334 611703 211335 611704
rect 211933 611703 211934 611704
rect 211946 611692 211980 612316
rect 211992 612304 211993 612305
rect 212591 612304 212592 612305
rect 211991 612303 211992 612304
rect 212592 612303 212593 612304
rect 211991 611704 211992 611705
rect 212592 611704 212593 611705
rect 211992 611703 211993 611704
rect 212591 611703 212592 611704
rect 212604 611692 212638 612316
rect 212650 612304 212651 612305
rect 213249 612304 213250 612305
rect 212649 612303 212650 612304
rect 213250 612303 213251 612304
rect 212649 611704 212650 611705
rect 213250 611704 213251 611705
rect 212650 611703 212651 611704
rect 213249 611703 213250 611704
rect 213262 611692 213296 612316
rect 213308 612304 213309 612305
rect 213307 612303 213308 612304
rect 213630 612288 213702 612326
rect 213668 611720 213702 612288
rect 213307 611704 213308 611705
rect 213308 611703 213309 611704
rect 213618 611692 213629 611703
rect 211174 611658 213629 611692
rect 211174 611034 211208 611658
rect 211288 611034 211322 611658
rect 211334 611646 211335 611647
rect 211933 611646 211934 611647
rect 211333 611645 211334 611646
rect 211934 611645 211935 611646
rect 211333 611046 211334 611047
rect 211934 611046 211935 611047
rect 211334 611045 211335 611046
rect 211933 611045 211934 611046
rect 211946 611034 211980 611658
rect 211992 611646 211993 611647
rect 212591 611646 212592 611647
rect 211991 611645 211992 611646
rect 212592 611645 212593 611646
rect 211991 611046 211992 611047
rect 212592 611046 212593 611047
rect 211992 611045 211993 611046
rect 212591 611045 212592 611046
rect 212604 611034 212638 611658
rect 212650 611646 212651 611647
rect 213249 611646 213250 611647
rect 212649 611645 212650 611646
rect 213250 611645 213251 611646
rect 212649 611046 212650 611047
rect 213250 611046 213251 611047
rect 212650 611045 212651 611046
rect 213249 611045 213250 611046
rect 213262 611034 213296 611658
rect 213308 611646 213309 611647
rect 213307 611645 213308 611646
rect 213630 611630 213702 611668
rect 213668 611062 213702 611630
rect 213307 611046 213308 611047
rect 213308 611045 213309 611046
rect 213618 611034 213629 611045
rect 211174 611000 213629 611034
rect 211174 610376 211208 611000
rect 211288 610376 211322 611000
rect 211334 610988 211335 610989
rect 211933 610988 211934 610989
rect 211333 610987 211334 610988
rect 211934 610987 211935 610988
rect 211333 610388 211334 610389
rect 211934 610388 211935 610389
rect 211334 610387 211335 610388
rect 211933 610387 211934 610388
rect 211946 610376 211980 611000
rect 211992 610988 211993 610989
rect 212591 610988 212592 610989
rect 211991 610987 211992 610988
rect 212592 610987 212593 610988
rect 211991 610388 211992 610389
rect 212592 610388 212593 610389
rect 211992 610387 211993 610388
rect 212591 610387 212592 610388
rect 212604 610376 212638 611000
rect 212650 610988 212651 610989
rect 213249 610988 213250 610989
rect 212649 610987 212650 610988
rect 213250 610987 213251 610988
rect 212649 610388 212650 610389
rect 213250 610388 213251 610389
rect 212650 610387 212651 610388
rect 213249 610387 213250 610388
rect 213262 610376 213296 611000
rect 213308 610988 213309 610989
rect 213307 610987 213308 610988
rect 213630 610972 213702 611010
rect 213668 610404 213702 610972
rect 213307 610388 213308 610389
rect 213308 610387 213309 610388
rect 213618 610376 213629 610387
rect 211174 610342 213629 610376
rect 211174 609718 211208 610342
rect 211288 609718 211322 610342
rect 211334 610330 211335 610331
rect 211933 610330 211934 610331
rect 211333 610329 211334 610330
rect 211934 610329 211935 610330
rect 211333 609730 211334 609731
rect 211934 609730 211935 609731
rect 211334 609729 211335 609730
rect 211933 609729 211934 609730
rect 211946 609718 211980 610342
rect 211992 610330 211993 610331
rect 212591 610330 212592 610331
rect 211991 610329 211992 610330
rect 212592 610329 212593 610330
rect 212604 610194 212638 610342
rect 212650 610330 212651 610331
rect 213249 610330 213250 610331
rect 212649 610329 212650 610330
rect 213250 610329 213251 610330
rect 212586 609742 212660 610194
rect 211991 609730 211992 609731
rect 211992 609729 211993 609730
rect 212190 609718 212660 609742
rect 213250 609730 213251 609731
rect 213249 609729 213250 609730
rect 213262 609718 213296 610342
rect 213308 610330 213309 610331
rect 213307 610329 213308 610330
rect 213630 610314 213702 610352
rect 213668 609746 213702 610314
rect 213307 609730 213308 609731
rect 213308 609729 213309 609730
rect 213618 609718 213629 609729
rect 211174 609684 213629 609718
rect 211174 609604 211208 609684
rect 211288 609604 211322 609684
rect 211946 609604 211980 609684
rect 212190 609650 212660 609684
rect 212586 609604 212660 609650
rect 213262 609604 213296 609684
rect 213770 609604 213804 613088
rect 214692 610698 214726 615632
rect 215148 615142 215520 615632
rect 217628 615388 217640 615670
rect 217662 615422 217674 615644
rect 214778 615014 215520 615142
rect 214778 614822 215220 615014
rect 226746 614020 226946 614042
rect 213884 610360 213898 610382
rect 215336 610006 215370 610698
rect 215450 610006 215474 610040
rect 215242 609972 215536 610006
rect 215336 609938 215370 609972
rect 215336 609870 215394 609938
rect 215468 609877 215484 609972
rect 215336 609614 215370 609870
rect 215388 609619 215404 609827
rect 215416 609811 215422 609827
rect 215412 609635 215422 609811
rect 215416 609619 215422 609635
rect 215438 609623 215488 609877
rect 215310 609610 215374 609614
rect 215310 609604 215394 609610
rect 205456 609570 213804 609604
rect 203868 609140 203914 609172
rect 203868 608838 203888 609140
rect 203924 609112 203942 609172
rect 205128 609104 205142 609172
rect 205822 609132 205856 609166
rect 205936 609132 205970 609570
rect 206067 609534 209691 609570
rect 206390 609474 206424 609534
rect 206746 609474 206780 609534
rect 206875 609482 206909 609534
rect 206390 609440 206780 609474
rect 206144 609396 206216 609438
rect 206808 609396 206909 609482
rect 206144 609362 206230 609396
rect 206154 609324 206230 609362
rect 206372 609198 206794 609390
rect 206372 609172 206840 609198
rect 206372 609170 206794 609172
rect 205598 609098 206050 609132
rect 199429 608824 199475 608836
rect 205598 608816 205632 609098
rect 205822 609018 205856 609098
rect 205936 609024 205970 609098
rect 205936 609018 205972 609024
rect 205662 608974 205734 609012
rect 205784 609004 205972 609018
rect 205784 608984 205970 609004
rect 205700 608940 205734 608974
rect 205809 608972 205810 608973
rect 205810 608971 205811 608972
rect 205810 608942 205811 608943
rect 205809 608941 205810 608942
rect 205822 608930 205856 608984
rect 205936 608930 205970 608984
rect 205784 608896 205970 608930
rect 205822 608870 205856 608896
rect 205810 608838 205868 608870
rect 205822 608834 205856 608838
rect 205694 608816 205828 608834
rect 205936 608816 205970 608896
rect 205598 608782 206050 608816
rect 205936 608760 205970 608782
rect 206067 608746 206182 609168
rect 206372 609150 206840 609170
rect 206232 609116 206840 609150
rect 206232 609088 206266 609116
rect 206198 609054 206266 609088
rect 206232 608856 206285 609054
rect 206287 608974 206368 609021
rect 206334 608936 206368 608974
rect 206232 608794 206266 608856
rect 206372 608811 206798 609116
rect 206875 608836 206909 609396
rect 209507 608836 209541 609534
rect 211174 609288 211208 609570
rect 212586 609540 212660 609570
rect 215336 609542 215394 609604
rect 215450 609597 215460 609623
rect 215450 609585 215456 609597
rect 215336 609484 215370 609542
rect 215396 609488 215400 609576
rect 215424 609508 215456 609576
rect 215468 609508 215484 609623
rect 215336 609474 215374 609484
rect 215424 609474 215484 609508
rect 215502 609474 215536 609972
rect 248056 609972 248446 610006
rect 215242 609440 215536 609474
rect 215674 609462 215694 609576
rect 248056 609474 248090 609972
rect 248270 609904 248317 609951
rect 248232 609870 248317 609904
rect 248159 609811 248204 609822
rect 248287 609811 248332 609822
rect 248170 609635 248204 609811
rect 248298 609635 248332 609811
rect 248270 609576 248317 609623
rect 248232 609542 248317 609576
rect 248412 609474 248446 609972
rect 248056 609440 248446 609474
rect 215336 609390 215374 609440
rect 215424 609432 215456 609440
rect 215424 609390 215428 609432
rect 215300 609288 215550 609390
rect 209590 609268 211232 609288
rect 215300 609282 215682 609288
rect 216036 609282 217398 609288
rect 211174 609232 211208 609268
rect 215300 609232 215550 609282
rect 215674 609232 215694 609276
rect 209590 609212 211232 609232
rect 215300 609226 215694 609232
rect 216036 609226 217342 609232
rect 206328 608794 206798 608811
rect 206232 608760 206798 608794
rect 211174 608760 211208 609212
rect 212506 609084 212520 609172
rect 213256 609104 213270 609172
rect 214046 609104 214070 609172
rect 215300 609026 215550 609226
rect 215674 609204 215694 609226
rect 215674 609092 215694 609158
rect 215366 608976 215400 608986
rect 215382 608942 215434 608952
rect 215348 608908 215372 608942
rect 215382 608874 215406 608942
rect 215480 608840 215514 608852
rect 215258 608806 215514 608840
rect 248038 608770 248460 609390
rect 179764 608329 180384 608714
rect 180434 608666 181000 608700
rect 180434 608534 180468 608666
rect 180589 608596 180626 608620
rect 180806 608597 180845 608620
rect 180805 608596 180845 608597
rect 180805 608592 180816 608596
rect 180489 608534 180570 608571
rect 180617 608568 180626 608592
rect 180805 608586 180817 608592
rect 180629 608571 180817 608586
rect 180629 608568 180898 608571
rect 180629 608552 180816 608568
rect 180817 608534 180898 608568
rect 180966 608534 181000 608666
rect 180434 608513 181090 608534
rect 180400 608479 181090 608513
rect 180434 608467 181090 608479
rect 180436 608460 181090 608467
rect 180613 608445 180821 608458
rect 180617 608433 180817 608445
rect 180434 608406 180468 608433
rect 180613 608424 180821 608433
rect 180617 608412 180817 608424
rect 180966 608406 181000 608433
rect 180579 608398 180855 608399
rect 180468 608365 180966 608398
rect 180468 608331 180966 608344
rect 183086 608329 184232 608572
rect 256394 608420 256406 608702
rect 256428 608454 256440 608676
rect 176310 608210 176338 608266
rect 182742 607910 183290 607944
rect 183376 607926 183410 607944
rect 183908 607926 183942 607944
rect 182782 607876 183324 607890
rect 183340 607856 183978 607926
rect 205648 607858 205794 607876
rect 214404 607858 214550 607876
rect 179658 607440 179692 607794
rect 182536 607736 182918 607760
rect 205738 607754 205800 607800
rect 205866 607754 205950 607800
rect 182564 607708 182918 607732
rect 205738 607726 205828 607750
rect 205838 607726 205894 607750
rect 186136 607694 187240 607720
rect 186108 607666 187268 607692
rect 179220 607406 187472 607440
rect 179270 607258 179290 607360
rect 179298 607286 179346 607332
rect 179270 606600 179290 606702
rect 179298 606628 179346 606674
rect 179658 606542 179692 607406
rect 179729 607330 179832 607338
rect 179722 607326 179832 607330
rect 187286 607326 187297 607337
rect 179722 607292 187297 607326
rect 179744 607280 179832 607292
rect 179742 607210 179754 607250
rect 179714 607182 179754 607194
rect 179760 607146 179794 607280
rect 187298 607264 187370 607302
rect 179800 607210 182742 607250
rect 182942 607210 183142 607250
rect 183342 607210 187330 607250
rect 179800 607182 182742 607194
rect 182942 607182 183142 607194
rect 183342 607182 187330 607194
rect 187336 607130 187370 607264
rect 187438 607250 187472 607406
rect 187376 607210 187472 607250
rect 187376 607182 187408 607194
rect 187298 607118 187386 607130
rect 187438 607118 187472 607210
rect 179722 607056 179794 607094
rect 179844 607084 187386 607118
rect 187404 607084 187472 607118
rect 205886 607108 205894 607726
rect 187298 607072 187386 607084
rect 179760 606680 179794 607056
rect 187336 606696 187370 607072
rect 179744 606672 179832 606680
rect 179722 606668 179832 606672
rect 187286 606668 187297 606679
rect 179722 606634 187297 606668
rect 179744 606622 179832 606634
rect 179736 606558 179754 606598
rect 140869 606258 144717 606269
rect 140869 606246 144706 606258
rect 140869 606235 144717 606246
rect 144758 606235 149271 606269
rect 139388 606152 140078 606162
rect 128126 605362 128746 605784
rect 128796 605732 129362 605766
rect 128796 605410 128830 605732
rect 129167 605652 129178 605663
rect 128851 605590 128932 605637
rect 128991 605618 129178 605652
rect 129179 605590 129260 605637
rect 128898 605552 128932 605590
rect 129226 605552 129260 605590
rect 129167 605524 129178 605535
rect 128991 605490 129178 605524
rect 129328 605410 129362 605732
rect 128796 605376 129362 605410
rect 129526 605378 129552 606150
rect 129560 605344 129586 606150
rect 126854 604616 130166 604654
rect 126910 604560 130110 604598
rect 129560 604511 129594 604545
rect 132618 604511 132652 604545
rect 135676 604511 135710 604545
rect 135790 604511 135824 606150
rect 139336 606138 140524 606152
rect 139416 606124 140050 606134
rect 139280 606082 140580 606124
rect 144758 606066 144792 606235
rect 148680 606199 149271 606235
rect 179326 606094 179346 606542
rect 179658 606502 179754 606542
rect 179270 605942 179290 606044
rect 179298 605970 179346 606016
rect 179658 605884 179692 606502
rect 179760 606488 179794 606622
rect 187298 606606 187370 606644
rect 179800 606558 187330 606598
rect 179800 606502 187330 606542
rect 187336 606472 187370 606606
rect 187438 606598 187472 607084
rect 187376 606558 187472 606598
rect 187376 606502 187412 606542
rect 187298 606460 187386 606472
rect 187438 606460 187472 606558
rect 179722 606398 179794 606436
rect 179844 606426 187386 606460
rect 187404 606426 187472 606460
rect 187298 606414 187386 606426
rect 179760 606022 179794 606398
rect 187336 606038 187370 606414
rect 179744 606014 179832 606022
rect 179722 606010 179832 606014
rect 187286 606010 187297 606021
rect 179722 605976 187297 606010
rect 179744 605964 179832 605976
rect 179748 605894 179754 605912
rect 179658 605838 179754 605884
rect 179270 605284 179290 605386
rect 179298 605312 179346 605358
rect 179270 604626 179290 604728
rect 179298 604654 179346 604700
rect 179658 604568 179692 605838
rect 179760 605830 179794 605964
rect 187298 605948 187370 605986
rect 179804 605912 187330 605940
rect 179800 605894 187330 605912
rect 179800 605838 187330 605884
rect 187336 605814 187370 605948
rect 187438 605940 187472 606426
rect 187376 605894 187472 605940
rect 187376 605838 187408 605884
rect 187298 605802 187386 605814
rect 187438 605802 187472 605894
rect 179722 605740 179794 605778
rect 179844 605768 187386 605802
rect 187404 605768 187472 605802
rect 187298 605756 187386 605768
rect 179760 605364 179794 605740
rect 187336 605380 187370 605756
rect 179744 605356 179832 605364
rect 179722 605352 179832 605356
rect 187286 605352 187297 605363
rect 179722 605318 187297 605352
rect 179744 605306 179832 605318
rect 179760 605172 179794 605306
rect 187298 605290 187370 605328
rect 179860 605236 187330 605276
rect 179804 605180 187330 605220
rect 187336 605156 187370 605290
rect 187438 605276 187472 605768
rect 187376 605236 187472 605276
rect 187376 605180 187396 605220
rect 187298 605144 187386 605156
rect 187438 605144 187472 605236
rect 179722 605082 179794 605120
rect 179844 605110 187386 605144
rect 187404 605110 187472 605144
rect 187298 605098 187386 605110
rect 179760 604706 179794 605082
rect 187336 604722 187370 605098
rect 179744 604698 179832 604706
rect 179722 604694 179832 604698
rect 187286 604694 187297 604705
rect 179722 604660 187297 604694
rect 179744 604648 179832 604660
rect 179748 604584 179754 604596
rect 179658 604528 179754 604568
rect 127897 604477 136167 604511
rect 127897 601934 127931 604477
rect 129560 604397 129594 604477
rect 132618 604397 132652 604477
rect 135676 604397 135710 604477
rect 135790 604397 135824 604477
rect 127952 604335 128033 604382
rect 128092 604363 135824 604397
rect 129547 604351 129548 604352
rect 129548 604350 129549 604351
rect 127999 603767 128033 604335
rect 129258 604322 129314 604336
rect 129258 604266 129314 604280
rect 129548 603751 129549 603752
rect 129547 603750 129548 603751
rect 129560 603739 129594 604363
rect 129606 604351 129607 604352
rect 132605 604351 132606 604352
rect 129605 604350 129606 604351
rect 132606 604350 132607 604351
rect 129605 603751 129606 603752
rect 132606 603751 132607 603752
rect 129606 603750 129607 603751
rect 132605 603750 132606 603751
rect 132618 603739 132652 604363
rect 132664 604351 132665 604352
rect 135663 604351 135664 604352
rect 132663 604350 132664 604351
rect 135664 604350 135665 604351
rect 135392 603832 135448 603838
rect 135392 603776 135448 603782
rect 132663 603751 132664 603752
rect 135664 603751 135665 603752
rect 132664 603750 132665 603751
rect 135663 603750 135664 603751
rect 135676 603739 135710 604363
rect 135790 603739 135824 604363
rect 179658 604372 179692 604528
rect 179760 604514 179794 604648
rect 187298 604632 187370 604670
rect 179800 604584 183276 604596
rect 183476 604584 183676 604596
rect 183876 604584 187330 604596
rect 179800 604528 183276 604568
rect 183476 604528 183676 604568
rect 183876 604528 187330 604568
rect 187336 604498 187370 604632
rect 187376 604584 187430 604596
rect 187376 604528 187402 604568
rect 187298 604486 187386 604498
rect 187438 604486 187472 605110
rect 179844 604455 187386 604486
rect 179844 604452 187401 604455
rect 187404 604452 187472 604486
rect 187298 604440 187401 604452
rect 183736 604372 183742 604410
rect 187438 604372 187472 604452
rect 179658 604338 187910 604372
rect 179270 603968 179290 604070
rect 183098 604046 183452 604070
rect 179298 603996 179346 604042
rect 183070 604018 183452 604042
rect 183736 604028 183742 604338
rect 185574 604086 186734 604112
rect 185602 604058 186706 604084
rect 187438 603984 187472 604338
rect 127952 603677 128033 603724
rect 128092 603705 135824 603739
rect 129258 603699 129362 603700
rect 129547 603693 129548 603694
rect 129548 603692 129549 603693
rect 127999 603109 128033 603677
rect 129258 603643 129306 603644
rect 129258 603174 129314 603178
rect 129258 603118 129314 603122
rect 129548 603093 129549 603094
rect 129547 603092 129548 603093
rect 129560 603081 129594 603705
rect 129606 603693 129607 603694
rect 132605 603693 132606 603694
rect 129605 603692 129606 603693
rect 132606 603692 132607 603693
rect 129605 603093 129606 603094
rect 132606 603093 132607 603094
rect 129606 603092 129607 603093
rect 132605 603092 132606 603093
rect 132618 603081 132652 603705
rect 132664 603693 132665 603694
rect 135663 603693 135664 603694
rect 132663 603692 132664 603693
rect 135664 603692 135665 603693
rect 135392 603654 135448 603678
rect 135392 603598 135448 603622
rect 132663 603093 132664 603094
rect 135664 603093 135665 603094
rect 132664 603092 132665 603093
rect 135663 603092 135664 603093
rect 135676 603081 135710 603705
rect 135790 603081 135824 603705
rect 177554 603614 177598 603964
rect 177610 603614 177654 603964
rect 183222 603888 184530 603922
rect 183316 603854 183824 603868
rect 183874 603852 184512 603888
rect 183276 603553 183310 603571
rect 183790 603553 183824 603571
rect 183240 603517 183860 603553
rect 184006 603517 184380 603530
rect 179215 603483 185078 603517
rect 127952 603019 128033 603066
rect 128092 603047 135824 603081
rect 179230 603064 179850 603483
rect 183240 603482 183860 603483
rect 179900 603449 180434 603468
rect 179934 603434 180432 603449
rect 179900 603409 180466 603415
rect 179900 603406 179934 603409
rect 180432 603406 180466 603409
rect 179866 603403 179968 603406
rect 180398 603403 180500 603406
rect 179866 603400 180500 603403
rect 179866 603369 179934 603400
rect 180057 603388 180309 603392
rect 180045 603369 180321 603388
rect 180398 603369 180500 603400
rect 179900 603112 179934 603369
rect 180271 603354 180282 603357
rect 180079 603339 180287 603354
rect 180294 603339 180402 603346
rect 179955 603292 180036 603339
rect 180079 603335 180402 603339
rect 180095 603320 180282 603335
rect 180283 603328 180402 603335
rect 180283 603318 180364 603328
rect 180283 603300 180374 603318
rect 180283 603292 180364 603300
rect 180002 603254 180036 603292
rect 180330 603254 180364 603292
rect 180271 603226 180282 603237
rect 180095 603192 180282 603226
rect 180432 603112 180466 603369
rect 179900 603078 180466 603112
rect 129547 603035 129548 603036
rect 129548 603034 129549 603035
rect 127999 602451 128033 603019
rect 129258 603014 129314 603016
rect 129258 602958 129314 602960
rect 129548 602435 129549 602436
rect 129547 602434 129548 602435
rect 129560 602423 129594 603047
rect 129606 603035 129607 603036
rect 132605 603035 132606 603036
rect 129605 603034 129606 603035
rect 132606 603034 132607 603035
rect 129605 602435 129606 602436
rect 132606 602435 132607 602436
rect 129606 602434 129607 602435
rect 132605 602434 132606 602435
rect 132618 602423 132652 603047
rect 132664 603035 132665 603036
rect 135663 603035 135664 603036
rect 132663 603034 132664 603035
rect 135664 603034 135665 603035
rect 135392 602512 135448 602528
rect 135392 602456 135448 602472
rect 132663 602435 132664 602436
rect 135664 602435 135665 602436
rect 132664 602434 132665 602435
rect 135663 602434 135664 602435
rect 135676 602423 135710 603047
rect 135790 602423 135824 603047
rect 183692 602819 183714 603108
rect 183720 602819 183770 603080
rect 186080 602838 187052 602844
rect 187451 602819 187485 603421
rect 179635 602785 187905 602819
rect 179274 602677 179290 602779
rect 179302 602705 179346 602751
rect 127952 602361 128033 602408
rect 128092 602389 135824 602423
rect 129547 602377 129548 602378
rect 129548 602376 129549 602377
rect 127999 601934 128033 602361
rect 129560 601993 129594 602389
rect 129606 602377 129607 602378
rect 132605 602377 132606 602378
rect 129605 602376 129606 602377
rect 132606 602376 132607 602377
rect 132618 601993 132652 602389
rect 132664 602377 132665 602378
rect 135663 602377 135664 602378
rect 132663 602376 132664 602377
rect 135664 602376 135665 602377
rect 135392 602288 135448 602290
rect 135676 601993 135710 602389
rect 128079 601981 128080 601982
rect 128080 601980 128081 601981
rect 129532 601934 129579 601981
rect 132590 601934 132637 601981
rect 135648 601934 135695 601981
rect 127897 601900 129579 601934
rect 129622 601900 132637 601934
rect 132680 601900 135695 601934
rect 127897 601832 127931 601900
rect 127999 601832 128033 601900
rect 135790 601832 135824 602389
rect 179274 602019 179290 602121
rect 179302 602047 179346 602093
rect 149330 601872 149388 601934
rect 149390 601872 149448 601874
rect 126484 601798 135824 601832
rect 127897 601055 127931 601798
rect 128382 601786 129314 601798
rect 179274 601361 179290 601463
rect 179302 601389 179346 601435
rect 179274 600703 179290 600805
rect 179302 600731 179346 600777
rect 140356 600218 141276 600222
rect 141546 600218 142466 600222
rect 142856 600210 143776 600222
rect 132136 600168 132774 600204
rect 144024 600202 144944 600222
rect 145184 600198 148736 600222
rect 125638 600134 132774 600168
rect 145150 600164 148770 600168
rect 127058 595908 127060 596210
rect 127114 595964 127116 596210
rect 127172 595434 127206 599982
rect 131538 599944 131572 600134
rect 131640 600068 131674 600118
rect 131684 600066 131704 600072
rect 131712 600066 131730 600100
rect 131782 600070 131934 600092
rect 131766 600066 131934 600070
rect 131950 600068 131984 600118
rect 131602 600032 131704 600066
rect 131708 600058 131742 600066
rect 131712 600048 131732 600058
rect 131766 600048 132022 600066
rect 131712 600032 132022 600048
rect 131684 600026 131704 600032
rect 131708 600024 131912 600032
rect 131712 600012 131912 600024
rect 131714 599998 131732 600012
rect 131720 599990 131754 599998
rect 131720 599944 131754 599978
rect 132052 599944 132086 600134
rect 131538 599910 132086 599944
rect 132136 599856 132774 600134
rect 135062 600092 135262 600104
rect 135034 600064 135290 600076
rect 128688 599440 128722 599474
rect 129446 599440 129480 599474
rect 130204 599440 130238 599474
rect 130962 599440 130996 599474
rect 131720 599440 131754 599474
rect 132478 599440 132512 599474
rect 133236 599440 133270 599474
rect 133994 599440 134028 599474
rect 134752 599440 134786 599474
rect 135510 599440 135544 599474
rect 127920 599406 136268 599440
rect 127920 599378 127954 599406
rect 127920 599304 127988 599378
rect 128688 599326 128722 599406
rect 129446 599326 129480 599406
rect 130204 599326 130238 599406
rect 130962 599326 130996 599406
rect 131720 599326 131754 599406
rect 132478 599326 132512 599406
rect 133236 599326 133270 599406
rect 133994 599326 134028 599406
rect 134752 599326 134786 599406
rect 135510 599326 135544 599406
rect 136082 599326 136093 599337
rect 127920 599302 128010 599304
rect 127920 599276 128056 599302
rect 127920 599264 128062 599276
rect 127920 599194 128010 599264
rect 128016 599194 128062 599264
rect 128068 599194 128090 599304
rect 128106 599292 136093 599326
rect 128675 599280 128676 599281
rect 128676 599279 128677 599280
rect 127920 598746 127988 599194
rect 128022 598746 128056 599194
rect 127920 598656 128010 598746
rect 128016 598696 128062 598746
rect 128016 598684 128038 598696
rect 128040 598684 128062 598696
rect 128068 598656 128090 598746
rect 128676 598680 128677 598681
rect 128675 598679 128676 598680
rect 128688 598668 128722 599292
rect 128734 599280 128735 599281
rect 129433 599280 129434 599281
rect 128733 599279 128734 599280
rect 129434 599279 129435 599280
rect 128733 598680 128734 598681
rect 129434 598680 129435 598681
rect 128734 598679 128735 598680
rect 129433 598679 129434 598680
rect 129446 598668 129480 599292
rect 129492 599280 129493 599281
rect 130191 599280 130192 599281
rect 129491 599279 129492 599280
rect 130192 599279 130193 599280
rect 129491 598680 129492 598681
rect 130192 598680 130193 598681
rect 129492 598679 129493 598680
rect 130191 598679 130192 598680
rect 130204 598668 130238 599292
rect 130250 599280 130251 599281
rect 130949 599280 130950 599281
rect 130249 599279 130250 599280
rect 130950 599279 130951 599280
rect 130249 598680 130250 598681
rect 130950 598680 130951 598681
rect 130250 598679 130251 598680
rect 130949 598679 130950 598680
rect 130962 598668 130996 599292
rect 131008 599280 131009 599281
rect 131707 599280 131708 599281
rect 131007 599279 131008 599280
rect 131708 599279 131709 599280
rect 131007 598680 131008 598681
rect 131708 598680 131709 598681
rect 131008 598679 131009 598680
rect 131707 598679 131708 598680
rect 131720 598668 131754 599292
rect 131766 599280 131767 599281
rect 132465 599280 132466 599281
rect 131765 599279 131766 599280
rect 132466 599279 132467 599280
rect 131765 598680 131766 598681
rect 132466 598680 132467 598681
rect 131766 598679 131767 598680
rect 132465 598679 132466 598680
rect 132478 598668 132512 599292
rect 132524 599280 132525 599281
rect 133223 599280 133224 599281
rect 132523 599279 132524 599280
rect 133224 599279 133225 599280
rect 132523 598680 132524 598681
rect 133224 598680 133225 598681
rect 132524 598679 132525 598680
rect 133223 598679 133224 598680
rect 133236 598668 133270 599292
rect 133282 599280 133283 599281
rect 133981 599280 133982 599281
rect 133281 599279 133282 599280
rect 133982 599279 133983 599280
rect 133281 598680 133282 598681
rect 133982 598680 133983 598681
rect 133282 598679 133283 598680
rect 133981 598679 133982 598680
rect 133994 598668 134028 599292
rect 134040 599280 134041 599281
rect 134739 599280 134740 599281
rect 134039 599279 134040 599280
rect 134740 599279 134741 599280
rect 134039 598680 134040 598681
rect 134740 598680 134741 598681
rect 134040 598679 134041 598680
rect 134739 598679 134740 598680
rect 134752 598668 134786 599292
rect 134798 599280 134799 599281
rect 135497 599280 135498 599281
rect 134797 599279 134798 599280
rect 135498 599279 135499 599280
rect 134797 598680 134798 598681
rect 135498 598680 135499 598681
rect 134798 598679 134799 598680
rect 135497 598679 135498 598680
rect 135510 598668 135544 599292
rect 135556 599280 135557 599281
rect 135555 599279 135556 599280
rect 136094 599264 136166 599302
rect 136132 598696 136166 599264
rect 135555 598680 135556 598681
rect 135556 598679 135557 598680
rect 136082 598668 136093 598679
rect 127920 598646 127988 598656
rect 127920 598644 128010 598646
rect 127920 598618 128056 598644
rect 127920 598606 128062 598618
rect 127920 598488 128010 598606
rect 127920 597986 127988 598488
rect 128016 598460 128062 598606
rect 128022 598038 128062 598460
rect 128040 598026 128062 598038
rect 128068 597998 128090 598646
rect 128106 598634 136093 598668
rect 128675 598622 128676 598623
rect 128676 598621 128677 598622
rect 128676 598022 128677 598023
rect 128675 598021 128676 598022
rect 128688 598010 128722 598634
rect 128734 598622 128735 598623
rect 129433 598622 129434 598623
rect 128733 598621 128734 598622
rect 129434 598621 129435 598622
rect 129446 598028 129480 598634
rect 129492 598622 129493 598623
rect 130191 598622 130192 598623
rect 129491 598621 129492 598622
rect 130192 598621 130193 598622
rect 128733 598022 128734 598023
rect 128734 598021 128735 598022
rect 128796 598010 129480 598028
rect 129491 598022 129492 598023
rect 130192 598022 130193 598023
rect 129492 598021 129493 598022
rect 130191 598021 130192 598022
rect 130204 598010 130238 598634
rect 130250 598622 130251 598623
rect 130949 598622 130950 598623
rect 130249 598621 130250 598622
rect 130950 598621 130951 598622
rect 130249 598022 130250 598023
rect 130950 598022 130951 598023
rect 130250 598021 130251 598022
rect 130949 598021 130950 598022
rect 130962 598010 130996 598634
rect 131008 598622 131009 598623
rect 131707 598622 131708 598623
rect 131007 598621 131008 598622
rect 131708 598621 131709 598622
rect 131007 598022 131008 598023
rect 131708 598022 131709 598023
rect 131008 598021 131009 598022
rect 131707 598021 131708 598022
rect 131720 598010 131754 598634
rect 131766 598622 131767 598623
rect 132465 598622 132466 598623
rect 131765 598621 131766 598622
rect 132466 598621 132467 598622
rect 131765 598022 131766 598023
rect 132466 598022 132467 598023
rect 131766 598021 131767 598022
rect 132465 598021 132466 598022
rect 131942 598010 132264 598012
rect 132478 598010 132512 598634
rect 132524 598622 132525 598623
rect 133223 598622 133224 598623
rect 132523 598621 132524 598622
rect 133224 598621 133225 598622
rect 132523 598022 132524 598023
rect 133224 598022 133225 598023
rect 132524 598021 132525 598022
rect 133223 598021 133224 598022
rect 133236 598010 133270 598634
rect 133282 598622 133283 598623
rect 133981 598622 133982 598623
rect 133281 598621 133282 598622
rect 133982 598621 133983 598622
rect 133281 598022 133282 598023
rect 133982 598022 133983 598023
rect 133282 598021 133283 598022
rect 133981 598021 133982 598022
rect 133994 598010 134028 598634
rect 134040 598622 134041 598623
rect 134739 598622 134740 598623
rect 134039 598621 134040 598622
rect 134740 598621 134741 598622
rect 134039 598022 134040 598023
rect 134740 598022 134741 598023
rect 134040 598021 134041 598022
rect 134739 598021 134740 598022
rect 134752 598010 134786 598634
rect 134798 598622 134799 598623
rect 135497 598622 135498 598623
rect 134797 598621 134798 598622
rect 135498 598621 135499 598622
rect 134797 598022 134798 598023
rect 135498 598022 135499 598023
rect 134798 598021 134799 598022
rect 135497 598021 135498 598022
rect 135510 598010 135544 598634
rect 135556 598622 135557 598623
rect 135555 598621 135556 598622
rect 136094 598606 136166 598644
rect 136132 598038 136166 598606
rect 135555 598022 135556 598023
rect 135556 598021 135557 598022
rect 136082 598010 136093 598021
rect 127920 597960 128056 597986
rect 127920 597948 128062 597960
rect 127920 597328 127988 597948
rect 128022 597884 128062 597948
rect 128068 597884 128090 597988
rect 128106 597976 136093 598010
rect 128675 597964 128676 597965
rect 128676 597963 128677 597964
rect 128022 597436 128056 597884
rect 128022 597380 128062 597436
rect 128040 597368 128062 597380
rect 128068 597340 128090 597436
rect 128676 597364 128677 597365
rect 128675 597363 128676 597364
rect 128688 597352 128722 597976
rect 128734 597964 128735 597965
rect 128733 597963 128734 597964
rect 128796 597954 129480 597976
rect 129492 597964 129493 597965
rect 130191 597964 130192 597965
rect 129491 597963 129492 597964
rect 130192 597963 130193 597964
rect 128902 597496 129224 597954
rect 128733 597364 128734 597365
rect 129434 597364 129435 597365
rect 128734 597363 128735 597364
rect 129433 597363 129434 597364
rect 129446 597352 129480 597954
rect 129491 597364 129492 597365
rect 130192 597364 130193 597365
rect 129492 597363 129493 597364
rect 130191 597363 130192 597364
rect 130204 597352 130238 597976
rect 130250 597964 130251 597965
rect 130949 597964 130950 597965
rect 130249 597963 130250 597964
rect 130950 597963 130951 597964
rect 130249 597364 130250 597365
rect 130950 597364 130951 597365
rect 130250 597363 130251 597364
rect 130949 597363 130950 597364
rect 130962 597352 130996 597976
rect 131008 597964 131009 597965
rect 131707 597964 131708 597965
rect 131007 597963 131008 597964
rect 131708 597963 131709 597964
rect 131007 597364 131008 597365
rect 131708 597364 131709 597365
rect 131008 597363 131009 597364
rect 131707 597363 131708 597364
rect 131720 597352 131754 597976
rect 131766 597964 131767 597965
rect 131765 597963 131766 597964
rect 131942 597768 132264 597976
rect 132465 597964 132466 597965
rect 132466 597963 132467 597964
rect 131794 597556 132264 597768
rect 131942 597504 132264 597556
rect 131765 597364 131766 597365
rect 132466 597364 132467 597365
rect 131766 597363 131767 597364
rect 132465 597363 132466 597364
rect 132478 597352 132512 597976
rect 132524 597964 132525 597965
rect 133223 597964 133224 597965
rect 132523 597963 132524 597964
rect 133224 597963 133225 597964
rect 132523 597364 132524 597365
rect 133224 597364 133225 597365
rect 132524 597363 132525 597364
rect 133223 597363 133224 597364
rect 133236 597352 133270 597976
rect 133282 597964 133283 597965
rect 133981 597964 133982 597965
rect 133281 597963 133282 597964
rect 133982 597963 133983 597964
rect 133281 597364 133282 597365
rect 133982 597364 133983 597365
rect 133282 597363 133283 597364
rect 133981 597363 133982 597364
rect 133994 597352 134028 597976
rect 134040 597964 134041 597965
rect 134739 597964 134740 597965
rect 134039 597963 134040 597964
rect 134740 597963 134741 597964
rect 134039 597364 134040 597365
rect 134740 597364 134741 597365
rect 134040 597363 134041 597364
rect 134739 597363 134740 597364
rect 134752 597352 134786 597976
rect 134798 597964 134799 597965
rect 135497 597964 135498 597965
rect 134797 597963 134798 597964
rect 135498 597963 135499 597964
rect 135510 597420 135544 597976
rect 135556 597964 135557 597965
rect 135555 597963 135556 597964
rect 136094 597948 136166 597986
rect 134797 597364 134798 597365
rect 134798 597363 134799 597364
rect 135476 597358 135500 597392
rect 135504 597358 135544 597420
rect 136132 597380 136166 597948
rect 135555 597364 135556 597365
rect 135556 597363 135557 597364
rect 135510 597352 135544 597358
rect 136082 597352 136093 597363
rect 127920 597302 128056 597328
rect 127920 597290 128062 597302
rect 127920 596670 127988 597290
rect 128022 597220 128062 597290
rect 128068 597220 128090 597330
rect 128106 597318 136093 597352
rect 128675 597306 128676 597307
rect 128676 597305 128677 597306
rect 128022 596772 128056 597220
rect 128022 596722 128062 596772
rect 128040 596710 128062 596722
rect 128068 596682 128090 596772
rect 128676 596706 128677 596707
rect 128675 596705 128676 596706
rect 128688 596694 128722 597318
rect 128734 597306 128735 597307
rect 129433 597306 129434 597307
rect 128733 597305 128734 597306
rect 129434 597305 129435 597306
rect 128733 596706 128734 596707
rect 129434 596706 129435 596707
rect 128734 596705 128735 596706
rect 129433 596705 129434 596706
rect 129446 596694 129480 597318
rect 129492 597306 129493 597307
rect 130191 597306 130192 597307
rect 129491 597305 129492 597306
rect 130192 597305 130193 597306
rect 129491 596706 129492 596707
rect 130192 596706 130193 596707
rect 129492 596705 129493 596706
rect 130191 596705 130192 596706
rect 130204 596694 130238 597318
rect 130250 597306 130251 597307
rect 130949 597306 130950 597307
rect 130249 597305 130250 597306
rect 130950 597305 130951 597306
rect 130249 596706 130250 596707
rect 130950 596706 130951 596707
rect 130250 596705 130251 596706
rect 130949 596705 130950 596706
rect 130962 596694 130996 597318
rect 131008 597306 131009 597307
rect 131707 597306 131708 597307
rect 131007 597305 131008 597306
rect 131708 597305 131709 597306
rect 131007 596706 131008 596707
rect 131708 596706 131709 596707
rect 131008 596705 131009 596706
rect 131707 596705 131708 596706
rect 131720 596694 131754 597318
rect 131766 597306 131767 597307
rect 132465 597306 132466 597307
rect 131765 597305 131766 597306
rect 132466 597305 132467 597306
rect 131765 596706 131766 596707
rect 132466 596706 132467 596707
rect 131766 596705 131767 596706
rect 132465 596705 132466 596706
rect 132478 596694 132512 597318
rect 132524 597306 132525 597307
rect 133223 597306 133224 597307
rect 132523 597305 132524 597306
rect 133224 597305 133225 597306
rect 132523 596706 132524 596707
rect 133224 596706 133225 596707
rect 132524 596705 132525 596706
rect 133223 596705 133224 596706
rect 133236 596694 133270 597318
rect 133282 597306 133283 597307
rect 133981 597306 133982 597307
rect 133281 597305 133282 597306
rect 133982 597305 133983 597306
rect 133281 596706 133282 596707
rect 133982 596706 133983 596707
rect 133282 596705 133283 596706
rect 133981 596705 133982 596706
rect 133994 596694 134028 597318
rect 134040 597306 134041 597307
rect 134739 597306 134740 597307
rect 134039 597305 134040 597306
rect 134740 597305 134741 597306
rect 134039 596706 134040 596707
rect 134740 596706 134741 596707
rect 134040 596705 134041 596706
rect 134739 596705 134740 596706
rect 134752 596694 134786 597318
rect 135510 597312 135544 597318
rect 134798 597306 134799 597307
rect 134797 597305 134798 597306
rect 135476 597256 135500 597312
rect 135504 597228 135544 597312
rect 135556 597306 135557 597307
rect 135555 597305 135556 597306
rect 136094 597290 136166 597328
rect 134797 596706 134798 596707
rect 135498 596706 135499 596707
rect 134798 596705 134799 596706
rect 135497 596705 135498 596706
rect 135510 596694 135544 597228
rect 136132 596722 136166 597290
rect 136190 596772 136192 597052
rect 136218 596744 136220 597024
rect 135555 596706 135556 596707
rect 135556 596705 135557 596706
rect 136082 596694 136093 596705
rect 127920 596644 128056 596670
rect 127920 596632 128062 596644
rect 127920 595984 127988 596632
rect 128022 596568 128062 596632
rect 128068 596568 128090 596672
rect 128106 596660 136093 596694
rect 128675 596648 128676 596649
rect 128676 596647 128677 596648
rect 128022 596120 128056 596568
rect 128022 596064 128062 596120
rect 128040 596052 128062 596064
rect 128068 596024 128090 596120
rect 128676 596048 128677 596049
rect 128675 596047 128676 596048
rect 128688 596036 128722 596660
rect 128734 596648 128735 596649
rect 129433 596648 129434 596649
rect 128733 596647 128734 596648
rect 129434 596647 129435 596648
rect 128733 596048 128734 596049
rect 129434 596048 129435 596049
rect 128734 596047 128735 596048
rect 129433 596047 129434 596048
rect 129446 596036 129480 596660
rect 129492 596648 129493 596649
rect 130191 596648 130192 596649
rect 129491 596647 129492 596648
rect 130192 596647 130193 596648
rect 129491 596048 129492 596049
rect 130192 596048 130193 596049
rect 129492 596047 129493 596048
rect 130191 596047 130192 596048
rect 130204 596036 130238 596660
rect 130250 596648 130251 596649
rect 130949 596648 130950 596649
rect 130249 596647 130250 596648
rect 130950 596647 130951 596648
rect 130249 596048 130250 596049
rect 130950 596048 130951 596049
rect 130250 596047 130251 596048
rect 130949 596047 130950 596048
rect 130962 596036 130996 596660
rect 131008 596648 131009 596649
rect 131707 596648 131708 596649
rect 131007 596647 131008 596648
rect 131708 596647 131709 596648
rect 131720 596302 131754 596660
rect 131766 596648 131767 596649
rect 132465 596648 132466 596649
rect 131765 596647 131766 596648
rect 132466 596647 132467 596648
rect 131776 596302 132224 596456
rect 131676 596244 132224 596302
rect 131676 596154 131796 596244
rect 131007 596048 131008 596049
rect 131708 596048 131709 596049
rect 131008 596047 131009 596048
rect 131707 596047 131708 596048
rect 131720 596036 131754 596154
rect 131765 596048 131766 596049
rect 132466 596048 132467 596049
rect 131766 596047 131767 596048
rect 132465 596047 132466 596048
rect 132478 596036 132512 596660
rect 132524 596648 132525 596649
rect 133223 596648 133224 596649
rect 132523 596647 132524 596648
rect 133224 596647 133225 596648
rect 132523 596048 132524 596049
rect 133224 596048 133225 596049
rect 132524 596047 132525 596048
rect 133223 596047 133224 596048
rect 133236 596036 133270 596660
rect 133282 596648 133283 596649
rect 133981 596648 133982 596649
rect 133281 596647 133282 596648
rect 133982 596647 133983 596648
rect 133281 596048 133282 596049
rect 133982 596048 133983 596049
rect 133282 596047 133283 596048
rect 133981 596047 133982 596048
rect 133994 596036 134028 596660
rect 134040 596648 134041 596649
rect 134739 596648 134740 596649
rect 134039 596647 134040 596648
rect 134740 596647 134741 596648
rect 134039 596048 134040 596049
rect 134740 596048 134741 596049
rect 134040 596047 134041 596048
rect 134739 596047 134740 596048
rect 134752 596036 134786 596660
rect 134798 596648 134799 596649
rect 135497 596648 135498 596649
rect 134797 596647 134798 596648
rect 135498 596647 135499 596648
rect 135510 596112 135544 596660
rect 135556 596648 135557 596649
rect 135555 596647 135556 596648
rect 136094 596632 136166 596670
rect 134797 596048 134798 596049
rect 134798 596047 134799 596048
rect 135476 596042 135502 596084
rect 135504 596042 135544 596112
rect 136132 596064 136166 596632
rect 136190 596120 136198 596568
rect 136218 596092 136226 596596
rect 135555 596048 135556 596049
rect 135556 596047 135557 596048
rect 135510 596036 135544 596042
rect 136082 596036 136093 596047
rect 128106 596002 136093 596036
rect 127920 595922 127964 595984
rect 128688 595922 128722 596002
rect 129446 595922 129480 596002
rect 130204 595922 130238 596002
rect 130962 595922 130996 596002
rect 131720 595922 131754 596002
rect 132478 595922 132512 596002
rect 133236 595922 133270 596002
rect 133994 595922 134028 596002
rect 134752 595922 134786 596002
rect 135510 595996 135544 596002
rect 135476 595948 135502 595996
rect 135504 595922 135544 595996
rect 136234 595922 136268 599406
rect 139922 599210 140090 599324
rect 139922 599154 140134 599210
rect 140014 599062 140134 599154
rect 140074 599034 140092 599058
rect 140070 598730 140092 599034
rect 140108 598898 140216 599024
rect 140108 598768 140130 598898
rect 140296 598596 142604 600034
rect 142874 598590 145182 600028
rect 145364 598322 145398 599982
rect 144830 598010 146480 598322
rect 141044 597826 141366 597966
rect 142554 597826 142876 598000
rect 144076 597826 144398 598002
rect 141044 597494 144398 597826
rect 144824 597502 146480 598010
rect 141044 597464 144284 597494
rect 140970 597458 144284 597464
rect 140970 597294 141138 597458
rect 141318 596888 144284 597458
rect 144830 596884 146480 597502
rect 146916 596886 148566 598324
rect 149020 596884 152370 600204
rect 167170 600102 168684 600116
rect 166904 600050 166928 600086
rect 166882 600040 166928 600050
rect 179274 600045 179290 600147
rect 179302 600073 179346 600119
rect 174054 599984 174124 600030
rect 179635 599999 179669 602785
rect 183692 602754 183714 602785
rect 183720 602754 183770 602785
rect 187343 602761 187389 602785
rect 187349 602757 187383 602761
rect 179792 602739 187290 602743
rect 179780 602717 187306 602739
rect 187315 602733 187417 602756
rect 179780 602711 187417 602717
rect 187302 602705 187417 602711
rect 187451 602705 187485 602785
rect 179814 602699 187383 602705
rect 179690 602643 179771 602690
rect 179814 602677 187399 602699
rect 179830 602671 187399 602677
rect 187417 602671 187519 602705
rect 179922 602665 179956 602671
rect 179724 602140 179731 602156
rect 179696 602112 179731 602128
rect 179737 602099 179771 602643
rect 179922 602637 179928 602660
rect 187302 602659 187399 602671
rect 179777 602140 181056 602156
rect 179777 602112 181028 602128
rect 187349 602115 187383 602659
rect 179721 602087 179818 602099
rect 180030 602087 180684 602108
rect 187290 602093 187301 602098
rect 186080 602087 187302 602093
rect 179721 602084 187302 602087
rect 179721 602081 187301 602084
rect 179721 602060 187306 602081
rect 179721 602059 187383 602060
rect 179780 602053 187417 602059
rect 180030 602047 181180 602053
rect 187302 602047 187417 602053
rect 187451 602047 187485 602671
rect 179814 602041 187383 602047
rect 179690 602025 179771 602032
rect 179690 602020 179805 602025
rect 179690 601997 179771 602020
rect 179814 602019 187399 602041
rect 179830 602013 187399 602019
rect 187417 602013 187519 602047
rect 179690 601992 179777 601997
rect 180526 601994 181180 602013
rect 187302 602001 187399 602013
rect 179690 601985 179771 601992
rect 179737 601441 179771 601985
rect 180120 601976 181522 601994
rect 180092 601948 181550 601966
rect 185622 601488 187030 601506
rect 185650 601460 187002 601478
rect 187349 601462 187383 602001
rect 187343 601445 187389 601462
rect 179721 601429 179818 601441
rect 187290 601429 187301 601440
rect 179721 601423 187301 601429
rect 179721 601402 187306 601423
rect 187315 601417 187417 601434
rect 179721 601401 187383 601402
rect 179780 601395 187417 601401
rect 187302 601389 187417 601395
rect 187451 601389 187485 602013
rect 199468 601434 199469 607108
rect 205942 607052 205950 607754
rect 205952 602866 206658 602902
rect 206755 602866 206789 607795
rect 214494 607754 214556 607800
rect 214622 607754 214706 607800
rect 214494 607726 214584 607750
rect 214594 607726 214650 607750
rect 214698 607052 214706 607754
rect 212564 603092 212570 603292
rect 212592 603064 212598 603320
rect 205952 602832 207354 602866
rect 179814 601383 187383 601389
rect 179690 601327 179771 601374
rect 179814 601361 187399 601383
rect 179830 601355 187399 601361
rect 187417 601355 187519 601389
rect 187302 601343 187399 601355
rect 179724 600818 179731 600836
rect 179696 600790 179731 600808
rect 179737 600783 179771 601327
rect 186166 601306 187343 601324
rect 186138 601278 187343 601296
rect 179777 600818 181034 600836
rect 179777 600790 181006 600808
rect 187349 600799 187383 601343
rect 187389 601306 187430 601324
rect 187389 601278 187402 601296
rect 179721 600771 179818 600783
rect 180010 600771 180664 600790
rect 187290 600771 187301 600782
rect 179721 600765 187301 600771
rect 179721 600744 187306 600765
rect 179721 600743 187383 600744
rect 179780 600737 187417 600743
rect 180010 600731 181200 600737
rect 187302 600731 187417 600737
rect 187451 600731 187485 601355
rect 179814 600725 187383 600731
rect 179690 600709 179771 600716
rect 179690 600700 179805 600709
rect 179814 600703 187399 600725
rect 179690 600681 179771 600700
rect 179830 600697 187399 600703
rect 187417 600697 187519 600731
rect 179690 600672 179777 600681
rect 180546 600676 181200 600697
rect 185564 600691 187028 600697
rect 187302 600685 187399 600697
rect 179690 600669 179771 600672
rect 179737 600125 179771 600669
rect 180142 600656 181544 600672
rect 180114 600628 181572 600644
rect 187349 600152 187383 600685
rect 187343 600129 187389 600152
rect 179721 600113 179818 600125
rect 187290 600113 187301 600124
rect 179721 600107 187301 600113
rect 179721 600085 187306 600107
rect 187315 600101 187417 600124
rect 179780 600079 187306 600085
rect 179814 600045 187340 600073
rect 179830 600041 187328 600045
rect 179737 600011 179771 600033
rect 187451 599999 187485 600697
rect 174054 599956 174068 599978
rect 179215 599965 187485 599999
rect 199468 600032 199496 601434
rect 169948 599400 170220 599404
rect 166932 599386 173264 599400
rect 169932 599384 170232 599386
rect 169932 599380 170230 599384
rect 166960 599352 173264 599372
rect 179635 599363 179669 599965
rect 186104 599940 187028 599946
rect 199468 599723 199469 600032
rect 200708 600010 200724 601412
rect 199429 599720 199469 599723
rect 199423 599708 199469 599720
rect 204244 599512 205182 601880
rect 205952 600664 206658 602832
rect 206755 602752 206789 602832
rect 206869 602752 206903 602832
rect 207159 602752 207170 602763
rect 206721 602718 207170 602752
rect 206755 602094 206789 602718
rect 206869 602688 206903 602718
rect 206915 602706 206916 602707
rect 206914 602705 206915 602706
rect 207171 602690 207252 602737
rect 206869 602658 206909 602688
rect 206928 602686 206937 602688
rect 206869 602094 206903 602658
rect 207218 602122 207252 602690
rect 206914 602106 206915 602107
rect 206915 602105 206916 602106
rect 207159 602094 207170 602105
rect 206721 602060 207170 602094
rect 206755 601436 206789 602060
rect 206869 601436 206903 602060
rect 206915 602048 206916 602049
rect 206914 602047 206915 602048
rect 207171 602032 207252 602079
rect 207218 601464 207252 602032
rect 206914 601448 206915 601449
rect 206915 601447 206916 601448
rect 207159 601436 207170 601447
rect 206721 601402 207170 601436
rect 206755 600778 206789 601402
rect 206869 601080 206903 601402
rect 206915 601390 206916 601391
rect 206914 601389 206915 601390
rect 207171 601374 207252 601421
rect 207218 601080 207252 601374
rect 206869 600858 206914 601080
rect 207218 600903 207299 601080
rect 207171 600890 207299 600903
rect 207320 600890 207354 602832
rect 207538 601886 208958 602878
rect 214538 601978 214562 602178
rect 214566 601950 214590 602206
rect 207996 601734 208126 601754
rect 208850 601688 208877 601720
rect 206869 600778 206903 600858
rect 207042 600856 207432 600890
rect 206914 600790 206915 600791
rect 206915 600789 206916 600790
rect 207042 600778 207076 600856
rect 207218 600790 207252 600856
rect 207159 600778 207170 600789
rect 207256 600788 207303 600835
rect 206721 600744 207175 600778
rect 207202 600756 207303 600788
rect 207202 600754 207209 600756
rect 207218 600754 207303 600756
rect 206755 600664 206789 600744
rect 206869 600664 206903 600744
rect 207042 600664 207076 600744
rect 207156 600706 207190 600711
rect 207286 600706 207318 600711
rect 207145 600695 207190 600706
rect 207273 600695 207318 600706
rect 207156 600664 207190 600695
rect 207284 600664 207318 600695
rect 207320 600664 207354 600856
rect 205952 600630 207354 600664
rect 205952 600594 206658 600630
rect 205946 600288 206658 600324
rect 206755 600288 206789 600630
rect 207042 600358 207076 600630
rect 207156 600519 207190 600630
rect 207284 600519 207318 600630
rect 207256 600460 207303 600507
rect 207218 600426 207303 600460
rect 207398 600358 207432 600856
rect 207538 600696 208958 601688
rect 214538 601578 214562 601778
rect 214566 601550 214590 601806
rect 208164 600436 208238 600696
rect 208850 600652 208877 600696
rect 208884 600686 208911 600696
rect 209501 600378 209535 600416
rect 207042 600324 207432 600358
rect 205946 600274 207348 600288
rect 205946 600254 207446 600274
rect 205946 599512 206658 600254
rect 206755 600174 206789 600254
rect 206869 600174 206903 600254
rect 207024 600174 207446 600254
rect 206721 600140 207446 600174
rect 206755 599559 206789 600140
rect 206869 599730 206903 600140
rect 206915 600128 206916 600129
rect 206914 600127 206915 600128
rect 206869 599720 206914 599730
rect 207024 599708 207446 600140
rect 206884 599661 207446 599708
rect 206931 599654 207446 599661
rect 206931 599627 207348 599654
rect 207212 599559 207246 599627
rect 207314 599559 207348 599627
rect 207530 599559 209550 600378
rect 206755 599525 209550 599559
rect 166960 599330 169932 599352
rect 170232 599330 173264 599352
rect 182724 599301 183344 599302
rect 179731 599267 185078 599301
rect 181752 599262 181864 599267
rect 182724 599231 183344 599267
rect 183490 599254 183864 599267
rect 166750 599182 167750 599186
rect 168186 599182 169836 599184
rect 170290 599182 173914 599186
rect 166312 599022 166896 599048
rect 166312 599014 166880 599022
rect 164746 598960 164752 598963
rect 164746 598774 164772 598960
rect 166880 598816 166902 598958
rect 167532 598944 167544 598946
rect 167560 598916 167572 598946
rect 164746 598463 164752 598774
rect 166880 598694 167512 598816
rect 167680 598798 167714 599054
rect 166892 598394 167512 598694
rect 167562 598764 167612 598798
rect 167658 598764 168032 598798
rect 167562 598692 167596 598764
rect 167562 598516 167606 598692
rect 167610 598544 167634 598664
rect 167680 598656 167714 598764
rect 167745 598684 167768 598696
rect 167680 598584 167732 598656
rect 167741 598650 167768 598684
rect 167745 598638 167768 598650
rect 167562 598442 167596 598516
rect 167680 598442 167714 598584
rect 167745 598556 167768 598568
rect 167741 598522 167768 598556
rect 167745 598510 167768 598522
rect 167562 598408 167612 598442
rect 167658 598408 168032 598442
rect 167680 597880 167714 598408
rect 168186 598372 168418 599088
rect 166373 597748 167750 597833
rect 168186 597746 169836 597833
rect 161238 597528 161412 597560
rect 161272 597494 161446 597526
rect 161548 597474 161572 597492
rect 161548 597438 161608 597474
rect 161566 597426 161626 597438
rect 161566 597390 161608 597426
rect 152428 597094 152450 597290
rect 161602 596610 161636 597342
rect 164996 597046 165018 597256
rect 164204 596706 164214 596760
rect 164320 596706 164328 596740
rect 166382 596706 166416 597348
rect 166627 596742 166706 597579
rect 170326 597543 170360 599054
rect 173844 597543 173878 599054
rect 166759 597509 174933 597543
rect 170326 597429 170360 597509
rect 170440 597429 170474 597509
rect 171098 597429 171132 597509
rect 171756 597429 171790 597509
rect 172414 597429 172448 597509
rect 173072 597429 173106 597509
rect 173730 597429 173764 597509
rect 173844 597429 173878 597509
rect 166731 597182 166744 597417
rect 170292 597395 173878 597429
rect 166765 597182 166778 597383
rect 166822 596799 166842 596805
rect 166818 596749 166842 596799
rect 166663 596706 166697 596742
rect 166731 596726 166842 596749
rect 166846 596740 166870 596777
rect 170326 596771 170360 597395
rect 170440 596771 170474 597395
rect 170486 597383 170487 597384
rect 171085 597383 171086 597384
rect 170485 597382 170486 597383
rect 171086 597382 171087 597383
rect 170485 596783 170486 596784
rect 171086 596783 171087 596784
rect 170486 596782 170487 596783
rect 171085 596782 171086 596783
rect 171098 596771 171132 597395
rect 171144 597383 171145 597384
rect 171743 597383 171744 597384
rect 171143 597382 171144 597383
rect 171744 597382 171745 597383
rect 171143 596783 171144 596784
rect 171744 596783 171745 596784
rect 171144 596782 171145 596783
rect 171743 596782 171744 596783
rect 171756 596771 171790 597395
rect 171802 597383 171803 597384
rect 172401 597383 172402 597384
rect 171801 597382 171802 597383
rect 172402 597382 172403 597383
rect 171801 596783 171802 596784
rect 172402 596783 172403 596784
rect 171802 596782 171803 596783
rect 172401 596782 172402 596783
rect 172414 596771 172448 597395
rect 172460 597383 172461 597384
rect 173059 597383 173060 597384
rect 172459 597382 172460 597383
rect 173060 597382 173061 597383
rect 172459 596783 172460 596784
rect 173060 596783 173061 596784
rect 172460 596782 172461 596783
rect 173059 596782 173060 596783
rect 173072 596771 173106 597395
rect 173118 597383 173119 597384
rect 173717 597383 173718 597384
rect 173117 597382 173118 597383
rect 173718 597382 173719 597383
rect 173117 596783 173118 596784
rect 173718 596783 173719 596784
rect 173118 596782 173119 596783
rect 173717 596782 173718 596783
rect 173730 596771 173764 597395
rect 173844 596771 173878 597395
rect 174859 597312 174866 597407
rect 174887 597312 174894 597379
rect 185078 596982 187304 597016
rect 166846 596737 167748 596740
rect 170292 596737 173878 596771
rect 174859 596759 174866 596864
rect 174887 596787 174894 596864
rect 183950 596767 187415 596778
rect 183950 596755 187404 596767
rect 166846 596731 166870 596737
rect 166765 596721 166799 596726
rect 166759 596706 166805 596721
rect 162154 596670 163732 596704
rect 160778 596564 160824 596570
rect 160890 596564 160932 596570
rect 160778 596536 160852 596542
rect 160862 596536 160932 596542
rect 160774 596368 160920 596520
rect 160828 596264 160882 596368
rect 161602 596168 161646 596610
rect 127920 595888 136268 595922
rect 161612 595888 161646 596168
rect 162154 596106 162188 596670
rect 162283 596602 162538 596649
rect 162898 596602 162945 596649
rect 162290 596534 162314 596602
rect 162318 596568 162945 596602
rect 162318 596562 162342 596568
rect 162362 596521 162420 596568
rect 162948 596534 162966 596636
rect 163032 596618 163079 596649
rect 162976 596602 162994 596608
rect 163020 596602 163079 596618
rect 163556 596602 163603 596649
rect 162976 596568 163603 596602
rect 162976 596566 162994 596568
rect 163020 596566 163078 596568
rect 162976 596562 163078 596566
rect 163020 596538 163078 596562
rect 162996 596534 163078 596538
rect 162257 596509 162313 596520
rect 162268 596255 162313 596509
rect 162374 596267 162419 596521
rect 162915 596509 162960 596520
rect 162926 596255 162960 596509
rect 162968 596340 162990 596516
rect 162996 596312 163018 596534
rect 163020 596521 163078 596534
rect 163032 596267 163066 596521
rect 163573 596509 163618 596520
rect 163584 596255 163618 596509
rect 162256 596208 162538 596255
rect 162914 596208 162973 596255
rect 163004 596214 163051 596255
rect 162992 596208 163051 596214
rect 163572 596208 163630 596255
rect 162256 596174 162393 596208
rect 162436 596174 163051 596208
rect 163094 596174 163630 596208
rect 163664 596174 163678 596208
rect 162256 596158 162314 596174
rect 162338 596168 162358 596174
rect 162256 596143 162271 596158
rect 162366 596140 162386 596174
rect 162914 596158 162972 596174
rect 162992 596168 163016 596174
rect 163020 596140 163044 596174
rect 163572 596158 163630 596174
rect 163615 596143 163630 596158
rect 162268 596106 162302 596140
rect 162926 596106 162960 596140
rect 163584 596106 163618 596140
rect 163698 596106 163732 596670
rect 164258 596650 164268 596706
rect 164282 596672 167810 596706
rect 164282 596650 164292 596672
rect 164258 596112 164292 596650
rect 164294 596257 164326 596650
rect 164952 596620 164999 596651
rect 164940 596610 164999 596620
rect 165002 596610 165049 596651
rect 165610 596620 165657 596651
rect 164940 596604 165049 596610
rect 165598 596604 165657 596620
rect 165660 596604 165707 596651
rect 166268 596620 166314 596651
rect 166382 596638 166416 596672
rect 166256 596604 166314 596620
rect 166374 596604 166416 596638
rect 164434 596570 165049 596604
rect 165092 596570 165707 596604
rect 165750 596570 166314 596604
rect 164940 596564 165014 596570
rect 164338 596522 164362 596551
rect 164940 596523 164998 596564
rect 165598 596523 165656 596570
rect 166256 596523 166314 596570
rect 166318 596570 166336 596604
rect 166318 596564 166330 596570
rect 166382 596545 166388 596577
rect 166392 596545 166416 596604
rect 166382 596534 166416 596545
rect 164366 596522 164390 596523
rect 164338 596511 164406 596522
rect 164338 596268 164362 596511
rect 164366 596261 164406 596511
rect 164952 596304 164992 596523
rect 165019 596518 165064 596522
rect 165002 596511 165064 596518
rect 165002 596332 165020 596511
rect 164952 596273 164986 596304
rect 165030 596261 165064 596511
rect 165610 596273 165644 596523
rect 165677 596511 165722 596522
rect 165688 596261 165722 596511
rect 166268 596273 166302 596523
rect 166318 596511 166416 596534
rect 166318 596508 166380 596511
rect 164360 596214 164419 596261
rect 164924 596214 164971 596261
rect 165018 596214 165077 596261
rect 165582 596214 165629 596261
rect 165676 596214 165735 596261
rect 166240 596214 166287 596261
rect 164360 596180 164971 596214
rect 165014 596180 165629 596214
rect 165672 596180 166287 596214
rect 164360 596164 164418 596180
rect 165018 596164 165076 596180
rect 165676 596164 165734 596180
rect 164360 596149 164375 596164
rect 164372 596112 164406 596146
rect 165030 596112 165064 596146
rect 165066 596112 165070 596164
rect 165688 596112 165722 596146
rect 166312 596112 166318 596312
rect 166340 596112 166374 596312
rect 166382 596112 166416 596511
rect 161698 596072 163742 596106
rect 164258 596078 166416 596112
rect 166663 596604 166697 596672
rect 166731 596604 166744 596650
rect 166765 596604 166799 596672
rect 166976 596604 167023 596651
rect 167634 596604 167681 596651
rect 166663 596570 167023 596604
rect 167066 596570 167681 596604
rect 162154 595968 162188 596072
rect 162048 595948 162710 595968
rect 162090 595928 162656 595948
rect 162154 595924 162188 595928
rect 162118 595900 162656 595924
rect 162154 595888 162188 595900
rect 163698 595888 163732 596072
rect 164258 595896 164292 596078
rect 165066 595896 165070 596078
rect 127930 595778 127964 595888
rect 127930 595692 128030 595778
rect 127930 595434 127964 595692
rect 128564 595586 128572 595616
rect 128592 595614 128600 595616
rect 128654 595614 128678 595616
rect 128682 595586 128706 595616
rect 128062 595416 128610 595450
rect 128062 595388 128096 595416
rect 128576 595388 128610 595416
rect 128028 595384 128130 595388
rect 128542 595384 128644 595388
rect 128062 595282 128096 595384
rect 128102 595382 128610 595384
rect 128210 595370 128462 595374
rect 128198 595350 128474 595370
rect 128576 595350 128610 595382
rect 128106 595348 128256 595350
rect 128416 595348 128610 595350
rect 128106 595344 128610 595348
rect 128106 595334 128566 595344
rect 128164 595282 128198 595308
rect 128232 595302 128440 595334
rect 128470 595316 128560 595322
rect 128474 595282 128508 595308
rect 128576 595282 128610 595344
rect 128660 595282 129298 595504
rect 161590 595304 161682 595888
rect 162118 595492 162582 595888
rect 162118 595302 162596 595492
rect 162600 595440 162656 595458
rect 162710 595440 162762 595458
rect 125638 595260 129298 595282
rect 125638 595259 128214 595260
rect 125638 595258 128225 595259
rect 128236 595258 129298 595260
rect 125638 595248 129298 595258
rect 128062 595196 128096 595248
rect 128576 595196 128610 595248
rect 128660 595212 129298 595248
rect 137740 594852 140332 594932
rect 162558 594860 162596 595302
rect 162618 594920 162656 595432
rect 162710 595412 162734 595430
rect 162780 595302 163768 595888
rect 137672 594294 140332 594852
rect 137740 594038 140332 594294
rect 164222 593876 165082 595896
rect 165258 593884 166250 595904
rect 164398 593706 164412 593876
rect 164426 593734 164440 593876
rect 163756 592368 163782 593292
rect 163790 592368 163816 593258
rect 165066 592538 165070 593876
rect 165688 593870 165722 593884
rect 165592 593776 165926 593870
rect 165592 593692 166156 593776
rect 165030 592535 165070 592538
rect 165688 592535 165722 593692
rect 166312 592722 166318 596078
rect 166340 592722 166374 596078
rect 166663 595908 166697 596570
rect 166731 596098 166744 596570
rect 166765 596141 166799 596570
rect 166846 596523 166847 596524
rect 166845 596522 166846 596523
rect 166993 596511 167038 596522
rect 167651 596511 167696 596522
rect 166765 596125 166778 596141
rect 166992 596125 166993 596126
rect 166991 596124 166992 596125
rect 167004 596113 167038 596511
rect 167049 596125 167050 596126
rect 167650 596125 167651 596126
rect 167050 596124 167051 596125
rect 167649 596124 167650 596125
rect 167662 596113 167696 596511
rect 167776 596113 167810 596672
rect 170326 596113 170360 596737
rect 170440 596113 170474 596737
rect 170486 596725 170487 596726
rect 171085 596725 171086 596726
rect 170485 596724 170486 596725
rect 171086 596724 171087 596725
rect 170485 596125 170486 596126
rect 171086 596125 171087 596126
rect 170486 596124 170487 596125
rect 171085 596124 171086 596125
rect 171098 596113 171132 596737
rect 171144 596725 171145 596726
rect 171743 596725 171744 596726
rect 171143 596724 171144 596725
rect 171744 596724 171745 596725
rect 171143 596125 171144 596126
rect 171744 596125 171745 596126
rect 171144 596124 171145 596125
rect 171743 596124 171744 596125
rect 171756 596113 171790 596737
rect 171802 596725 171803 596726
rect 172401 596725 172402 596726
rect 171801 596724 171802 596725
rect 172402 596724 172403 596725
rect 171801 596125 171802 596126
rect 172402 596125 172403 596126
rect 171802 596124 171803 596125
rect 172401 596124 172402 596125
rect 172414 596113 172448 596737
rect 172460 596725 172461 596726
rect 173059 596725 173060 596726
rect 172459 596724 172460 596725
rect 173060 596724 173061 596725
rect 172459 596125 172460 596126
rect 173060 596125 173061 596126
rect 172460 596124 172461 596125
rect 173059 596124 173060 596125
rect 173072 596113 173106 596737
rect 173118 596725 173119 596726
rect 173717 596725 173718 596726
rect 173117 596724 173118 596725
rect 173718 596724 173719 596725
rect 173117 596125 173118 596126
rect 173718 596125 173719 596126
rect 173118 596124 173119 596125
rect 173717 596124 173718 596125
rect 173730 596113 173764 596737
rect 173844 596113 173878 596737
rect 174859 596654 174866 596749
rect 183950 596744 187415 596755
rect 174887 596654 174894 596721
rect 183950 596358 183984 596744
rect 184694 596676 184732 596714
rect 185352 596676 185390 596714
rect 186010 596676 186048 596714
rect 186668 596676 186706 596714
rect 187354 596710 187364 596714
rect 184126 596642 184732 596676
rect 184784 596642 185390 596676
rect 185442 596642 186048 596676
rect 186100 596642 186706 596676
rect 186758 596642 187342 596676
rect 187354 596608 187376 596710
rect 187456 596682 187490 598350
rect 206546 598202 206658 598206
rect 207314 598148 207348 599525
rect 207530 599489 209550 599525
rect 207734 597936 208140 597940
rect 204412 597576 204418 597622
rect 204440 597548 204446 597622
rect 204462 597572 204614 597626
rect 204640 597572 204732 597588
rect 204462 597566 204732 597572
rect 204412 597468 204418 597510
rect 204440 597468 204446 597538
rect 204462 597518 204718 597566
rect 204462 597480 204614 597518
rect 208646 597202 209900 597210
rect 203640 596788 204814 596798
rect 205094 596788 205678 596810
rect 203640 596764 205678 596788
rect 204372 596754 205678 596764
rect 205094 596718 205678 596754
rect 187315 596604 187316 596605
rect 187354 596604 187364 596608
rect 187316 596603 187317 596604
rect 184053 596592 184098 596603
rect 184711 596592 184756 596603
rect 185369 596592 185414 596603
rect 186027 596594 186072 596603
rect 184064 596358 184098 596592
rect 184109 596370 184110 596371
rect 184710 596370 184711 596371
rect 184110 596369 184111 596370
rect 184709 596369 184710 596370
rect 184722 596358 184756 596592
rect 184767 596370 184768 596371
rect 185368 596370 185369 596371
rect 184768 596369 184769 596370
rect 185367 596369 185368 596370
rect 185380 596358 185414 596592
rect 186012 596382 186092 596594
rect 186685 596592 186730 596603
rect 185425 596370 185426 596371
rect 185426 596369 185427 596370
rect 185888 596358 186346 596382
rect 186684 596370 186685 596371
rect 186683 596369 186684 596370
rect 186696 596358 186730 596592
rect 187342 596392 187400 596604
rect 186741 596370 186742 596371
rect 187324 596370 187400 596392
rect 186742 596369 186743 596370
rect 187304 596364 187315 596369
rect 187296 596358 187316 596364
rect 183950 596324 187316 596358
rect 166718 596051 166799 596098
rect 166858 596079 167810 596113
rect 170292 596079 173878 596113
rect 174859 596101 174866 596206
rect 174887 596129 174894 596206
rect 166991 596067 166992 596068
rect 166992 596066 166993 596067
rect 166731 596016 166744 596051
rect 166765 595908 166799 596051
rect 167004 595908 167038 596079
rect 167050 596067 167051 596068
rect 167649 596067 167650 596068
rect 167049 596066 167050 596067
rect 167650 596066 167651 596067
rect 167596 596046 167656 596048
rect 167662 595908 167696 596079
rect 167776 596048 167810 596079
rect 167702 596046 167868 596048
rect 167776 595908 167810 596046
rect 166418 594797 170042 595908
rect 170326 595455 170360 596079
rect 170440 595455 170474 596079
rect 170486 596067 170487 596068
rect 171085 596067 171086 596068
rect 170485 596066 170486 596067
rect 171086 596066 171087 596067
rect 170485 595467 170486 595468
rect 171086 595467 171087 595468
rect 170486 595466 170487 595467
rect 171085 595466 171086 595467
rect 171098 595455 171132 596079
rect 171144 596067 171145 596068
rect 171743 596067 171744 596068
rect 171143 596066 171144 596067
rect 171744 596066 171745 596067
rect 171134 595461 171138 595544
rect 171143 595467 171144 595468
rect 171744 595467 171745 595468
rect 171144 595466 171145 595467
rect 171743 595466 171744 595467
rect 171756 595455 171790 596079
rect 171802 596067 171803 596068
rect 172401 596067 172402 596068
rect 171801 596066 171802 596067
rect 172402 596066 172403 596067
rect 171801 595467 171802 595468
rect 172402 595467 172403 595468
rect 171802 595466 171803 595467
rect 172401 595466 172402 595467
rect 172414 595455 172448 596079
rect 172460 596067 172461 596068
rect 173059 596067 173060 596068
rect 172459 596066 172460 596067
rect 173060 596066 173061 596067
rect 172459 595467 172460 595468
rect 173060 595467 173061 595468
rect 172460 595466 172461 595467
rect 173059 595466 173060 595467
rect 173072 595455 173106 596079
rect 173118 596067 173119 596068
rect 173717 596067 173718 596068
rect 173117 596066 173118 596067
rect 173718 596066 173719 596067
rect 173117 595467 173118 595468
rect 173718 595467 173719 595468
rect 173118 595466 173119 595467
rect 173717 595466 173718 595467
rect 173730 595455 173764 596079
rect 173844 595455 173878 596079
rect 174859 595992 174866 596091
rect 174887 595992 174894 596063
rect 179526 595778 180358 595792
rect 179260 595740 179284 595762
rect 179238 595716 179284 595740
rect 183950 595700 183984 596324
rect 184064 595700 184098 596324
rect 184110 596312 184111 596313
rect 184709 596312 184710 596313
rect 184109 596311 184110 596312
rect 184710 596311 184711 596312
rect 184109 595712 184110 595713
rect 184710 595712 184711 595713
rect 184110 595711 184111 595712
rect 184709 595711 184710 595712
rect 184722 595700 184756 596324
rect 184768 596312 184769 596313
rect 185367 596312 185368 596313
rect 184767 596311 184768 596312
rect 185368 596311 185369 596312
rect 184767 595712 184768 595713
rect 185368 595712 185369 595713
rect 184768 595711 184769 595712
rect 185367 595711 185368 595712
rect 185380 595700 185414 596324
rect 185426 596312 185427 596313
rect 185425 596311 185426 596312
rect 185888 596290 186346 596324
rect 186683 596312 186684 596313
rect 186684 596311 186685 596312
rect 185425 595712 185426 595713
rect 186026 595712 186027 595713
rect 185426 595711 185427 595712
rect 186025 595711 186026 595712
rect 186038 595700 186072 596290
rect 186083 595712 186084 595713
rect 186684 595712 186685 595713
rect 186084 595711 186085 595712
rect 186683 595711 186684 595712
rect 186696 595700 186730 596324
rect 187296 596318 187316 596324
rect 186742 596312 186743 596313
rect 187324 596312 187344 596370
rect 187385 596355 187400 596370
rect 187385 596312 187400 596327
rect 186741 596311 186742 596312
rect 187324 596290 187400 596312
rect 186741 595712 186742 595713
rect 187342 595712 187400 596290
rect 186742 595711 186743 595712
rect 187304 595700 187315 595711
rect 183950 595666 187315 595700
rect 187348 595684 187372 595712
rect 187385 595697 187400 595712
rect 180302 595628 180414 595630
rect 170292 595421 173878 595455
rect 170326 594818 170360 595421
rect 170440 594979 170474 595421
rect 170486 595409 170487 595410
rect 171085 595409 171086 595410
rect 170485 595408 170486 595409
rect 171086 595408 171087 595409
rect 171098 594979 171132 595421
rect 171134 595322 171138 595415
rect 171144 595409 171145 595410
rect 171743 595409 171744 595410
rect 171143 595408 171144 595409
rect 171744 595408 171745 595409
rect 171756 595030 171790 595421
rect 171802 595409 171803 595410
rect 172401 595409 172402 595410
rect 171801 595408 171802 595409
rect 172402 595408 172403 595409
rect 172414 595030 172448 595421
rect 172460 595409 172461 595410
rect 173059 595409 173060 595410
rect 172459 595408 172460 595409
rect 173060 595408 173061 595409
rect 173072 595030 173106 595421
rect 173118 595409 173119 595410
rect 173717 595409 173718 595410
rect 173117 595408 173118 595409
rect 173718 595408 173719 595409
rect 173730 595030 173764 595421
rect 171756 594979 171801 595030
rect 172414 594979 172459 595030
rect 173072 594979 173117 595030
rect 173730 594979 173775 595030
rect 171070 594920 171117 594967
rect 171704 594920 173749 594967
rect 170502 594886 171117 594920
rect 171160 594886 171775 594920
rect 171818 594886 172433 594920
rect 172476 594886 173091 594920
rect 173134 594886 173749 594920
rect 170422 594818 173782 594831
rect 173844 594818 173878 595421
rect 183088 595232 183422 595410
rect 181622 595156 182542 595190
rect 181622 595042 181656 595156
rect 182366 595088 182404 595126
rect 181798 595076 182404 595088
rect 181782 595054 182404 595076
rect 181782 595042 182382 595054
rect 182508 595042 182542 595156
rect 182790 595148 183710 595182
rect 182790 595042 182824 595148
rect 183534 595080 183572 595118
rect 182966 595076 183572 595080
rect 182950 595046 183572 595076
rect 182950 595042 183550 595046
rect 183676 595042 183710 595148
rect 183950 595042 183984 595666
rect 184064 595042 184098 595666
rect 184110 595654 184111 595655
rect 184709 595654 184710 595655
rect 184109 595653 184110 595654
rect 184710 595653 184711 595654
rect 184109 595054 184110 595055
rect 184710 595054 184711 595055
rect 184110 595053 184111 595054
rect 184709 595053 184710 595054
rect 184722 595042 184756 595666
rect 184768 595654 184769 595655
rect 185367 595654 185368 595655
rect 184767 595653 184768 595654
rect 185368 595653 185369 595654
rect 184767 595054 184768 595055
rect 185368 595054 185369 595055
rect 184768 595053 184769 595054
rect 185367 595053 185368 595054
rect 185380 595042 185414 595666
rect 185426 595654 185427 595655
rect 186025 595654 186026 595655
rect 185425 595653 185426 595654
rect 186026 595653 186027 595654
rect 185425 595054 185426 595055
rect 186026 595054 186027 595055
rect 185426 595053 185427 595054
rect 186025 595053 186026 595054
rect 186038 595042 186072 595666
rect 186084 595654 186085 595655
rect 186683 595654 186684 595655
rect 186083 595653 186084 595654
rect 186684 595653 186685 595654
rect 186083 595054 186084 595055
rect 186684 595054 186685 595055
rect 186084 595053 186085 595054
rect 186683 595053 186684 595054
rect 186696 595042 186730 595666
rect 186742 595654 186743 595655
rect 187385 595654 187400 595669
rect 186741 595653 186742 595654
rect 186741 595054 186742 595055
rect 187342 595054 187400 595654
rect 186742 595053 186743 595054
rect 187304 595042 187315 595053
rect 179328 595008 187315 595042
rect 187385 595039 187400 595054
rect 170326 594797 173878 594818
rect 174855 594797 174864 594936
rect 174893 594825 174902 594974
rect 180576 594928 180958 595008
rect 181622 594928 181656 595008
rect 181736 594970 181770 595004
rect 182394 594970 182428 595004
rect 181736 594928 181770 594962
rect 182394 594928 182428 594962
rect 182508 594928 182542 595008
rect 182790 594928 182824 595008
rect 182904 594936 182938 594996
rect 182904 594928 183540 594936
rect 183562 594928 183596 594996
rect 183676 594928 183710 595008
rect 183950 594928 183984 595008
rect 184064 594928 184098 595008
rect 184722 594928 184756 595008
rect 185380 594928 185414 595008
rect 186038 594928 186072 595008
rect 186696 594928 186730 595008
rect 187456 594990 187502 596682
rect 204876 596246 204910 596702
rect 208646 596544 208702 596546
rect 209844 596544 209900 596546
rect 208646 596488 208702 596490
rect 209844 596488 209900 596490
rect 205014 596310 205034 596352
rect 205014 596246 205054 596310
rect 205058 596246 205082 596282
rect 205094 596246 205680 596282
rect 187354 594928 187388 594962
rect 179238 594894 187422 594928
rect 180576 594832 180958 594894
rect 180542 594806 180958 594832
rect 166418 594763 174864 594797
rect 180494 594798 180958 594806
rect 166418 593955 170042 594763
rect 174855 594564 174864 594763
rect 174893 594526 174902 594735
rect 179798 594556 179816 594778
rect 179826 594556 179844 594750
rect 180494 594720 180576 594798
rect 181622 594612 181656 594894
rect 182508 594612 182542 594894
rect 182790 594612 182824 594894
rect 182904 594798 183540 594894
rect 183562 594798 183596 594894
rect 182904 594612 183620 594798
rect 183676 594612 183710 594894
rect 181586 594600 182578 594612
rect 179324 594462 179866 594490
rect 179284 594422 179832 594456
rect 179250 594360 179270 594394
rect 173164 594166 174516 594182
rect 179284 594140 179318 594422
rect 179646 594342 179657 594353
rect 179348 594298 179420 594336
rect 179470 594308 179657 594342
rect 179658 594298 179730 594336
rect 179386 594264 179420 594298
rect 179646 594254 179657 594265
rect 179696 594264 179730 594298
rect 179470 594220 179657 594254
rect 179798 594140 179832 594422
rect 179882 594408 180078 594510
rect 179880 594168 180078 594408
rect 179284 594106 179832 594140
rect 179882 594048 180078 594168
rect 180276 594048 180520 594510
rect 165024 592523 165070 592535
rect 166312 592495 166318 592584
rect 166340 592538 166374 592584
rect 166340 592535 166380 592538
rect 166340 592523 166386 592535
rect 166418 592472 167846 593955
rect 167872 592498 167930 592526
rect 168530 592498 168588 592526
rect 169188 592498 169246 592526
rect 169846 592498 169904 592526
rect 167884 592494 167918 592498
rect 168542 592494 168576 592498
rect 169200 592494 169234 592498
rect 169858 592494 169892 592498
rect 169972 592472 170006 593955
rect 171395 593251 171540 593350
rect 181622 593338 181656 594600
rect 182508 593338 182542 594600
rect 182754 594594 183746 594612
rect 182790 594556 182824 594594
rect 182904 594564 183620 594594
rect 182904 594556 182938 594564
rect 183562 594556 183596 594564
rect 183676 594556 183710 594594
rect 182698 594538 183802 594556
rect 182790 593330 182824 594538
rect 182904 593420 182938 594538
rect 183562 593420 183596 594538
rect 183676 593330 183710 594538
rect 183950 593326 183984 594894
rect 184754 593404 184762 594496
rect 185474 593756 185476 594496
rect 185474 593372 185500 593428
rect 185430 593348 185476 593372
rect 187468 593326 187502 594990
rect 204278 596212 205680 596246
rect 204278 594702 204312 596212
rect 204727 596132 204839 596144
rect 204876 596132 204910 596212
rect 204473 596129 204839 596132
rect 204333 596110 204414 596117
rect 204333 596086 204448 596110
rect 204473 596098 204824 596129
rect 204842 596098 204910 596132
rect 204727 596086 204824 596098
rect 204333 596082 204414 596086
rect 204333 596070 204420 596082
rect 204374 596058 204420 596070
rect 204774 596062 204808 596086
rect 204380 596039 204414 596058
rect 204768 596042 204814 596062
rect 204333 596038 204414 596039
rect 204333 596026 204461 596038
rect 204715 596026 204726 596037
rect 204333 595992 204726 596026
rect 204740 596014 204842 596034
rect 204364 595980 204461 595992
rect 204380 595502 204414 595980
rect 204727 595964 204808 596011
rect 204774 595487 204808 595964
rect 204727 595486 204808 595487
rect 204727 595474 204824 595486
rect 204876 595474 204910 596098
rect 205014 595744 205054 596212
rect 205058 595744 205082 596212
rect 205094 595842 205680 596212
rect 208646 595886 208702 595888
rect 209844 595886 209900 595888
rect 205094 595818 206122 595842
rect 208646 595830 208702 595832
rect 209844 595830 209900 595832
rect 205490 595804 206122 595818
rect 205524 595744 205542 595800
rect 205550 595744 206062 595782
rect 205014 595690 205034 595744
rect 205524 595638 205542 595690
rect 205552 595666 205570 595690
rect 204333 595452 204414 595459
rect 204333 595434 204448 595452
rect 204473 595440 204824 595474
rect 204842 595440 204910 595474
rect 204333 595424 204414 595434
rect 204333 595412 204420 595424
rect 204374 595406 204420 595412
rect 204466 595410 204642 595432
rect 204727 595428 204824 595440
rect 204774 595408 204808 595428
rect 204380 595381 204414 595406
rect 204333 595380 204414 595381
rect 204416 595380 204420 595406
rect 204444 595382 204670 595404
rect 204768 595384 204814 595408
rect 204444 595380 204448 595382
rect 204333 595368 204461 595380
rect 204715 595368 204726 595379
rect 204333 595334 204726 595368
rect 204740 595356 204842 595380
rect 204364 595322 204461 595334
rect 204380 594844 204414 595322
rect 204727 595306 204808 595353
rect 204774 594829 204808 595306
rect 204727 594828 204808 594829
rect 204727 594816 204824 594828
rect 204876 594816 204910 595440
rect 204473 594785 204824 594816
rect 204473 594782 204839 594785
rect 204842 594782 204910 594816
rect 204727 594770 204839 594782
rect 204774 594738 204808 594740
rect 204774 594722 204808 594736
rect 204876 594702 204910 594782
rect 205094 594702 205680 595620
rect 204278 594668 205680 594702
rect 208646 594670 208702 594672
rect 209844 594670 209900 594672
rect 204876 594658 204910 594668
rect 205094 594632 205680 594668
rect 207690 594618 208614 594644
rect 208646 594614 208702 594616
rect 209844 594614 209900 594616
rect 207724 594584 208614 594610
rect 204222 594186 204870 594196
rect 205086 594142 207106 594178
rect 204372 594140 207106 594142
rect 204332 594118 207106 594140
rect 204276 594108 207106 594118
rect 204276 594080 204310 594108
rect 204332 594080 204725 594106
rect 204242 594074 204725 594080
rect 204242 594072 204344 594074
rect 171649 592888 171794 593251
rect 179122 593250 180042 593274
rect 180312 593250 180362 593274
rect 180387 593251 181232 593269
rect 181622 593251 182542 593269
rect 182790 593268 182824 593269
rect 183676 593268 183710 593269
rect 182790 593251 183710 593268
rect 183950 593264 183984 593269
rect 187468 593264 187502 593274
rect 183950 593251 184046 593264
rect 180387 593250 181268 593251
rect 179088 593216 180076 593220
rect 180278 593216 180308 593220
rect 180405 593214 181268 593250
rect 181586 593206 182578 593251
rect 182754 593198 183746 593251
rect 183914 593230 184046 593251
rect 185458 593230 187502 593264
rect 183914 593194 184029 593230
rect 185512 593196 187536 593220
rect 173828 593124 173906 593147
rect 173823 593096 173906 593119
rect 171649 592472 175070 592508
rect 166418 592460 175070 592472
rect 177494 592470 177498 593074
rect 177522 593034 177568 593046
rect 177522 593022 177562 593034
rect 179062 593030 180344 593066
rect 180441 593030 180475 593119
rect 177522 592470 177554 593022
rect 179062 592996 181334 593030
rect 166418 592449 167872 592460
rect 167930 592449 168530 592460
rect 168588 592449 169188 592460
rect 169246 592449 175070 592460
rect 166418 592438 167883 592449
rect 167919 592438 168541 592449
rect 168577 592438 169199 592449
rect 169235 592438 175070 592449
rect 166418 592422 167846 592438
rect 169972 592428 170006 592438
rect 169554 592426 170042 592428
rect 166418 592420 167868 592422
rect 167934 592420 168526 592422
rect 169972 592420 170006 592426
rect 166418 592394 167846 592420
rect 166418 592392 167896 592394
rect 167906 592392 168554 592394
rect 166418 592358 167846 592392
rect 169554 592370 170098 592400
rect 169972 592358 170006 592370
rect 166418 592336 170006 592358
rect 166418 592324 170482 592336
rect 166418 592312 168030 592324
rect 168440 592318 170482 592324
rect 168440 592312 168558 592318
rect 166418 592304 168558 592312
rect 157844 591810 158880 591818
rect 158800 591730 158880 591738
rect 161190 591138 161198 592280
rect 166686 590538 166720 592304
rect 167156 592286 168558 592304
rect 168030 592280 168440 592284
rect 167128 592258 168586 592280
rect 167162 591070 168564 591084
rect 171649 588884 175070 592438
rect 173340 588774 173552 588884
rect 176870 585058 176904 590538
rect 177494 588926 177498 591366
rect 177522 590538 177554 591366
rect 177654 591310 177676 592526
rect 178844 592056 178878 592076
rect 178920 592056 178940 592452
rect 178844 592028 178982 592056
rect 178820 591800 179020 592028
rect 177522 588870 177562 590538
rect 177528 585058 177562 588870
rect 178186 585058 178220 590538
rect 178844 585058 178878 591800
rect 178920 591760 178940 591782
rect 179062 591698 180344 592996
rect 180441 591698 180475 592996
rect 180555 592990 180589 592996
rect 180500 592894 180509 592928
rect 180543 592894 180547 592975
rect 180549 592944 180589 592990
rect 180549 592934 180601 592944
rect 180555 592928 180601 592934
rect 181158 592928 181205 592975
rect 180555 592894 181205 592928
rect 180555 592847 180601 592894
rect 180492 592564 180518 592836
rect 180555 592835 180589 592847
rect 181175 592835 181201 592846
rect 181213 592835 181247 592996
rect 180528 591859 180589 592835
rect 181186 592204 181247 592835
rect 181186 592050 181266 592204
rect 181172 591862 181266 592050
rect 181186 591859 181266 591862
rect 180555 591847 180589 591859
rect 181196 591847 181266 591859
rect 180500 591766 180509 591800
rect 180543 591766 180547 591847
rect 180555 591800 180601 591847
rect 181158 591800 181266 591847
rect 180555 591766 181266 591800
rect 180555 591760 180601 591766
rect 180549 591750 180601 591760
rect 180549 591704 180589 591750
rect 181196 591748 181266 591766
rect 180555 591698 180589 591704
rect 181213 591698 181247 591748
rect 181300 591698 181334 592996
rect 179062 591664 181334 591698
rect 181676 592990 183891 593024
rect 181676 591692 181710 592990
rect 181871 592938 181918 592969
rect 181859 592922 181918 592938
rect 182420 592922 182467 592969
rect 182529 592938 182576 592969
rect 182517 592922 182576 592938
rect 183078 592922 183125 592969
rect 183187 592938 183234 592969
rect 183175 592922 183234 592938
rect 183736 592922 183783 592969
rect 181852 592888 182467 592922
rect 182510 592888 183125 592922
rect 183168 592897 183783 592922
rect 183156 592888 183783 592897
rect 181756 592834 181778 592869
rect 181859 592841 181917 592888
rect 181784 592840 181806 592841
rect 181779 592829 181824 592840
rect 181790 592538 181824 592829
rect 181837 592538 181858 592834
rect 181756 591813 181778 592538
rect 181784 591853 181824 592538
rect 181865 592510 181905 592841
rect 182414 592840 182440 592869
rect 182517 592841 182575 592888
rect 183156 592882 183234 592888
rect 183175 592841 183234 592882
rect 182442 592840 182488 592841
rect 182414 592829 182488 592840
rect 182414 592788 182440 592829
rect 181784 591841 181806 591853
rect 181871 591841 181905 592510
rect 182386 592056 182440 592788
rect 182442 592732 182488 592829
rect 182442 592420 182482 592732
rect 182529 592420 182563 592841
rect 183125 592840 183146 592841
rect 183181 592840 183234 592841
rect 183095 592829 183178 592840
rect 183106 592558 183178 592829
rect 183106 592420 183146 592558
rect 183181 592420 183221 592840
rect 183753 592829 183798 592840
rect 183764 592420 183798 592829
rect 183839 592702 183860 592897
rect 182442 592056 182493 592420
rect 182448 591853 182493 592056
rect 182508 591848 182516 592064
rect 182386 591841 182440 591846
rect 182442 591841 182468 591846
rect 182529 591841 182574 592420
rect 183106 591853 183151 592420
rect 183125 591841 183146 591853
rect 183181 591841 183232 592420
rect 183764 591853 183809 592420
rect 181859 591794 181918 591841
rect 182386 591794 183783 591841
rect 181852 591760 182467 591794
rect 182510 591760 183125 591794
rect 183156 591785 183783 591794
rect 181859 591744 181917 591760
rect 182424 591732 182440 591760
rect 182517 591744 182575 591760
rect 183156 591754 183166 591785
rect 183168 591760 183783 591785
rect 183175 591744 183233 591760
rect 183845 591692 183850 591726
rect 183878 591692 183891 592990
rect 179062 591628 180344 591664
rect 180084 590822 180344 590858
rect 180441 590822 180475 591664
rect 181676 591658 183891 591692
rect 183959 591318 183993 593119
rect 183632 591284 185078 591318
rect 180084 590788 183014 590822
rect 180084 589990 180344 590788
rect 180441 589990 180475 590788
rect 180555 590751 180602 590767
rect 180543 590720 180602 590751
rect 180864 590720 180911 590767
rect 181213 590736 181260 590767
rect 181201 590720 181260 590736
rect 181522 590720 181569 590767
rect 181871 590736 181918 590767
rect 181859 590720 181918 590736
rect 182180 590720 182227 590767
rect 182529 590736 182576 590767
rect 182517 590720 182576 590736
rect 182838 590720 182885 590767
rect 180543 590686 180911 590720
rect 180954 590686 181569 590720
rect 181612 590686 182227 590720
rect 182270 590686 182885 590720
rect 180543 590639 180601 590686
rect 181201 590639 181259 590686
rect 181859 590639 181917 590686
rect 182517 590639 182575 590686
rect 180555 590139 180589 590639
rect 180881 590627 180926 590638
rect 180892 590151 180926 590627
rect 181213 590139 181247 590639
rect 181539 590627 181584 590638
rect 181550 590151 181584 590627
rect 181871 590139 181905 590639
rect 182197 590627 182242 590638
rect 182208 590151 182242 590627
rect 182529 590139 182563 590639
rect 182855 590627 182900 590638
rect 182866 590151 182900 590627
rect 180543 590092 180602 590139
rect 180864 590092 180911 590139
rect 181201 590092 181260 590139
rect 181522 590092 181569 590139
rect 181859 590092 181918 590139
rect 182180 590092 182227 590139
rect 182517 590092 182576 590139
rect 182838 590092 182885 590139
rect 180543 590058 180911 590092
rect 180954 590058 181569 590092
rect 181612 590058 182227 590092
rect 182270 590058 182885 590092
rect 180543 590042 180601 590058
rect 181201 590042 181259 590058
rect 181859 590042 181917 590058
rect 182517 590042 182575 590058
rect 180543 590027 180558 590042
rect 182980 589990 183014 590788
rect 180084 589956 183014 589990
rect 183632 589986 183666 591284
rect 183761 591216 183891 591263
rect 183808 591182 183891 591216
rect 183833 591135 183891 591182
rect 183735 591123 183791 591134
rect 183746 591102 183791 591123
rect 183845 591102 183890 591135
rect 183746 590147 183780 591102
rect 183845 590135 183879 591102
rect 183833 590088 183891 590135
rect 183808 590054 183891 590088
rect 183833 590038 183891 590054
rect 183876 590023 183891 590038
rect 183959 589986 183993 591284
rect 185518 591004 185564 591020
rect 183632 589980 185078 589986
rect 180084 589920 180344 589956
rect 180441 584945 180475 589956
rect 183632 589952 185246 589980
rect 180728 586180 181118 586214
rect 180728 585682 180762 586180
rect 180942 586112 180989 586159
rect 180904 586078 180989 586112
rect 180831 586019 180876 586030
rect 180959 586019 181004 586030
rect 180842 585843 180876 586019
rect 180970 585843 181004 586019
rect 180942 585784 180989 585831
rect 180904 585750 180989 585784
rect 181084 585682 181118 586180
rect 180728 585648 181118 585682
rect 180710 584978 181132 585598
rect 183959 584945 183993 589952
rect 184380 589916 185246 589952
rect 185682 589918 187332 591356
rect 187676 591348 187696 592452
rect 187600 589490 187634 590538
rect 187786 589916 189100 593256
rect 204276 592018 204310 594072
rect 204431 594038 204714 594062
rect 204768 594044 204802 594062
rect 204721 594034 204833 594040
rect 204459 594025 204833 594034
rect 204870 594028 204904 594108
rect 204331 593966 204412 594013
rect 204459 594010 204818 594025
rect 204471 593994 204818 594010
rect 204836 593994 204904 594028
rect 204721 593982 204818 593994
rect 204378 593461 204412 593966
rect 204768 593476 204802 593982
rect 204331 593460 204412 593461
rect 204331 593448 204459 593460
rect 204709 593448 204720 593459
rect 204331 593414 204720 593448
rect 204362 593408 204678 593414
rect 204362 593402 204459 593408
rect 204378 593398 204412 593402
rect 204464 593380 204650 593398
rect 204721 593386 204802 593433
rect 204768 593383 204802 593386
rect 204721 593382 204802 593383
rect 204721 593370 204818 593382
rect 204870 593370 204904 593994
rect 204331 593308 204412 593355
rect 204471 593336 204818 593370
rect 204836 593336 204904 593370
rect 204721 593324 204818 593336
rect 204378 592803 204412 593308
rect 204768 592818 204802 593324
rect 204331 592802 204412 592803
rect 204331 592790 204459 592802
rect 204709 592790 204720 592801
rect 204331 592756 204720 592790
rect 204362 592744 204459 592756
rect 204378 592740 204418 592744
rect 204410 592728 204418 592740
rect 204438 592718 204446 592744
rect 204721 592728 204802 592775
rect 204768 592725 204802 592728
rect 204721 592724 204802 592725
rect 204721 592712 204818 592724
rect 204870 592712 204904 593336
rect 205086 594002 207106 594108
rect 205086 593988 207276 594002
rect 205086 593974 207106 593988
rect 205086 593960 207248 593974
rect 205086 593318 207106 593960
rect 204331 592650 204412 592697
rect 204471 592678 204818 592712
rect 204836 592678 204904 592712
rect 204721 592666 204818 592678
rect 204378 592145 204412 592650
rect 204768 592160 204802 592666
rect 204331 592144 204412 592145
rect 204331 592132 204459 592144
rect 204709 592132 204720 592143
rect 204331 592098 204720 592132
rect 204347 592092 204698 592098
rect 204347 592088 204459 592092
rect 204347 592086 204670 592088
rect 204448 592064 204670 592086
rect 204344 592018 204446 592026
rect 204471 592020 204842 592052
rect 204870 592018 204904 592678
rect 205078 592712 207098 593142
rect 205078 592678 208447 592712
rect 205078 592150 207098 592678
rect 203634 591984 204904 592018
rect 204276 590686 204310 591984
rect 205074 590554 208678 591982
rect 205212 590528 205246 590554
rect 205308 590532 205636 590554
rect 187732 589746 187754 589750
rect 187704 589718 187726 589722
rect 187704 589492 187728 589718
rect 187704 589490 187726 589492
rect 187732 589490 187756 589746
rect 187410 589478 187756 589490
rect 187600 585058 187634 589478
rect 187732 589464 187756 589478
rect 187732 589460 187754 589464
<< metal2 >>
rect 524 -800 636 480
rect 1706 -800 1818 480
rect 2888 -800 3000 480
rect 4070 -800 4182 480
rect 5252 -800 5364 480
rect 6434 -800 6546 480
rect 7616 -800 7728 480
rect 8798 -800 8910 480
rect 9980 -800 10092 480
rect 11162 -800 11274 480
rect 12344 -800 12456 480
rect 13526 -800 13638 480
rect 14708 -800 14820 480
rect 15890 -800 16002 480
rect 17072 -800 17184 480
rect 18254 -800 18366 480
rect 19436 -800 19548 480
rect 20618 -800 20730 480
rect 21800 -800 21912 480
rect 22982 -800 23094 480
rect 24164 -800 24276 480
rect 25346 -800 25458 480
rect 26528 -800 26640 480
rect 27710 -800 27822 480
rect 28892 -800 29004 480
rect 30074 -800 30186 480
rect 31256 -800 31368 480
rect 32438 -800 32550 480
rect 33620 -800 33732 480
rect 34802 -800 34914 480
rect 35984 -800 36096 480
rect 37166 -800 37278 480
rect 38348 -800 38460 480
rect 39530 -800 39642 480
rect 40712 -800 40824 480
rect 41894 -800 42006 480
rect 43076 -800 43188 480
rect 44258 -800 44370 480
rect 45440 -800 45552 480
rect 46622 -800 46734 480
rect 47804 -800 47916 480
rect 48986 -800 49098 480
rect 50168 -800 50280 480
rect 51350 -800 51462 480
rect 52532 -800 52644 480
rect 53714 -800 53826 480
rect 54896 -800 55008 480
rect 56078 -800 56190 480
rect 57260 -800 57372 480
rect 58442 -800 58554 480
rect 59624 -800 59736 480
rect 60806 -800 60918 480
rect 61988 -800 62100 480
rect 63170 -800 63282 480
rect 64352 -800 64464 480
rect 65534 -800 65646 480
rect 66716 -800 66828 480
rect 67898 -800 68010 480
rect 69080 -800 69192 480
rect 70262 -800 70374 480
rect 71444 -800 71556 480
rect 72626 -800 72738 480
rect 73808 -800 73920 480
rect 74990 -800 75102 480
rect 76172 -800 76284 480
rect 77354 -800 77466 480
rect 78536 -800 78648 480
rect 79718 -800 79830 480
rect 80900 -800 81012 480
rect 82082 -800 82194 480
rect 83264 -800 83376 480
rect 84446 -800 84558 480
rect 85628 -800 85740 480
rect 86810 -800 86922 480
rect 87992 -800 88104 480
rect 89174 -800 89286 480
rect 90356 -800 90468 480
rect 91538 -800 91650 480
rect 92720 -800 92832 480
rect 93902 -800 94014 480
rect 95084 -800 95196 480
rect 96266 -800 96378 480
rect 97448 -800 97560 480
rect 98630 -800 98742 480
rect 99812 -800 99924 480
rect 100994 -800 101106 480
rect 102176 -800 102288 480
rect 103358 -800 103470 480
rect 104540 -800 104652 480
rect 105722 -800 105834 480
rect 106904 -800 107016 480
rect 108086 -800 108198 480
rect 109268 -800 109380 480
rect 110450 -800 110562 480
rect 111632 -800 111744 480
rect 112814 -800 112926 480
rect 113996 -800 114108 480
rect 115178 -800 115290 480
rect 116360 -800 116472 480
rect 117542 -800 117654 480
rect 118724 -800 118836 480
rect 119906 -800 120018 480
rect 121088 -800 121200 480
rect 122270 -800 122382 480
rect 123452 -800 123564 480
rect 124634 -800 124746 480
rect 125816 -800 125928 480
rect 126998 -800 127110 480
rect 128180 -800 128292 480
rect 129362 -800 129474 480
rect 130544 -800 130656 480
rect 131726 -800 131838 480
rect 132908 -800 133020 480
rect 134090 -800 134202 480
rect 135272 -800 135384 480
rect 136454 -800 136566 480
rect 137636 -800 137748 480
rect 138818 -800 138930 480
rect 140000 -800 140112 480
rect 141182 -800 141294 480
rect 142364 -800 142476 480
rect 143546 -800 143658 480
rect 144728 -800 144840 480
rect 145910 -800 146022 480
rect 147092 -800 147204 480
rect 148274 -800 148386 480
rect 149456 -800 149568 480
rect 150638 -800 150750 480
rect 151820 -800 151932 480
rect 153002 -800 153114 480
rect 154184 -800 154296 480
rect 155366 -800 155478 480
rect 156548 -800 156660 480
rect 157730 -800 157842 480
rect 158912 -800 159024 480
rect 160094 -800 160206 480
rect 161276 -800 161388 480
rect 162458 -800 162570 480
rect 163640 -800 163752 480
rect 164822 -800 164934 480
rect 166004 -800 166116 480
rect 167186 -800 167298 480
rect 168368 -800 168480 480
rect 169550 -800 169662 480
rect 170732 -800 170844 480
rect 171914 -800 172026 480
rect 173096 -800 173208 480
rect 174278 -800 174390 480
rect 175460 -800 175572 480
rect 176642 -800 176754 480
rect 177824 -800 177936 480
rect 179006 -800 179118 480
rect 180188 -800 180300 480
rect 181370 -800 181482 480
rect 182552 -800 182664 480
rect 183734 -800 183846 480
rect 184916 -800 185028 480
rect 186098 -800 186210 480
rect 187280 -800 187392 480
rect 188462 -800 188574 480
rect 189644 -800 189756 480
rect 190826 -800 190938 480
rect 192008 -800 192120 480
rect 193190 -800 193302 480
rect 194372 -800 194484 480
rect 195554 -800 195666 480
rect 196736 -800 196848 480
rect 197918 -800 198030 480
rect 199100 -800 199212 480
rect 200282 -800 200394 480
rect 201464 -800 201576 480
rect 202646 -800 202758 480
rect 203828 -800 203940 480
rect 205010 -800 205122 480
rect 206192 -800 206304 480
rect 207374 -800 207486 480
rect 208556 -800 208668 480
rect 209738 -800 209850 480
rect 210920 -800 211032 480
rect 212102 -800 212214 480
rect 213284 -800 213396 480
rect 214466 -800 214578 480
rect 215648 -800 215760 480
rect 216830 -800 216942 480
rect 218012 -800 218124 480
rect 219194 -800 219306 480
rect 220376 -800 220488 480
rect 221558 -800 221670 480
rect 222740 -800 222852 480
rect 223922 -800 224034 480
rect 225104 -800 225216 480
rect 226286 -800 226398 480
rect 227468 -800 227580 480
rect 228650 -800 228762 480
rect 229832 -800 229944 480
rect 231014 -800 231126 480
rect 232196 -800 232308 480
rect 233378 -800 233490 480
rect 234560 -800 234672 480
rect 235742 -800 235854 480
rect 236924 -800 237036 480
rect 238106 -800 238218 480
rect 239288 -800 239400 480
rect 240470 -800 240582 480
rect 241652 -800 241764 480
rect 242834 -800 242946 480
rect 244016 -800 244128 480
rect 245198 -800 245310 480
rect 246380 -800 246492 480
rect 247562 -800 247674 480
rect 248744 -800 248856 480
rect 249926 -800 250038 480
rect 251108 -800 251220 480
rect 252290 -800 252402 480
rect 253472 -800 253584 480
rect 254654 -800 254766 480
rect 255836 -800 255948 480
rect 257018 -800 257130 480
rect 258200 -800 258312 480
rect 259382 -800 259494 480
rect 260564 -800 260676 480
rect 261746 -800 261858 480
rect 262928 -800 263040 480
rect 264110 -800 264222 480
rect 265292 -800 265404 480
rect 266474 -800 266586 480
rect 267656 -800 267768 480
rect 268838 -800 268950 480
rect 270020 -800 270132 480
rect 271202 -800 271314 480
rect 272384 -800 272496 480
rect 273566 -800 273678 480
rect 274748 -800 274860 480
rect 275930 -800 276042 480
rect 277112 -800 277224 480
rect 278294 -800 278406 480
rect 279476 -800 279588 480
rect 280658 -800 280770 480
rect 281840 -800 281952 480
rect 283022 -800 283134 480
rect 284204 -800 284316 480
rect 285386 -800 285498 480
rect 286568 -800 286680 480
rect 287750 -800 287862 480
rect 288932 -800 289044 480
rect 290114 -800 290226 480
rect 291296 -800 291408 480
rect 292478 -800 292590 480
rect 293660 -800 293772 480
rect 294842 -800 294954 480
rect 296024 -800 296136 480
rect 297206 -800 297318 480
rect 298388 -800 298500 480
rect 299570 -800 299682 480
rect 300752 -800 300864 480
rect 301934 -800 302046 480
rect 303116 -800 303228 480
rect 304298 -800 304410 480
rect 305480 -800 305592 480
rect 306662 -800 306774 480
rect 307844 -800 307956 480
rect 309026 -800 309138 480
rect 310208 -800 310320 480
rect 311390 -800 311502 480
rect 312572 -800 312684 480
rect 313754 -800 313866 480
rect 314936 -800 315048 480
rect 316118 -800 316230 480
rect 317300 -800 317412 480
rect 318482 -800 318594 480
rect 319664 -800 319776 480
rect 320846 -800 320958 480
rect 322028 -800 322140 480
rect 323210 -800 323322 480
rect 324392 -800 324504 480
rect 325574 -800 325686 480
rect 326756 -800 326868 480
rect 327938 -800 328050 480
rect 329120 -800 329232 480
rect 330302 -800 330414 480
rect 331484 -800 331596 480
rect 332666 -800 332778 480
rect 333848 -800 333960 480
rect 335030 -800 335142 480
rect 336212 -800 336324 480
rect 337394 -800 337506 480
rect 338576 -800 338688 480
rect 339758 -800 339870 480
rect 340940 -800 341052 480
rect 342122 -800 342234 480
rect 343304 -800 343416 480
rect 344486 -800 344598 480
rect 345668 -800 345780 480
rect 346850 -800 346962 480
rect 348032 -800 348144 480
rect 349214 -800 349326 480
rect 350396 -800 350508 480
rect 351578 -800 351690 480
rect 352760 -800 352872 480
rect 353942 -800 354054 480
rect 355124 -800 355236 480
rect 356306 -800 356418 480
rect 357488 -800 357600 480
rect 358670 -800 358782 480
rect 359852 -800 359964 480
rect 361034 -800 361146 480
rect 362216 -800 362328 480
rect 363398 -800 363510 480
rect 364580 -800 364692 480
rect 365762 -800 365874 480
rect 366944 -800 367056 480
rect 368126 -800 368238 480
rect 369308 -800 369420 480
rect 370490 -800 370602 480
rect 371672 -800 371784 480
rect 372854 -800 372966 480
rect 374036 -800 374148 480
rect 375218 -800 375330 480
rect 376400 -800 376512 480
rect 377582 -800 377694 480
rect 378764 -800 378876 480
rect 379946 -800 380058 480
rect 381128 -800 381240 480
rect 382310 -800 382422 480
rect 383492 -800 383604 480
rect 384674 -800 384786 480
rect 385856 -800 385968 480
rect 387038 -800 387150 480
rect 388220 -800 388332 480
rect 389402 -800 389514 480
rect 390584 -800 390696 480
rect 391766 -800 391878 480
rect 392948 -800 393060 480
rect 394130 -800 394242 480
rect 395312 -800 395424 480
rect 396494 -800 396606 480
rect 397676 -800 397788 480
rect 398858 -800 398970 480
rect 400040 -800 400152 480
rect 401222 -800 401334 480
rect 402404 -800 402516 480
rect 403586 -800 403698 480
rect 404768 -800 404880 480
rect 405950 -800 406062 480
rect 407132 -800 407244 480
rect 408314 -800 408426 480
rect 409496 -800 409608 480
rect 410678 -800 410790 480
rect 411860 -800 411972 480
rect 413042 -800 413154 480
rect 414224 -800 414336 480
rect 415406 -800 415518 480
rect 416588 -800 416700 480
rect 417770 -800 417882 480
rect 418952 -800 419064 480
rect 420134 -800 420246 480
rect 421316 -800 421428 480
rect 422498 -800 422610 480
rect 423680 -800 423792 480
rect 424862 -800 424974 480
rect 426044 -800 426156 480
rect 427226 -800 427338 480
rect 428408 -800 428520 480
rect 429590 -800 429702 480
rect 430772 -800 430884 480
rect 431954 -800 432066 480
rect 433136 -800 433248 480
rect 434318 -800 434430 480
rect 435500 -800 435612 480
rect 436682 -800 436794 480
rect 437864 -800 437976 480
rect 439046 -800 439158 480
rect 440228 -800 440340 480
rect 441410 -800 441522 480
rect 442592 -800 442704 480
rect 443774 -800 443886 480
rect 444956 -800 445068 480
rect 446138 -800 446250 480
rect 447320 -800 447432 480
rect 448502 -800 448614 480
rect 449684 -800 449796 480
rect 450866 -800 450978 480
rect 452048 -800 452160 480
rect 453230 -800 453342 480
rect 454412 -800 454524 480
rect 455594 -800 455706 480
rect 456776 -800 456888 480
rect 457958 -800 458070 480
rect 459140 -800 459252 480
rect 460322 -800 460434 480
rect 461504 -800 461616 480
rect 462686 -800 462798 480
rect 463868 -800 463980 480
rect 465050 -800 465162 480
rect 466232 -800 466344 480
rect 467414 -800 467526 480
rect 468596 -800 468708 480
rect 469778 -800 469890 480
rect 470960 -800 471072 480
rect 472142 -800 472254 480
rect 473324 -800 473436 480
rect 474506 -800 474618 480
rect 475688 -800 475800 480
rect 476870 -800 476982 480
rect 478052 -800 478164 480
rect 479234 -800 479346 480
rect 480416 -800 480528 480
rect 481598 -800 481710 480
rect 482780 -800 482892 480
rect 483962 -800 484074 480
rect 485144 -800 485256 480
rect 486326 -800 486438 480
rect 487508 -800 487620 480
rect 488690 -800 488802 480
rect 489872 -800 489984 480
rect 491054 -800 491166 480
rect 492236 -800 492348 480
rect 493418 -800 493530 480
rect 494600 -800 494712 480
rect 495782 -800 495894 480
rect 496964 -800 497076 480
rect 498146 -800 498258 480
rect 499328 -800 499440 480
rect 500510 -800 500622 480
rect 501692 -800 501804 480
rect 502874 -800 502986 480
rect 504056 -800 504168 480
rect 505238 -800 505350 480
rect 506420 -800 506532 480
rect 507602 -800 507714 480
rect 508784 -800 508896 480
rect 509966 -800 510078 480
rect 511148 -800 511260 480
rect 512330 -800 512442 480
rect 513512 -800 513624 480
rect 514694 -800 514806 480
rect 515876 -800 515988 480
rect 517058 -800 517170 480
rect 518240 -800 518352 480
rect 519422 -800 519534 480
rect 520604 -800 520716 480
rect 521786 -800 521898 480
rect 522968 -800 523080 480
rect 524150 -800 524262 480
rect 525332 -800 525444 480
rect 526514 -800 526626 480
rect 527696 -800 527808 480
rect 528878 -800 528990 480
rect 530060 -800 530172 480
rect 531242 -800 531354 480
rect 532424 -800 532536 480
rect 533606 -800 533718 480
rect 534788 -800 534900 480
rect 535970 -800 536082 480
rect 537152 -800 537264 480
rect 538334 -800 538446 480
rect 539516 -800 539628 480
rect 540698 -800 540810 480
rect 541880 -800 541992 480
rect 543062 -800 543174 480
rect 544244 -800 544356 480
rect 545426 -800 545538 480
rect 546608 -800 546720 480
rect 547790 -800 547902 480
rect 548972 -800 549084 480
rect 550154 -800 550266 480
rect 551336 -800 551448 480
rect 552518 -800 552630 480
rect 553700 -800 553812 480
rect 554882 -800 554994 480
rect 556064 -800 556176 480
rect 557246 -800 557358 480
rect 558428 -800 558540 480
rect 559610 -800 559722 480
rect 560792 -800 560904 480
rect 561974 -800 562086 480
rect 563156 -800 563268 480
rect 564338 -800 564450 480
rect 565520 -800 565632 480
rect 566702 -800 566814 480
rect 567884 -800 567996 480
rect 569066 -800 569178 480
rect 570248 -800 570360 480
rect 571430 -800 571542 480
rect 572612 -800 572724 480
rect 573794 -800 573906 480
rect 574976 -800 575088 480
rect 576158 -800 576270 480
rect 577340 -800 577452 480
rect 578522 -800 578634 480
rect 579704 -800 579816 480
rect 580886 -800 580998 480
rect 582068 -800 582180 480
rect 583250 -800 583362 480
<< metal3 >>
rect 16194 702300 21194 704800
rect 68194 702300 73194 704800
rect 120194 702300 125194 704800
rect 165594 702300 170594 704800
rect 170894 702300 173094 704800
rect 173394 702300 175594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 222594 702300 224794 704800
rect 225094 702300 227294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 324294 702300 326494 704800
rect 326794 702300 328994 704800
rect 329294 702300 334294 704800
rect 413394 702300 418394 704800
rect 465394 702300 470394 704800
rect 510594 702340 515394 704800
rect 520594 702340 525394 704800
rect 566594 702300 571594 704800
rect -800 680242 1700 685242
rect 582300 677984 584800 682984
rect -800 643842 1660 648642
rect 582340 639784 584800 644584
rect -800 633842 1660 638642
rect 582340 629784 584800 634584
rect 583520 589472 584800 589584
rect 583520 588290 584800 588402
rect 583520 587108 584800 587220
rect 583520 585926 584800 586038
rect 583520 584744 584800 584856
rect 583520 583562 584800 583674
rect -800 559442 1660 564242
rect -800 549442 1660 554242
rect 582340 550562 584800 555362
rect 582340 540562 584800 545362
rect -800 511530 480 511642
rect -800 510348 480 510460
rect -800 509166 480 509278
rect -800 507984 480 508096
rect -800 506802 480 506914
rect -800 505620 480 505732
rect 583520 500050 584800 500162
rect 583520 498868 584800 498980
rect 583520 497686 584800 497798
rect 583520 496504 584800 496616
rect 583520 495322 584800 495434
rect 583520 494140 584800 494252
rect -800 468308 480 468420
rect -800 467126 480 467238
rect -800 465944 480 466056
rect -800 464762 480 464874
rect -800 463580 480 463692
rect -800 462398 480 462510
rect 583520 455628 584800 455740
rect 583520 454446 584800 454558
rect 583520 453264 584800 453376
rect 583520 452082 584800 452194
rect 583520 450900 584800 451012
rect 583520 449718 584800 449830
rect -800 425086 480 425198
rect -800 423904 480 424016
rect -800 422722 480 422834
rect -800 421540 480 421652
rect -800 420358 480 420470
rect -800 419176 480 419288
rect 583520 411206 584800 411318
rect 583520 410024 584800 410136
rect 583520 408842 584800 408954
rect 583520 407660 584800 407772
rect 583520 406478 584800 406590
rect 583520 405296 584800 405408
rect -800 381864 480 381976
rect -800 380682 480 380794
rect -800 379500 480 379612
rect -800 378318 480 378430
rect -800 377136 480 377248
rect -800 375954 480 376066
rect 583520 364784 584800 364896
rect 583520 363602 584800 363714
rect 583520 362420 584800 362532
rect 583520 361238 584800 361350
rect 583520 360056 584800 360168
rect 583520 358874 584800 358986
rect -800 338642 480 338754
rect -800 337460 480 337572
rect -800 336278 480 336390
rect -800 335096 480 335208
rect -800 333914 480 334026
rect -800 332732 480 332844
rect 583520 319562 584800 319674
rect 583520 318380 584800 318492
rect 583520 317198 584800 317310
rect 583520 316016 584800 316128
rect 583520 314834 584800 314946
rect 583520 313652 584800 313764
rect -800 295420 480 295532
rect -800 294238 480 294350
rect -800 293056 480 293168
rect -800 291874 480 291986
rect -800 290692 480 290804
rect -800 289510 480 289622
rect 583520 275140 584800 275252
rect 583520 273958 584800 274070
rect 583520 272776 584800 272888
rect 583520 271594 584800 271706
rect 583520 270412 584800 270524
rect 583520 269230 584800 269342
rect -800 252398 480 252510
rect -800 251216 480 251328
rect -800 250034 480 250146
rect -800 248852 480 248964
rect -800 247670 480 247782
rect -800 246488 480 246600
rect 582340 235230 584800 240030
rect 582340 225230 584800 230030
rect -800 214888 1660 219688
rect -800 204888 1660 209688
rect 582340 191430 584800 196230
rect 582340 181430 584800 186230
rect -800 172888 1660 177688
rect -800 162888 1660 167688
rect 582340 146830 584800 151630
rect 582340 136830 584800 141630
rect -800 124776 480 124888
rect -800 123594 480 123706
rect -800 122412 480 122524
rect -800 121230 480 121342
rect -800 120048 480 120160
rect -800 118866 480 118978
rect 583520 95118 584800 95230
rect 583520 93936 584800 94048
rect 583520 92754 584800 92866
rect 583520 91572 584800 91684
rect -800 81554 480 81666
rect -800 80372 480 80484
rect -800 79190 480 79302
rect -800 78008 480 78120
rect -800 76826 480 76938
rect -800 75644 480 75756
rect 583520 50460 584800 50572
rect 583520 49278 584800 49390
rect 583520 48096 584800 48208
rect 583520 46914 584800 47026
rect -800 38332 480 38444
rect -800 37150 480 37262
rect -800 35968 480 36080
rect -800 34786 480 34898
rect -800 33604 480 33716
rect -800 32422 480 32534
rect 583520 24002 584800 24114
rect 583520 22820 584800 22932
rect 583520 21638 584800 21750
rect 583520 20456 584800 20568
rect 583520 19274 584800 19386
rect 583520 18092 584800 18204
rect -800 16910 480 17022
rect 583520 16910 584800 17022
rect -800 15728 480 15840
rect 583520 15728 584800 15840
rect -800 14546 480 14658
rect 583520 14546 584800 14658
rect -800 13364 480 13476
rect 583520 13364 584800 13476
rect -800 12182 480 12294
rect 583520 12182 584800 12294
rect -800 11000 480 11112
rect 583520 11000 584800 11112
rect -800 9818 480 9930
rect 583520 9818 584800 9930
rect -800 8636 480 8748
rect 583520 8636 584800 8748
rect -800 7454 480 7566
rect 583520 7454 584800 7566
rect -800 6272 480 6384
rect 583520 6272 584800 6384
rect -800 5090 480 5202
rect 583520 5090 584800 5202
rect -800 3908 480 4020
rect 583520 3908 584800 4020
rect -800 2726 480 2838
rect 583520 2726 584800 2838
rect -800 1544 480 1656
rect 583520 1544 584800 1656
<< metal4 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
<< metal5 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
<< comment >>
rect -100 704000 584100 704100
rect -100 0 0 704000
rect 584000 0 584100 704000
rect -100 -100 584100 0
use sky130_fd_pr__res_generic_m3_DPAT6Q  R1
timestamp 1695698273
transform 1 0 1100 0 1 687
box -1100 -87 1100 87
use sky130_fd_pr__res_generic_m3_DPAT6Q  R2
timestamp 1695698273
transform 1 0 3300 0 1 687
box -1100 -87 1100 87
use sky130_fd_pr__res_generic_m3_DPAT6Q  R4
timestamp 1695698273
transform 1 0 5500 0 1 687
box -1100 -87 1100 87
use sky130_fd_pr__res_generic_m3_DPAT6Q  R5
timestamp 1695698273
transform 1 0 7700 0 1 687
box -1100 -87 1100 87
use sky130_fd_pr__res_generic_m3_DPAT6Q  R6
timestamp 1695698273
transform 1 0 9900 0 1 687
box -1100 -87 1100 87
use sky130_fd_pr__res_generic_m3_DPAT6Q  R7
timestamp 1695698273
transform 1 0 12100 0 1 687
box -1100 -87 1100 87
use sky130_fd_pr__res_generic_m3_2QNVX3  R8
timestamp 1695698273
transform 1 0 13256 0 1 706
box -56 -106 56 106
use sky130_fd_pr__res_generic_m3_SS5VKG  R9
timestamp 1695698273
transform 1 0 13368 0 1 688
box -56 -88 56 88
use sky130_fd_pr__res_generic_m3_HK2ST4  R11
timestamp 1695698273
transform 1 0 13480 0 1 715
box -56 -115 56 115
use sky130_fd_pr__res_generic_m3_BHQV68  R12
timestamp 1695698273
transform 1 0 13592 0 1 717
box -56 -117 56 117
use ColROs  x3
timestamp 1695698273
transform 1 0 84278 0 1 590538
box -27400 -18560 183690 52740
<< labels >>
flabel metal3 s 583520 269230 584800 269342 0 FreeSans 1120 0 0 0 gpio_analog[0]
port 0 nsew signal bidirectional
flabel metal3 s -800 381864 480 381976 0 FreeSans 1120 0 0 0 gpio_analog[10]
port 1 nsew signal bidirectional
flabel metal3 s -800 338642 480 338754 0 FreeSans 1120 0 0 0 gpio_analog[11]
port 2 nsew signal bidirectional
flabel metal3 s -800 295420 480 295532 0 FreeSans 1120 0 0 0 gpio_analog[12]
port 3 nsew signal bidirectional
flabel metal3 s -800 252398 480 252510 0 FreeSans 1120 0 0 0 gpio_analog[13]
port 4 nsew signal bidirectional
flabel metal3 s -800 124776 480 124888 0 FreeSans 1120 0 0 0 gpio_analog[14]
port 5 nsew signal bidirectional
flabel metal3 s -800 81554 480 81666 0 FreeSans 1120 0 0 0 gpio_analog[15]
port 6 nsew signal bidirectional
flabel metal3 s -800 38332 480 38444 0 FreeSans 1120 0 0 0 gpio_analog[16]
port 7 nsew signal bidirectional
flabel metal3 s -800 16910 480 17022 0 FreeSans 1120 0 0 0 gpio_analog[17]
port 8 nsew signal bidirectional
flabel metal3 s 583520 313652 584800 313764 0 FreeSans 1120 0 0 0 gpio_analog[1]
port 9 nsew signal bidirectional
flabel metal3 s 583520 358874 584800 358986 0 FreeSans 1120 0 0 0 gpio_analog[2]
port 10 nsew signal bidirectional
flabel metal3 s 583520 405296 584800 405408 0 FreeSans 1120 0 0 0 gpio_analog[3]
port 11 nsew signal bidirectional
flabel metal3 s 583520 449718 584800 449830 0 FreeSans 1120 0 0 0 gpio_analog[4]
port 12 nsew signal bidirectional
flabel metal3 s 583520 494140 584800 494252 0 FreeSans 1120 0 0 0 gpio_analog[5]
port 13 nsew signal bidirectional
flabel metal3 s 583520 583562 584800 583674 0 FreeSans 1120 0 0 0 gpio_analog[6]
port 14 nsew signal bidirectional
flabel metal3 s -800 511530 480 511642 0 FreeSans 1120 0 0 0 gpio_analog[7]
port 15 nsew signal bidirectional
flabel metal3 s -800 468308 480 468420 0 FreeSans 1120 0 0 0 gpio_analog[8]
port 16 nsew signal bidirectional
flabel metal3 s -800 425086 480 425198 0 FreeSans 1120 0 0 0 gpio_analog[9]
port 17 nsew signal bidirectional
flabel metal3 s 583520 270412 584800 270524 0 FreeSans 1120 0 0 0 gpio_noesd[0]
port 18 nsew signal bidirectional
flabel metal3 s -800 380682 480 380794 0 FreeSans 1120 0 0 0 gpio_noesd[10]
port 19 nsew signal bidirectional
flabel metal3 s -800 337460 480 337572 0 FreeSans 1120 0 0 0 gpio_noesd[11]
port 20 nsew signal bidirectional
flabel metal3 s -800 294238 480 294350 0 FreeSans 1120 0 0 0 gpio_noesd[12]
port 21 nsew signal bidirectional
flabel metal3 s -800 251216 480 251328 0 FreeSans 1120 0 0 0 gpio_noesd[13]
port 22 nsew signal bidirectional
flabel metal3 s -800 123594 480 123706 0 FreeSans 1120 0 0 0 gpio_noesd[14]
port 23 nsew signal bidirectional
flabel metal3 s -800 80372 480 80484 0 FreeSans 1120 0 0 0 gpio_noesd[15]
port 24 nsew signal bidirectional
flabel metal3 s -800 37150 480 37262 0 FreeSans 1120 0 0 0 gpio_noesd[16]
port 25 nsew signal bidirectional
flabel metal3 s -800 15728 480 15840 0 FreeSans 1120 0 0 0 gpio_noesd[17]
port 26 nsew signal bidirectional
flabel metal3 s 583520 314834 584800 314946 0 FreeSans 1120 0 0 0 gpio_noesd[1]
port 27 nsew signal bidirectional
flabel metal3 s 583520 360056 584800 360168 0 FreeSans 1120 0 0 0 gpio_noesd[2]
port 28 nsew signal bidirectional
flabel metal3 s 583520 406478 584800 406590 0 FreeSans 1120 0 0 0 gpio_noesd[3]
port 29 nsew signal bidirectional
flabel metal3 s 583520 450900 584800 451012 0 FreeSans 1120 0 0 0 gpio_noesd[4]
port 30 nsew signal bidirectional
flabel metal3 s 583520 495322 584800 495434 0 FreeSans 1120 0 0 0 gpio_noesd[5]
port 31 nsew signal bidirectional
flabel metal3 s 583520 584744 584800 584856 0 FreeSans 1120 0 0 0 gpio_noesd[6]
port 32 nsew signal bidirectional
flabel metal3 s -800 510348 480 510460 0 FreeSans 1120 0 0 0 gpio_noesd[7]
port 33 nsew signal bidirectional
flabel metal3 s -800 467126 480 467238 0 FreeSans 1120 0 0 0 gpio_noesd[8]
port 34 nsew signal bidirectional
flabel metal3 s -800 423904 480 424016 0 FreeSans 1120 0 0 0 gpio_noesd[9]
port 35 nsew signal bidirectional
flabel metal3 s 582300 677984 584800 682984 0 FreeSans 1120 0 0 0 io_analog[0]
port 36 nsew signal bidirectional
flabel metal3 s 0 680242 1700 685242 0 FreeSans 1120 0 0 0 io_analog[10]
port 37 nsew signal bidirectional
flabel metal3 s 566594 702300 571594 704800 0 FreeSans 1920 180 0 0 io_analog[1]
port 38 nsew signal bidirectional
flabel metal3 s 465394 702300 470394 704800 0 FreeSans 1920 180 0 0 io_analog[2]
port 39 nsew signal bidirectional
flabel metal3 s 413394 702300 418394 704800 0 FreeSans 1920 180 0 0 io_analog[3]
port 40 nsew signal bidirectional
flabel metal3 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal4 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal5 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal3 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal4 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal5 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal3 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal4 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal5 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal3 s 120194 702300 125194 704800 0 FreeSans 1920 180 0 0 io_analog[7]
port 44 nsew signal bidirectional
flabel metal3 s 68194 702300 73194 704800 0 FreeSans 1920 180 0 0 io_analog[8]
port 45 nsew signal bidirectional
flabel metal3 s 16194 702300 21194 704800 0 FreeSans 1920 180 0 0 io_analog[9]
port 46 nsew signal bidirectional
flabel metal3 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal4 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal5 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal3 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal4 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal5 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal3 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal4 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal5 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal3 s 326794 702300 328994 704800 0 FreeSans 1920 180 0 0 io_clamp_high[0]
port 50 nsew signal bidirectional
flabel metal3 s 225094 702300 227294 704800 0 FreeSans 1920 180 0 0 io_clamp_high[1]
port 51 nsew signal bidirectional
flabel metal3 s 173394 702300 175594 704800 0 FreeSans 1920 180 0 0 io_clamp_high[2]
port 52 nsew signal bidirectional
flabel metal3 s 324294 702300 326494 704800 0 FreeSans 1920 180 0 0 io_clamp_low[0]
port 53 nsew signal bidirectional
flabel metal3 s 222594 702300 224794 704800 0 FreeSans 1920 180 0 0 io_clamp_low[1]
port 54 nsew signal bidirectional
flabel metal3 s 170894 702300 173094 704800 0 FreeSans 1920 180 0 0 io_clamp_low[2]
port 55 nsew signal bidirectional
flabel metal3 s 583520 2726 584800 2838 0 FreeSans 1120 0 0 0 io_in[0]
port 56 nsew signal input
flabel metal3 s 583520 408842 584800 408954 0 FreeSans 1120 0 0 0 io_in[10]
port 57 nsew signal input
flabel metal3 s 583520 453264 584800 453376 0 FreeSans 1120 0 0 0 io_in[11]
port 58 nsew signal input
flabel metal3 s 583520 497686 584800 497798 0 FreeSans 1120 0 0 0 io_in[12]
port 59 nsew signal input
flabel metal3 s 583520 587108 584800 587220 0 FreeSans 1120 0 0 0 io_in[13]
port 60 nsew signal input
flabel metal3 s -800 507984 480 508096 0 FreeSans 1120 0 0 0 io_in[14]
port 61 nsew signal input
flabel metal3 s -800 464762 480 464874 0 FreeSans 1120 0 0 0 io_in[15]
port 62 nsew signal input
flabel metal3 s -800 421540 480 421652 0 FreeSans 1120 0 0 0 io_in[16]
port 63 nsew signal input
flabel metal3 s -800 378318 480 378430 0 FreeSans 1120 0 0 0 io_in[17]
port 64 nsew signal input
flabel metal3 s -800 335096 480 335208 0 FreeSans 1120 0 0 0 io_in[18]
port 65 nsew signal input
flabel metal3 s -800 291874 480 291986 0 FreeSans 1120 0 0 0 io_in[19]
port 66 nsew signal input
flabel metal3 s 583520 7454 584800 7566 0 FreeSans 1120 0 0 0 io_in[1]
port 67 nsew signal input
flabel metal3 s -800 248852 480 248964 0 FreeSans 1120 0 0 0 io_in[20]
port 68 nsew signal input
flabel metal3 s -800 121230 480 121342 0 FreeSans 1120 0 0 0 io_in[21]
port 69 nsew signal input
flabel metal3 s -800 78008 480 78120 0 FreeSans 1120 0 0 0 io_in[22]
port 70 nsew signal input
flabel metal3 s -800 34786 480 34898 0 FreeSans 1120 0 0 0 io_in[23]
port 71 nsew signal input
flabel metal3 s -800 13364 480 13476 0 FreeSans 1120 0 0 0 io_in[24]
port 72 nsew signal input
flabel metal3 s -800 8636 480 8748 0 FreeSans 1120 0 0 0 io_in[25]
port 73 nsew signal input
flabel metal3 s -800 3908 480 4020 0 FreeSans 1120 0 0 0 io_in[26]
port 74 nsew signal input
flabel metal3 s 583520 12182 584800 12294 0 FreeSans 1120 0 0 0 io_in[2]
port 75 nsew signal input
flabel metal3 s 583520 16910 584800 17022 0 FreeSans 1120 0 0 0 io_in[3]
port 76 nsew signal input
flabel metal3 s 583520 21638 584800 21750 0 FreeSans 1120 0 0 0 io_in[4]
port 77 nsew signal input
flabel metal3 s 583520 48096 584800 48208 0 FreeSans 1120 0 0 0 io_in[5]
port 78 nsew signal input
flabel metal3 s 583520 92754 584800 92866 0 FreeSans 1120 0 0 0 io_in[6]
port 79 nsew signal input
flabel metal3 s 583520 272776 584800 272888 0 FreeSans 1120 0 0 0 io_in[7]
port 80 nsew signal input
flabel metal3 s 583520 317198 584800 317310 0 FreeSans 1120 0 0 0 io_in[8]
port 81 nsew signal input
flabel metal3 s 583520 362420 584800 362532 0 FreeSans 1120 0 0 0 io_in[9]
port 82 nsew signal input
flabel metal3 s 583520 1544 584800 1656 0 FreeSans 1120 0 0 0 io_in_3v3[0]
port 83 nsew signal input
flabel metal3 s 583520 407660 584800 407772 0 FreeSans 1120 0 0 0 io_in_3v3[10]
port 84 nsew signal input
flabel metal3 s 583520 452082 584800 452194 0 FreeSans 1120 0 0 0 io_in_3v3[11]
port 85 nsew signal input
flabel metal3 s 583520 496504 584800 496616 0 FreeSans 1120 0 0 0 io_in_3v3[12]
port 86 nsew signal input
flabel metal3 s 583520 585926 584800 586038 0 FreeSans 1120 0 0 0 io_in_3v3[13]
port 87 nsew signal input
flabel metal3 s -800 509166 480 509278 0 FreeSans 1120 0 0 0 io_in_3v3[14]
port 88 nsew signal input
flabel metal3 s -800 465944 480 466056 0 FreeSans 1120 0 0 0 io_in_3v3[15]
port 89 nsew signal input
flabel metal3 s -800 422722 480 422834 0 FreeSans 1120 0 0 0 io_in_3v3[16]
port 90 nsew signal input
flabel metal3 s -800 379500 480 379612 0 FreeSans 1120 0 0 0 io_in_3v3[17]
port 91 nsew signal input
flabel metal3 s -800 336278 480 336390 0 FreeSans 1120 0 0 0 io_in_3v3[18]
port 92 nsew signal input
flabel metal3 s -800 293056 480 293168 0 FreeSans 1120 0 0 0 io_in_3v3[19]
port 93 nsew signal input
flabel metal3 s 583520 6272 584800 6384 0 FreeSans 1120 0 0 0 io_in_3v3[1]
port 94 nsew signal input
flabel metal3 s -800 250034 480 250146 0 FreeSans 1120 0 0 0 io_in_3v3[20]
port 95 nsew signal input
flabel metal3 s -800 122412 480 122524 0 FreeSans 1120 0 0 0 io_in_3v3[21]
port 96 nsew signal input
flabel metal3 s -800 79190 480 79302 0 FreeSans 1120 0 0 0 io_in_3v3[22]
port 97 nsew signal input
flabel metal3 s -800 35968 480 36080 0 FreeSans 1120 0 0 0 io_in_3v3[23]
port 98 nsew signal input
flabel metal3 s -800 14546 480 14658 0 FreeSans 1120 0 0 0 io_in_3v3[24]
port 99 nsew signal input
flabel metal3 s -800 9818 480 9930 0 FreeSans 1120 0 0 0 io_in_3v3[25]
port 100 nsew signal input
flabel metal3 s -800 5090 480 5202 0 FreeSans 1120 0 0 0 io_in_3v3[26]
port 101 nsew signal input
flabel metal3 s 583520 11000 584800 11112 0 FreeSans 1120 0 0 0 io_in_3v3[2]
port 102 nsew signal input
flabel metal3 s 583520 15728 584800 15840 0 FreeSans 1120 0 0 0 io_in_3v3[3]
port 103 nsew signal input
flabel metal3 s 583520 20456 584800 20568 0 FreeSans 1120 0 0 0 io_in_3v3[4]
port 104 nsew signal input
flabel metal3 s 583520 46914 584800 47026 0 FreeSans 1120 0 0 0 io_in_3v3[5]
port 105 nsew signal input
flabel metal3 s 583520 91572 584800 91684 0 FreeSans 1120 0 0 0 io_in_3v3[6]
port 106 nsew signal input
flabel metal3 s 583520 271594 584800 271706 0 FreeSans 1120 0 0 0 io_in_3v3[7]
port 107 nsew signal input
flabel metal3 s 583520 316016 584800 316128 0 FreeSans 1120 0 0 0 io_in_3v3[8]
port 108 nsew signal input
flabel metal3 s 583520 361238 584800 361350 0 FreeSans 1120 0 0 0 io_in_3v3[9]
port 109 nsew signal input
flabel metal3 s 583520 5090 584800 5202 0 FreeSans 1120 0 0 0 io_oeb[0]
port 110 nsew signal tristate
flabel metal3 s 583520 411206 584800 411318 0 FreeSans 1120 0 0 0 io_oeb[10]
port 111 nsew signal tristate
flabel metal3 s 583520 455628 584800 455740 0 FreeSans 1120 0 0 0 io_oeb[11]
port 112 nsew signal tristate
flabel metal3 s 583520 500050 584800 500162 0 FreeSans 1120 0 0 0 io_oeb[12]
port 113 nsew signal tristate
flabel metal3 s 583520 589472 584800 589584 0 FreeSans 1120 0 0 0 io_oeb[13]
port 114 nsew signal tristate
flabel metal3 s -800 505620 480 505732 0 FreeSans 1120 0 0 0 io_oeb[14]
port 115 nsew signal tristate
flabel metal3 s -800 462398 480 462510 0 FreeSans 1120 0 0 0 io_oeb[15]
port 116 nsew signal tristate
flabel metal3 s -800 419176 480 419288 0 FreeSans 1120 0 0 0 io_oeb[16]
port 117 nsew signal tristate
flabel metal3 s -800 375954 480 376066 0 FreeSans 1120 0 0 0 io_oeb[17]
port 118 nsew signal tristate
flabel metal3 s -800 332732 480 332844 0 FreeSans 1120 0 0 0 io_oeb[18]
port 119 nsew signal tristate
flabel metal3 s -800 289510 480 289622 0 FreeSans 1120 0 0 0 io_oeb[19]
port 120 nsew signal tristate
flabel metal3 s 583520 9818 584800 9930 0 FreeSans 1120 0 0 0 io_oeb[1]
port 121 nsew signal tristate
flabel metal3 s -800 246488 480 246600 0 FreeSans 1120 0 0 0 io_oeb[20]
port 122 nsew signal tristate
flabel metal3 s -800 118866 480 118978 0 FreeSans 1120 0 0 0 io_oeb[21]
port 123 nsew signal tristate
flabel metal3 s -800 75644 480 75756 0 FreeSans 1120 0 0 0 io_oeb[22]
port 124 nsew signal tristate
flabel metal3 s -800 32422 480 32534 0 FreeSans 1120 0 0 0 io_oeb[23]
port 125 nsew signal tristate
flabel metal3 s -800 11000 480 11112 0 FreeSans 1120 0 0 0 io_oeb[24]
port 126 nsew signal tristate
flabel metal3 s -800 6272 480 6384 0 FreeSans 1120 0 0 0 io_oeb[25]
port 127 nsew signal tristate
flabel metal3 s -800 1544 480 1656 0 FreeSans 1120 0 0 0 io_oeb[26]
port 128 nsew signal tristate
flabel metal3 s 583520 14546 584800 14658 0 FreeSans 1120 0 0 0 io_oeb[2]
port 129 nsew signal tristate
flabel metal3 s 583520 19274 584800 19386 0 FreeSans 1120 0 0 0 io_oeb[3]
port 130 nsew signal tristate
flabel metal3 s 583520 24002 584800 24114 0 FreeSans 1120 0 0 0 io_oeb[4]
port 131 nsew signal tristate
flabel metal3 s 583520 50460 584800 50572 0 FreeSans 1120 0 0 0 io_oeb[5]
port 132 nsew signal tristate
flabel metal3 s 583520 95118 584800 95230 0 FreeSans 1120 0 0 0 io_oeb[6]
port 133 nsew signal tristate
flabel metal3 s 583520 275140 584800 275252 0 FreeSans 1120 0 0 0 io_oeb[7]
port 134 nsew signal tristate
flabel metal3 s 583520 319562 584800 319674 0 FreeSans 1120 0 0 0 io_oeb[8]
port 135 nsew signal tristate
flabel metal3 s 583520 364784 584800 364896 0 FreeSans 1120 0 0 0 io_oeb[9]
port 136 nsew signal tristate
flabel metal3 s 583520 3908 584800 4020 0 FreeSans 1120 0 0 0 io_out[0]
port 137 nsew signal tristate
flabel metal3 s 583520 410024 584800 410136 0 FreeSans 1120 0 0 0 io_out[10]
port 138 nsew signal tristate
flabel metal3 s 583520 454446 584800 454558 0 FreeSans 1120 0 0 0 io_out[11]
port 139 nsew signal tristate
flabel metal3 s 583520 498868 584800 498980 0 FreeSans 1120 0 0 0 io_out[12]
port 140 nsew signal tristate
flabel metal3 s 583520 588290 584800 588402 0 FreeSans 1120 0 0 0 io_out[13]
port 141 nsew signal tristate
flabel metal3 s -800 506802 480 506914 0 FreeSans 1120 0 0 0 io_out[14]
port 142 nsew signal tristate
flabel metal3 s -800 463580 480 463692 0 FreeSans 1120 0 0 0 io_out[15]
port 143 nsew signal tristate
flabel metal3 s -800 420358 480 420470 0 FreeSans 1120 0 0 0 io_out[16]
port 144 nsew signal tristate
flabel metal3 s -800 377136 480 377248 0 FreeSans 1120 0 0 0 io_out[17]
port 145 nsew signal tristate
flabel metal3 s -800 333914 480 334026 0 FreeSans 1120 0 0 0 io_out[18]
port 146 nsew signal tristate
flabel metal3 s -800 290692 480 290804 0 FreeSans 1120 0 0 0 io_out[19]
port 147 nsew signal tristate
flabel metal3 s 583520 8636 584800 8748 0 FreeSans 1120 0 0 0 io_out[1]
port 148 nsew signal tristate
flabel metal3 s -800 247670 480 247782 0 FreeSans 1120 0 0 0 io_out[20]
port 149 nsew signal tristate
flabel metal3 s -800 120048 480 120160 0 FreeSans 1120 0 0 0 io_out[21]
port 150 nsew signal tristate
flabel metal3 s -800 76826 480 76938 0 FreeSans 1120 0 0 0 io_out[22]
port 151 nsew signal tristate
flabel metal3 s -800 33604 480 33716 0 FreeSans 1120 0 0 0 io_out[23]
port 152 nsew signal tristate
flabel metal3 s -800 12182 480 12294 0 FreeSans 1120 0 0 0 io_out[24]
port 153 nsew signal tristate
flabel metal3 s -800 7454 480 7566 0 FreeSans 1120 0 0 0 io_out[25]
port 154 nsew signal tristate
flabel metal3 s -800 2726 480 2838 0 FreeSans 1120 0 0 0 io_out[26]
port 155 nsew signal tristate
flabel metal3 s 583520 13364 584800 13476 0 FreeSans 1120 0 0 0 io_out[2]
port 156 nsew signal tristate
flabel metal3 s 583520 18092 584800 18204 0 FreeSans 1120 0 0 0 io_out[3]
port 157 nsew signal tristate
flabel metal3 s 583520 22820 584800 22932 0 FreeSans 1120 0 0 0 io_out[4]
port 158 nsew signal tristate
flabel metal3 s 583520 49278 584800 49390 0 FreeSans 1120 0 0 0 io_out[5]
port 159 nsew signal tristate
flabel metal3 s 583520 93936 584800 94048 0 FreeSans 1120 0 0 0 io_out[6]
port 160 nsew signal tristate
flabel metal3 s 583520 273958 584800 274070 0 FreeSans 1120 0 0 0 io_out[7]
port 161 nsew signal tristate
flabel metal3 s 583520 318380 584800 318492 0 FreeSans 1120 0 0 0 io_out[8]
port 162 nsew signal tristate
flabel metal3 s 583520 363602 584800 363714 0 FreeSans 1120 0 0 0 io_out[9]
port 163 nsew signal tristate
flabel metal2 s 125816 -800 125928 480 0 FreeSans 1120 90 0 0 la_data_in[0]
port 164 nsew signal input
flabel metal2 s 480416 -800 480528 480 0 FreeSans 1120 90 0 0 la_data_in[100]
port 165 nsew signal input
flabel metal2 s 483962 -800 484074 480 0 FreeSans 1120 90 0 0 la_data_in[101]
port 166 nsew signal input
flabel metal2 s 487508 -800 487620 480 0 FreeSans 1120 90 0 0 la_data_in[102]
port 167 nsew signal input
flabel metal2 s 491054 -800 491166 480 0 FreeSans 1120 90 0 0 la_data_in[103]
port 168 nsew signal input
flabel metal2 s 494600 -800 494712 480 0 FreeSans 1120 90 0 0 la_data_in[104]
port 169 nsew signal input
flabel metal2 s 498146 -800 498258 480 0 FreeSans 1120 90 0 0 la_data_in[105]
port 170 nsew signal input
flabel metal2 s 501692 -800 501804 480 0 FreeSans 1120 90 0 0 la_data_in[106]
port 171 nsew signal input
flabel metal2 s 505238 -800 505350 480 0 FreeSans 1120 90 0 0 la_data_in[107]
port 172 nsew signal input
flabel metal2 s 508784 -800 508896 480 0 FreeSans 1120 90 0 0 la_data_in[108]
port 173 nsew signal input
flabel metal2 s 512330 -800 512442 480 0 FreeSans 1120 90 0 0 la_data_in[109]
port 174 nsew signal input
flabel metal2 s 161276 -800 161388 480 0 FreeSans 1120 90 0 0 la_data_in[10]
port 175 nsew signal input
flabel metal2 s 515876 -800 515988 480 0 FreeSans 1120 90 0 0 la_data_in[110]
port 176 nsew signal input
flabel metal2 s 519422 -800 519534 480 0 FreeSans 1120 90 0 0 la_data_in[111]
port 177 nsew signal input
flabel metal2 s 522968 -800 523080 480 0 FreeSans 1120 90 0 0 la_data_in[112]
port 178 nsew signal input
flabel metal2 s 526514 -800 526626 480 0 FreeSans 1120 90 0 0 la_data_in[113]
port 179 nsew signal input
flabel metal2 s 530060 -800 530172 480 0 FreeSans 1120 90 0 0 la_data_in[114]
port 180 nsew signal input
flabel metal2 s 533606 -800 533718 480 0 FreeSans 1120 90 0 0 la_data_in[115]
port 181 nsew signal input
flabel metal2 s 537152 -800 537264 480 0 FreeSans 1120 90 0 0 la_data_in[116]
port 182 nsew signal input
flabel metal2 s 540698 -800 540810 480 0 FreeSans 1120 90 0 0 la_data_in[117]
port 183 nsew signal input
flabel metal2 s 544244 -800 544356 480 0 FreeSans 1120 90 0 0 la_data_in[118]
port 184 nsew signal input
flabel metal2 s 547790 -800 547902 480 0 FreeSans 1120 90 0 0 la_data_in[119]
port 185 nsew signal input
flabel metal2 s 164822 -800 164934 480 0 FreeSans 1120 90 0 0 la_data_in[11]
port 186 nsew signal input
flabel metal2 s 551336 -800 551448 480 0 FreeSans 1120 90 0 0 la_data_in[120]
port 187 nsew signal input
flabel metal2 s 554882 -800 554994 480 0 FreeSans 1120 90 0 0 la_data_in[121]
port 188 nsew signal input
flabel metal2 s 558428 -800 558540 480 0 FreeSans 1120 90 0 0 la_data_in[122]
port 189 nsew signal input
flabel metal2 s 561974 -800 562086 480 0 FreeSans 1120 90 0 0 la_data_in[123]
port 190 nsew signal input
flabel metal2 s 565520 -800 565632 480 0 FreeSans 1120 90 0 0 la_data_in[124]
port 191 nsew signal input
flabel metal2 s 569066 -800 569178 480 0 FreeSans 1120 90 0 0 la_data_in[125]
port 192 nsew signal input
flabel metal2 s 572612 -800 572724 480 0 FreeSans 1120 90 0 0 la_data_in[126]
port 193 nsew signal input
flabel metal2 s 576158 -800 576270 480 0 FreeSans 1120 90 0 0 la_data_in[127]
port 194 nsew signal input
flabel metal2 s 168368 -800 168480 480 0 FreeSans 1120 90 0 0 la_data_in[12]
port 195 nsew signal input
flabel metal2 s 171914 -800 172026 480 0 FreeSans 1120 90 0 0 la_data_in[13]
port 196 nsew signal input
flabel metal2 s 175460 -800 175572 480 0 FreeSans 1120 90 0 0 la_data_in[14]
port 197 nsew signal input
flabel metal2 s 179006 -800 179118 480 0 FreeSans 1120 90 0 0 la_data_in[15]
port 198 nsew signal input
flabel metal2 s 182552 -800 182664 480 0 FreeSans 1120 90 0 0 la_data_in[16]
port 199 nsew signal input
flabel metal2 s 186098 -800 186210 480 0 FreeSans 1120 90 0 0 la_data_in[17]
port 200 nsew signal input
flabel metal2 s 189644 -800 189756 480 0 FreeSans 1120 90 0 0 la_data_in[18]
port 201 nsew signal input
flabel metal2 s 193190 -800 193302 480 0 FreeSans 1120 90 0 0 la_data_in[19]
port 202 nsew signal input
flabel metal2 s 129362 -800 129474 480 0 FreeSans 1120 90 0 0 la_data_in[1]
port 203 nsew signal input
flabel metal2 s 196736 -800 196848 480 0 FreeSans 1120 90 0 0 la_data_in[20]
port 204 nsew signal input
flabel metal2 s 200282 -800 200394 480 0 FreeSans 1120 90 0 0 la_data_in[21]
port 205 nsew signal input
flabel metal2 s 203828 -800 203940 480 0 FreeSans 1120 90 0 0 la_data_in[22]
port 206 nsew signal input
flabel metal2 s 207374 -800 207486 480 0 FreeSans 1120 90 0 0 la_data_in[23]
port 207 nsew signal input
flabel metal2 s 210920 -800 211032 480 0 FreeSans 1120 90 0 0 la_data_in[24]
port 208 nsew signal input
flabel metal2 s 214466 -800 214578 480 0 FreeSans 1120 90 0 0 la_data_in[25]
port 209 nsew signal input
flabel metal2 s 218012 -800 218124 480 0 FreeSans 1120 90 0 0 la_data_in[26]
port 210 nsew signal input
flabel metal2 s 221558 -800 221670 480 0 FreeSans 1120 90 0 0 la_data_in[27]
port 211 nsew signal input
flabel metal2 s 225104 -800 225216 480 0 FreeSans 1120 90 0 0 la_data_in[28]
port 212 nsew signal input
flabel metal2 s 228650 -800 228762 480 0 FreeSans 1120 90 0 0 la_data_in[29]
port 213 nsew signal input
flabel metal2 s 132908 -800 133020 480 0 FreeSans 1120 90 0 0 la_data_in[2]
port 214 nsew signal input
flabel metal2 s 232196 -800 232308 480 0 FreeSans 1120 90 0 0 la_data_in[30]
port 215 nsew signal input
flabel metal2 s 235742 -800 235854 480 0 FreeSans 1120 90 0 0 la_data_in[31]
port 216 nsew signal input
flabel metal2 s 239288 -800 239400 480 0 FreeSans 1120 90 0 0 la_data_in[32]
port 217 nsew signal input
flabel metal2 s 242834 -800 242946 480 0 FreeSans 1120 90 0 0 la_data_in[33]
port 218 nsew signal input
flabel metal2 s 246380 -800 246492 480 0 FreeSans 1120 90 0 0 la_data_in[34]
port 219 nsew signal input
flabel metal2 s 249926 -800 250038 480 0 FreeSans 1120 90 0 0 la_data_in[35]
port 220 nsew signal input
flabel metal2 s 253472 -800 253584 480 0 FreeSans 1120 90 0 0 la_data_in[36]
port 221 nsew signal input
flabel metal2 s 257018 -800 257130 480 0 FreeSans 1120 90 0 0 la_data_in[37]
port 222 nsew signal input
flabel metal2 s 260564 -800 260676 480 0 FreeSans 1120 90 0 0 la_data_in[38]
port 223 nsew signal input
flabel metal2 s 264110 -800 264222 480 0 FreeSans 1120 90 0 0 la_data_in[39]
port 224 nsew signal input
flabel metal2 s 136454 -800 136566 480 0 FreeSans 1120 90 0 0 la_data_in[3]
port 225 nsew signal input
flabel metal2 s 267656 -800 267768 480 0 FreeSans 1120 90 0 0 la_data_in[40]
port 226 nsew signal input
flabel metal2 s 271202 -800 271314 480 0 FreeSans 1120 90 0 0 la_data_in[41]
port 227 nsew signal input
flabel metal2 s 274748 -800 274860 480 0 FreeSans 1120 90 0 0 la_data_in[42]
port 228 nsew signal input
flabel metal2 s 278294 -800 278406 480 0 FreeSans 1120 90 0 0 la_data_in[43]
port 229 nsew signal input
flabel metal2 s 281840 -800 281952 480 0 FreeSans 1120 90 0 0 la_data_in[44]
port 230 nsew signal input
flabel metal2 s 285386 -800 285498 480 0 FreeSans 1120 90 0 0 la_data_in[45]
port 231 nsew signal input
flabel metal2 s 288932 -800 289044 480 0 FreeSans 1120 90 0 0 la_data_in[46]
port 232 nsew signal input
flabel metal2 s 292478 -800 292590 480 0 FreeSans 1120 90 0 0 la_data_in[47]
port 233 nsew signal input
flabel metal2 s 296024 -800 296136 480 0 FreeSans 1120 90 0 0 la_data_in[48]
port 234 nsew signal input
flabel metal2 s 299570 -800 299682 480 0 FreeSans 1120 90 0 0 la_data_in[49]
port 235 nsew signal input
flabel metal2 s 140000 -800 140112 480 0 FreeSans 1120 90 0 0 la_data_in[4]
port 236 nsew signal input
flabel metal2 s 303116 -800 303228 480 0 FreeSans 1120 90 0 0 la_data_in[50]
port 237 nsew signal input
flabel metal2 s 306662 -800 306774 480 0 FreeSans 1120 90 0 0 la_data_in[51]
port 238 nsew signal input
flabel metal2 s 310208 -800 310320 480 0 FreeSans 1120 90 0 0 la_data_in[52]
port 239 nsew signal input
flabel metal2 s 313754 -800 313866 480 0 FreeSans 1120 90 0 0 la_data_in[53]
port 240 nsew signal input
flabel metal2 s 317300 -800 317412 480 0 FreeSans 1120 90 0 0 la_data_in[54]
port 241 nsew signal input
flabel metal2 s 320846 -800 320958 480 0 FreeSans 1120 90 0 0 la_data_in[55]
port 242 nsew signal input
flabel metal2 s 324392 -800 324504 480 0 FreeSans 1120 90 0 0 la_data_in[56]
port 243 nsew signal input
flabel metal2 s 327938 -800 328050 480 0 FreeSans 1120 90 0 0 la_data_in[57]
port 244 nsew signal input
flabel metal2 s 331484 -800 331596 480 0 FreeSans 1120 90 0 0 la_data_in[58]
port 245 nsew signal input
flabel metal2 s 335030 -800 335142 480 0 FreeSans 1120 90 0 0 la_data_in[59]
port 246 nsew signal input
flabel metal2 s 143546 -800 143658 480 0 FreeSans 1120 90 0 0 la_data_in[5]
port 247 nsew signal input
flabel metal2 s 338576 -800 338688 480 0 FreeSans 1120 90 0 0 la_data_in[60]
port 248 nsew signal input
flabel metal2 s 342122 -800 342234 480 0 FreeSans 1120 90 0 0 la_data_in[61]
port 249 nsew signal input
flabel metal2 s 345668 -800 345780 480 0 FreeSans 1120 90 0 0 la_data_in[62]
port 250 nsew signal input
flabel metal2 s 349214 -800 349326 480 0 FreeSans 1120 90 0 0 la_data_in[63]
port 251 nsew signal input
flabel metal2 s 352760 -800 352872 480 0 FreeSans 1120 90 0 0 la_data_in[64]
port 252 nsew signal input
flabel metal2 s 356306 -800 356418 480 0 FreeSans 1120 90 0 0 la_data_in[65]
port 253 nsew signal input
flabel metal2 s 359852 -800 359964 480 0 FreeSans 1120 90 0 0 la_data_in[66]
port 254 nsew signal input
flabel metal2 s 363398 -800 363510 480 0 FreeSans 1120 90 0 0 la_data_in[67]
port 255 nsew signal input
flabel metal2 s 366944 -800 367056 480 0 FreeSans 1120 90 0 0 la_data_in[68]
port 256 nsew signal input
flabel metal2 s 370490 -800 370602 480 0 FreeSans 1120 90 0 0 la_data_in[69]
port 257 nsew signal input
flabel metal2 s 147092 -800 147204 480 0 FreeSans 1120 90 0 0 la_data_in[6]
port 258 nsew signal input
flabel metal2 s 374036 -800 374148 480 0 FreeSans 1120 90 0 0 la_data_in[70]
port 259 nsew signal input
flabel metal2 s 377582 -800 377694 480 0 FreeSans 1120 90 0 0 la_data_in[71]
port 260 nsew signal input
flabel metal2 s 381128 -800 381240 480 0 FreeSans 1120 90 0 0 la_data_in[72]
port 261 nsew signal input
flabel metal2 s 384674 -800 384786 480 0 FreeSans 1120 90 0 0 la_data_in[73]
port 262 nsew signal input
flabel metal2 s 388220 -800 388332 480 0 FreeSans 1120 90 0 0 la_data_in[74]
port 263 nsew signal input
flabel metal2 s 391766 -800 391878 480 0 FreeSans 1120 90 0 0 la_data_in[75]
port 264 nsew signal input
flabel metal2 s 395312 -800 395424 480 0 FreeSans 1120 90 0 0 la_data_in[76]
port 265 nsew signal input
flabel metal2 s 398858 -800 398970 480 0 FreeSans 1120 90 0 0 la_data_in[77]
port 266 nsew signal input
flabel metal2 s 402404 -800 402516 480 0 FreeSans 1120 90 0 0 la_data_in[78]
port 267 nsew signal input
flabel metal2 s 405950 -800 406062 480 0 FreeSans 1120 90 0 0 la_data_in[79]
port 268 nsew signal input
flabel metal2 s 150638 -800 150750 480 0 FreeSans 1120 90 0 0 la_data_in[7]
port 269 nsew signal input
flabel metal2 s 409496 -800 409608 480 0 FreeSans 1120 90 0 0 la_data_in[80]
port 270 nsew signal input
flabel metal2 s 413042 -800 413154 480 0 FreeSans 1120 90 0 0 la_data_in[81]
port 271 nsew signal input
flabel metal2 s 416588 -800 416700 480 0 FreeSans 1120 90 0 0 la_data_in[82]
port 272 nsew signal input
flabel metal2 s 420134 -800 420246 480 0 FreeSans 1120 90 0 0 la_data_in[83]
port 273 nsew signal input
flabel metal2 s 423680 -800 423792 480 0 FreeSans 1120 90 0 0 la_data_in[84]
port 274 nsew signal input
flabel metal2 s 427226 -800 427338 480 0 FreeSans 1120 90 0 0 la_data_in[85]
port 275 nsew signal input
flabel metal2 s 430772 -800 430884 480 0 FreeSans 1120 90 0 0 la_data_in[86]
port 276 nsew signal input
flabel metal2 s 434318 -800 434430 480 0 FreeSans 1120 90 0 0 la_data_in[87]
port 277 nsew signal input
flabel metal2 s 437864 -800 437976 480 0 FreeSans 1120 90 0 0 la_data_in[88]
port 278 nsew signal input
flabel metal2 s 441410 -800 441522 480 0 FreeSans 1120 90 0 0 la_data_in[89]
port 279 nsew signal input
flabel metal2 s 154184 -800 154296 480 0 FreeSans 1120 90 0 0 la_data_in[8]
port 280 nsew signal input
flabel metal2 s 444956 -800 445068 480 0 FreeSans 1120 90 0 0 la_data_in[90]
port 281 nsew signal input
flabel metal2 s 448502 -800 448614 480 0 FreeSans 1120 90 0 0 la_data_in[91]
port 282 nsew signal input
flabel metal2 s 452048 -800 452160 480 0 FreeSans 1120 90 0 0 la_data_in[92]
port 283 nsew signal input
flabel metal2 s 455594 -800 455706 480 0 FreeSans 1120 90 0 0 la_data_in[93]
port 284 nsew signal input
flabel metal2 s 459140 -800 459252 480 0 FreeSans 1120 90 0 0 la_data_in[94]
port 285 nsew signal input
flabel metal2 s 462686 -800 462798 480 0 FreeSans 1120 90 0 0 la_data_in[95]
port 286 nsew signal input
flabel metal2 s 466232 -800 466344 480 0 FreeSans 1120 90 0 0 la_data_in[96]
port 287 nsew signal input
flabel metal2 s 469778 -800 469890 480 0 FreeSans 1120 90 0 0 la_data_in[97]
port 288 nsew signal input
flabel metal2 s 473324 -800 473436 480 0 FreeSans 1120 90 0 0 la_data_in[98]
port 289 nsew signal input
flabel metal2 s 476870 -800 476982 480 0 FreeSans 1120 90 0 0 la_data_in[99]
port 290 nsew signal input
flabel metal2 s 157730 -800 157842 480 0 FreeSans 1120 90 0 0 la_data_in[9]
port 291 nsew signal input
flabel metal2 s 126998 -800 127110 480 0 FreeSans 1120 90 0 0 la_data_out[0]
port 292 nsew signal tristate
flabel metal2 s 481598 -800 481710 480 0 FreeSans 1120 90 0 0 la_data_out[100]
port 293 nsew signal tristate
flabel metal2 s 485144 -800 485256 480 0 FreeSans 1120 90 0 0 la_data_out[101]
port 294 nsew signal tristate
flabel metal2 s 488690 -800 488802 480 0 FreeSans 1120 90 0 0 la_data_out[102]
port 295 nsew signal tristate
flabel metal2 s 492236 -800 492348 480 0 FreeSans 1120 90 0 0 la_data_out[103]
port 296 nsew signal tristate
flabel metal2 s 495782 -800 495894 480 0 FreeSans 1120 90 0 0 la_data_out[104]
port 297 nsew signal tristate
flabel metal2 s 499328 -800 499440 480 0 FreeSans 1120 90 0 0 la_data_out[105]
port 298 nsew signal tristate
flabel metal2 s 502874 -800 502986 480 0 FreeSans 1120 90 0 0 la_data_out[106]
port 299 nsew signal tristate
flabel metal2 s 506420 -800 506532 480 0 FreeSans 1120 90 0 0 la_data_out[107]
port 300 nsew signal tristate
flabel metal2 s 509966 -800 510078 480 0 FreeSans 1120 90 0 0 la_data_out[108]
port 301 nsew signal tristate
flabel metal2 s 513512 -800 513624 480 0 FreeSans 1120 90 0 0 la_data_out[109]
port 302 nsew signal tristate
flabel metal2 s 162458 -800 162570 480 0 FreeSans 1120 90 0 0 la_data_out[10]
port 303 nsew signal tristate
flabel metal2 s 517058 -800 517170 480 0 FreeSans 1120 90 0 0 la_data_out[110]
port 304 nsew signal tristate
flabel metal2 s 520604 -800 520716 480 0 FreeSans 1120 90 0 0 la_data_out[111]
port 305 nsew signal tristate
flabel metal2 s 524150 -800 524262 480 0 FreeSans 1120 90 0 0 la_data_out[112]
port 306 nsew signal tristate
flabel metal2 s 527696 -800 527808 480 0 FreeSans 1120 90 0 0 la_data_out[113]
port 307 nsew signal tristate
flabel metal2 s 531242 -800 531354 480 0 FreeSans 1120 90 0 0 la_data_out[114]
port 308 nsew signal tristate
flabel metal2 s 534788 -800 534900 480 0 FreeSans 1120 90 0 0 la_data_out[115]
port 309 nsew signal tristate
flabel metal2 s 538334 -800 538446 480 0 FreeSans 1120 90 0 0 la_data_out[116]
port 310 nsew signal tristate
flabel metal2 s 541880 -800 541992 480 0 FreeSans 1120 90 0 0 la_data_out[117]
port 311 nsew signal tristate
flabel metal2 s 545426 -800 545538 480 0 FreeSans 1120 90 0 0 la_data_out[118]
port 312 nsew signal tristate
flabel metal2 s 548972 -800 549084 480 0 FreeSans 1120 90 0 0 la_data_out[119]
port 313 nsew signal tristate
flabel metal2 s 166004 -800 166116 480 0 FreeSans 1120 90 0 0 la_data_out[11]
port 314 nsew signal tristate
flabel metal2 s 552518 -800 552630 480 0 FreeSans 1120 90 0 0 la_data_out[120]
port 315 nsew signal tristate
flabel metal2 s 556064 -800 556176 480 0 FreeSans 1120 90 0 0 la_data_out[121]
port 316 nsew signal tristate
flabel metal2 s 559610 -800 559722 480 0 FreeSans 1120 90 0 0 la_data_out[122]
port 317 nsew signal tristate
flabel metal2 s 563156 -800 563268 480 0 FreeSans 1120 90 0 0 la_data_out[123]
port 318 nsew signal tristate
flabel metal2 s 566702 -800 566814 480 0 FreeSans 1120 90 0 0 la_data_out[124]
port 319 nsew signal tristate
flabel metal2 s 570248 -800 570360 480 0 FreeSans 1120 90 0 0 la_data_out[125]
port 320 nsew signal tristate
flabel metal2 s 573794 -800 573906 480 0 FreeSans 1120 90 0 0 la_data_out[126]
port 321 nsew signal tristate
flabel metal2 s 577340 -800 577452 480 0 FreeSans 1120 90 0 0 la_data_out[127]
port 322 nsew signal tristate
flabel metal2 s 169550 -800 169662 480 0 FreeSans 1120 90 0 0 la_data_out[12]
port 323 nsew signal tristate
flabel metal2 s 173096 -800 173208 480 0 FreeSans 1120 90 0 0 la_data_out[13]
port 324 nsew signal tristate
flabel metal2 s 176642 -800 176754 480 0 FreeSans 1120 90 0 0 la_data_out[14]
port 325 nsew signal tristate
flabel metal2 s 180188 -800 180300 480 0 FreeSans 1120 90 0 0 la_data_out[15]
port 326 nsew signal tristate
flabel metal2 s 183734 -800 183846 480 0 FreeSans 1120 90 0 0 la_data_out[16]
port 327 nsew signal tristate
flabel metal2 s 187280 -800 187392 480 0 FreeSans 1120 90 0 0 la_data_out[17]
port 328 nsew signal tristate
flabel metal2 s 190826 -800 190938 480 0 FreeSans 1120 90 0 0 la_data_out[18]
port 329 nsew signal tristate
flabel metal2 s 194372 -800 194484 480 0 FreeSans 1120 90 0 0 la_data_out[19]
port 330 nsew signal tristate
flabel metal2 s 130544 -800 130656 480 0 FreeSans 1120 90 0 0 la_data_out[1]
port 331 nsew signal tristate
flabel metal2 s 197918 -800 198030 480 0 FreeSans 1120 90 0 0 la_data_out[20]
port 332 nsew signal tristate
flabel metal2 s 201464 -800 201576 480 0 FreeSans 1120 90 0 0 la_data_out[21]
port 333 nsew signal tristate
flabel metal2 s 205010 -800 205122 480 0 FreeSans 1120 90 0 0 la_data_out[22]
port 334 nsew signal tristate
flabel metal2 s 208556 -800 208668 480 0 FreeSans 1120 90 0 0 la_data_out[23]
port 335 nsew signal tristate
flabel metal2 s 212102 -800 212214 480 0 FreeSans 1120 90 0 0 la_data_out[24]
port 336 nsew signal tristate
flabel metal2 s 215648 -800 215760 480 0 FreeSans 1120 90 0 0 la_data_out[25]
port 337 nsew signal tristate
flabel metal2 s 219194 -800 219306 480 0 FreeSans 1120 90 0 0 la_data_out[26]
port 338 nsew signal tristate
flabel metal2 s 222740 -800 222852 480 0 FreeSans 1120 90 0 0 la_data_out[27]
port 339 nsew signal tristate
flabel metal2 s 226286 -800 226398 480 0 FreeSans 1120 90 0 0 la_data_out[28]
port 340 nsew signal tristate
flabel metal2 s 229832 -800 229944 480 0 FreeSans 1120 90 0 0 la_data_out[29]
port 341 nsew signal tristate
flabel metal2 s 134090 -800 134202 480 0 FreeSans 1120 90 0 0 la_data_out[2]
port 342 nsew signal tristate
flabel metal2 s 233378 -800 233490 480 0 FreeSans 1120 90 0 0 la_data_out[30]
port 343 nsew signal tristate
flabel metal2 s 236924 -800 237036 480 0 FreeSans 1120 90 0 0 la_data_out[31]
port 344 nsew signal tristate
flabel metal2 s 240470 -800 240582 480 0 FreeSans 1120 90 0 0 la_data_out[32]
port 345 nsew signal tristate
flabel metal2 s 244016 -800 244128 480 0 FreeSans 1120 90 0 0 la_data_out[33]
port 346 nsew signal tristate
flabel metal2 s 247562 -800 247674 480 0 FreeSans 1120 90 0 0 la_data_out[34]
port 347 nsew signal tristate
flabel metal2 s 251108 -800 251220 480 0 FreeSans 1120 90 0 0 la_data_out[35]
port 348 nsew signal tristate
flabel metal2 s 254654 -800 254766 480 0 FreeSans 1120 90 0 0 la_data_out[36]
port 349 nsew signal tristate
flabel metal2 s 258200 -800 258312 480 0 FreeSans 1120 90 0 0 la_data_out[37]
port 350 nsew signal tristate
flabel metal2 s 261746 -800 261858 480 0 FreeSans 1120 90 0 0 la_data_out[38]
port 351 nsew signal tristate
flabel metal2 s 265292 -800 265404 480 0 FreeSans 1120 90 0 0 la_data_out[39]
port 352 nsew signal tristate
flabel metal2 s 137636 -800 137748 480 0 FreeSans 1120 90 0 0 la_data_out[3]
port 353 nsew signal tristate
flabel metal2 s 268838 -800 268950 480 0 FreeSans 1120 90 0 0 la_data_out[40]
port 354 nsew signal tristate
flabel metal2 s 272384 -800 272496 480 0 FreeSans 1120 90 0 0 la_data_out[41]
port 355 nsew signal tristate
flabel metal2 s 275930 -800 276042 480 0 FreeSans 1120 90 0 0 la_data_out[42]
port 356 nsew signal tristate
flabel metal2 s 279476 -800 279588 480 0 FreeSans 1120 90 0 0 la_data_out[43]
port 357 nsew signal tristate
flabel metal2 s 283022 -800 283134 480 0 FreeSans 1120 90 0 0 la_data_out[44]
port 358 nsew signal tristate
flabel metal2 s 286568 -800 286680 480 0 FreeSans 1120 90 0 0 la_data_out[45]
port 359 nsew signal tristate
flabel metal2 s 290114 -800 290226 480 0 FreeSans 1120 90 0 0 la_data_out[46]
port 360 nsew signal tristate
flabel metal2 s 293660 -800 293772 480 0 FreeSans 1120 90 0 0 la_data_out[47]
port 361 nsew signal tristate
flabel metal2 s 297206 -800 297318 480 0 FreeSans 1120 90 0 0 la_data_out[48]
port 362 nsew signal tristate
flabel metal2 s 300752 -800 300864 480 0 FreeSans 1120 90 0 0 la_data_out[49]
port 363 nsew signal tristate
flabel metal2 s 141182 -800 141294 480 0 FreeSans 1120 90 0 0 la_data_out[4]
port 364 nsew signal tristate
flabel metal2 s 304298 -800 304410 480 0 FreeSans 1120 90 0 0 la_data_out[50]
port 365 nsew signal tristate
flabel metal2 s 307844 -800 307956 480 0 FreeSans 1120 90 0 0 la_data_out[51]
port 366 nsew signal tristate
flabel metal2 s 311390 -800 311502 480 0 FreeSans 1120 90 0 0 la_data_out[52]
port 367 nsew signal tristate
flabel metal2 s 314936 -800 315048 480 0 FreeSans 1120 90 0 0 la_data_out[53]
port 368 nsew signal tristate
flabel metal2 s 318482 -800 318594 480 0 FreeSans 1120 90 0 0 la_data_out[54]
port 369 nsew signal tristate
flabel metal2 s 322028 -800 322140 480 0 FreeSans 1120 90 0 0 la_data_out[55]
port 370 nsew signal tristate
flabel metal2 s 325574 -800 325686 480 0 FreeSans 1120 90 0 0 la_data_out[56]
port 371 nsew signal tristate
flabel metal2 s 329120 -800 329232 480 0 FreeSans 1120 90 0 0 la_data_out[57]
port 372 nsew signal tristate
flabel metal2 s 332666 -800 332778 480 0 FreeSans 1120 90 0 0 la_data_out[58]
port 373 nsew signal tristate
flabel metal2 s 336212 -800 336324 480 0 FreeSans 1120 90 0 0 la_data_out[59]
port 374 nsew signal tristate
flabel metal2 s 144728 -800 144840 480 0 FreeSans 1120 90 0 0 la_data_out[5]
port 375 nsew signal tristate
flabel metal2 s 339758 -800 339870 480 0 FreeSans 1120 90 0 0 la_data_out[60]
port 376 nsew signal tristate
flabel metal2 s 343304 -800 343416 480 0 FreeSans 1120 90 0 0 la_data_out[61]
port 377 nsew signal tristate
flabel metal2 s 346850 -800 346962 480 0 FreeSans 1120 90 0 0 la_data_out[62]
port 378 nsew signal tristate
flabel metal2 s 350396 -800 350508 480 0 FreeSans 1120 90 0 0 la_data_out[63]
port 379 nsew signal tristate
flabel metal2 s 353942 -800 354054 480 0 FreeSans 1120 90 0 0 la_data_out[64]
port 380 nsew signal tristate
flabel metal2 s 357488 -800 357600 480 0 FreeSans 1120 90 0 0 la_data_out[65]
port 381 nsew signal tristate
flabel metal2 s 361034 -800 361146 480 0 FreeSans 1120 90 0 0 la_data_out[66]
port 382 nsew signal tristate
flabel metal2 s 364580 -800 364692 480 0 FreeSans 1120 90 0 0 la_data_out[67]
port 383 nsew signal tristate
flabel metal2 s 368126 -800 368238 480 0 FreeSans 1120 90 0 0 la_data_out[68]
port 384 nsew signal tristate
flabel metal2 s 371672 -800 371784 480 0 FreeSans 1120 90 0 0 la_data_out[69]
port 385 nsew signal tristate
flabel metal2 s 148274 -800 148386 480 0 FreeSans 1120 90 0 0 la_data_out[6]
port 386 nsew signal tristate
flabel metal2 s 375218 -800 375330 480 0 FreeSans 1120 90 0 0 la_data_out[70]
port 387 nsew signal tristate
flabel metal2 s 378764 -800 378876 480 0 FreeSans 1120 90 0 0 la_data_out[71]
port 388 nsew signal tristate
flabel metal2 s 382310 -800 382422 480 0 FreeSans 1120 90 0 0 la_data_out[72]
port 389 nsew signal tristate
flabel metal2 s 385856 -800 385968 480 0 FreeSans 1120 90 0 0 la_data_out[73]
port 390 nsew signal tristate
flabel metal2 s 389402 -800 389514 480 0 FreeSans 1120 90 0 0 la_data_out[74]
port 391 nsew signal tristate
flabel metal2 s 392948 -800 393060 480 0 FreeSans 1120 90 0 0 la_data_out[75]
port 392 nsew signal tristate
flabel metal2 s 396494 -800 396606 480 0 FreeSans 1120 90 0 0 la_data_out[76]
port 393 nsew signal tristate
flabel metal2 s 400040 -800 400152 480 0 FreeSans 1120 90 0 0 la_data_out[77]
port 394 nsew signal tristate
flabel metal2 s 403586 -800 403698 480 0 FreeSans 1120 90 0 0 la_data_out[78]
port 395 nsew signal tristate
flabel metal2 s 407132 -800 407244 480 0 FreeSans 1120 90 0 0 la_data_out[79]
port 396 nsew signal tristate
flabel metal2 s 151820 -800 151932 480 0 FreeSans 1120 90 0 0 la_data_out[7]
port 397 nsew signal tristate
flabel metal2 s 410678 -800 410790 480 0 FreeSans 1120 90 0 0 la_data_out[80]
port 398 nsew signal tristate
flabel metal2 s 414224 -800 414336 480 0 FreeSans 1120 90 0 0 la_data_out[81]
port 399 nsew signal tristate
flabel metal2 s 417770 -800 417882 480 0 FreeSans 1120 90 0 0 la_data_out[82]
port 400 nsew signal tristate
flabel metal2 s 421316 -800 421428 480 0 FreeSans 1120 90 0 0 la_data_out[83]
port 401 nsew signal tristate
flabel metal2 s 424862 -800 424974 480 0 FreeSans 1120 90 0 0 la_data_out[84]
port 402 nsew signal tristate
flabel metal2 s 428408 -800 428520 480 0 FreeSans 1120 90 0 0 la_data_out[85]
port 403 nsew signal tristate
flabel metal2 s 431954 -800 432066 480 0 FreeSans 1120 90 0 0 la_data_out[86]
port 404 nsew signal tristate
flabel metal2 s 435500 -800 435612 480 0 FreeSans 1120 90 0 0 la_data_out[87]
port 405 nsew signal tristate
flabel metal2 s 439046 -800 439158 480 0 FreeSans 1120 90 0 0 la_data_out[88]
port 406 nsew signal tristate
flabel metal2 s 442592 -800 442704 480 0 FreeSans 1120 90 0 0 la_data_out[89]
port 407 nsew signal tristate
flabel metal2 s 155366 -800 155478 480 0 FreeSans 1120 90 0 0 la_data_out[8]
port 408 nsew signal tristate
flabel metal2 s 446138 -800 446250 480 0 FreeSans 1120 90 0 0 la_data_out[90]
port 409 nsew signal tristate
flabel metal2 s 449684 -800 449796 480 0 FreeSans 1120 90 0 0 la_data_out[91]
port 410 nsew signal tristate
flabel metal2 s 453230 -800 453342 480 0 FreeSans 1120 90 0 0 la_data_out[92]
port 411 nsew signal tristate
flabel metal2 s 456776 -800 456888 480 0 FreeSans 1120 90 0 0 la_data_out[93]
port 412 nsew signal tristate
flabel metal2 s 460322 -800 460434 480 0 FreeSans 1120 90 0 0 la_data_out[94]
port 413 nsew signal tristate
flabel metal2 s 463868 -800 463980 480 0 FreeSans 1120 90 0 0 la_data_out[95]
port 414 nsew signal tristate
flabel metal2 s 467414 -800 467526 480 0 FreeSans 1120 90 0 0 la_data_out[96]
port 415 nsew signal tristate
flabel metal2 s 470960 -800 471072 480 0 FreeSans 1120 90 0 0 la_data_out[97]
port 416 nsew signal tristate
flabel metal2 s 474506 -800 474618 480 0 FreeSans 1120 90 0 0 la_data_out[98]
port 417 nsew signal tristate
flabel metal2 s 478052 -800 478164 480 0 FreeSans 1120 90 0 0 la_data_out[99]
port 418 nsew signal tristate
flabel metal2 s 158912 -800 159024 480 0 FreeSans 1120 90 0 0 la_data_out[9]
port 419 nsew signal tristate
flabel metal2 s 128180 -800 128292 480 0 FreeSans 1120 90 0 0 la_oenb[0]
port 420 nsew signal input
flabel metal2 s 482780 -800 482892 480 0 FreeSans 1120 90 0 0 la_oenb[100]
port 421 nsew signal input
flabel metal2 s 486326 -800 486438 480 0 FreeSans 1120 90 0 0 la_oenb[101]
port 422 nsew signal input
flabel metal2 s 489872 -800 489984 480 0 FreeSans 1120 90 0 0 la_oenb[102]
port 423 nsew signal input
flabel metal2 s 493418 -800 493530 480 0 FreeSans 1120 90 0 0 la_oenb[103]
port 424 nsew signal input
flabel metal2 s 496964 -800 497076 480 0 FreeSans 1120 90 0 0 la_oenb[104]
port 425 nsew signal input
flabel metal2 s 500510 -800 500622 480 0 FreeSans 1120 90 0 0 la_oenb[105]
port 426 nsew signal input
flabel metal2 s 504056 -800 504168 480 0 FreeSans 1120 90 0 0 la_oenb[106]
port 427 nsew signal input
flabel metal2 s 507602 -800 507714 480 0 FreeSans 1120 90 0 0 la_oenb[107]
port 428 nsew signal input
flabel metal2 s 511148 -800 511260 480 0 FreeSans 1120 90 0 0 la_oenb[108]
port 429 nsew signal input
flabel metal2 s 514694 -800 514806 480 0 FreeSans 1120 90 0 0 la_oenb[109]
port 430 nsew signal input
flabel metal2 s 163640 -800 163752 480 0 FreeSans 1120 90 0 0 la_oenb[10]
port 431 nsew signal input
flabel metal2 s 518240 -800 518352 480 0 FreeSans 1120 90 0 0 la_oenb[110]
port 432 nsew signal input
flabel metal2 s 521786 -800 521898 480 0 FreeSans 1120 90 0 0 la_oenb[111]
port 433 nsew signal input
flabel metal2 s 525332 -800 525444 480 0 FreeSans 1120 90 0 0 la_oenb[112]
port 434 nsew signal input
flabel metal2 s 528878 -800 528990 480 0 FreeSans 1120 90 0 0 la_oenb[113]
port 435 nsew signal input
flabel metal2 s 532424 -800 532536 480 0 FreeSans 1120 90 0 0 la_oenb[114]
port 436 nsew signal input
flabel metal2 s 535970 -800 536082 480 0 FreeSans 1120 90 0 0 la_oenb[115]
port 437 nsew signal input
flabel metal2 s 539516 -800 539628 480 0 FreeSans 1120 90 0 0 la_oenb[116]
port 438 nsew signal input
flabel metal2 s 543062 -800 543174 480 0 FreeSans 1120 90 0 0 la_oenb[117]
port 439 nsew signal input
flabel metal2 s 546608 -800 546720 480 0 FreeSans 1120 90 0 0 la_oenb[118]
port 440 nsew signal input
flabel metal2 s 550154 -800 550266 480 0 FreeSans 1120 90 0 0 la_oenb[119]
port 441 nsew signal input
flabel metal2 s 167186 -800 167298 480 0 FreeSans 1120 90 0 0 la_oenb[11]
port 442 nsew signal input
flabel metal2 s 553700 -800 553812 480 0 FreeSans 1120 90 0 0 la_oenb[120]
port 443 nsew signal input
flabel metal2 s 557246 -800 557358 480 0 FreeSans 1120 90 0 0 la_oenb[121]
port 444 nsew signal input
flabel metal2 s 560792 -800 560904 480 0 FreeSans 1120 90 0 0 la_oenb[122]
port 445 nsew signal input
flabel metal2 s 564338 -800 564450 480 0 FreeSans 1120 90 0 0 la_oenb[123]
port 446 nsew signal input
flabel metal2 s 567884 -800 567996 480 0 FreeSans 1120 90 0 0 la_oenb[124]
port 447 nsew signal input
flabel metal2 s 571430 -800 571542 480 0 FreeSans 1120 90 0 0 la_oenb[125]
port 448 nsew signal input
flabel metal2 s 574976 -800 575088 480 0 FreeSans 1120 90 0 0 la_oenb[126]
port 449 nsew signal input
flabel metal2 s 578522 -800 578634 480 0 FreeSans 1120 90 0 0 la_oenb[127]
port 450 nsew signal input
flabel metal2 s 170732 -800 170844 480 0 FreeSans 1120 90 0 0 la_oenb[12]
port 451 nsew signal input
flabel metal2 s 174278 -800 174390 480 0 FreeSans 1120 90 0 0 la_oenb[13]
port 452 nsew signal input
flabel metal2 s 177824 -800 177936 480 0 FreeSans 1120 90 0 0 la_oenb[14]
port 453 nsew signal input
flabel metal2 s 181370 -800 181482 480 0 FreeSans 1120 90 0 0 la_oenb[15]
port 454 nsew signal input
flabel metal2 s 184916 -800 185028 480 0 FreeSans 1120 90 0 0 la_oenb[16]
port 455 nsew signal input
flabel metal2 s 188462 -800 188574 480 0 FreeSans 1120 90 0 0 la_oenb[17]
port 456 nsew signal input
flabel metal2 s 192008 -800 192120 480 0 FreeSans 1120 90 0 0 la_oenb[18]
port 457 nsew signal input
flabel metal2 s 195554 -800 195666 480 0 FreeSans 1120 90 0 0 la_oenb[19]
port 458 nsew signal input
flabel metal2 s 131726 -800 131838 480 0 FreeSans 1120 90 0 0 la_oenb[1]
port 459 nsew signal input
flabel metal2 s 199100 -800 199212 480 0 FreeSans 1120 90 0 0 la_oenb[20]
port 460 nsew signal input
flabel metal2 s 202646 -800 202758 480 0 FreeSans 1120 90 0 0 la_oenb[21]
port 461 nsew signal input
flabel metal2 s 206192 -800 206304 480 0 FreeSans 1120 90 0 0 la_oenb[22]
port 462 nsew signal input
flabel metal2 s 209738 -800 209850 480 0 FreeSans 1120 90 0 0 la_oenb[23]
port 463 nsew signal input
flabel metal2 s 213284 -800 213396 480 0 FreeSans 1120 90 0 0 la_oenb[24]
port 464 nsew signal input
flabel metal2 s 216830 -800 216942 480 0 FreeSans 1120 90 0 0 la_oenb[25]
port 465 nsew signal input
flabel metal2 s 220376 -800 220488 480 0 FreeSans 1120 90 0 0 la_oenb[26]
port 466 nsew signal input
flabel metal2 s 223922 -800 224034 480 0 FreeSans 1120 90 0 0 la_oenb[27]
port 467 nsew signal input
flabel metal2 s 227468 -800 227580 480 0 FreeSans 1120 90 0 0 la_oenb[28]
port 468 nsew signal input
flabel metal2 s 231014 -800 231126 480 0 FreeSans 1120 90 0 0 la_oenb[29]
port 469 nsew signal input
flabel metal2 s 135272 -800 135384 480 0 FreeSans 1120 90 0 0 la_oenb[2]
port 470 nsew signal input
flabel metal2 s 234560 -800 234672 480 0 FreeSans 1120 90 0 0 la_oenb[30]
port 471 nsew signal input
flabel metal2 s 238106 -800 238218 480 0 FreeSans 1120 90 0 0 la_oenb[31]
port 472 nsew signal input
flabel metal2 s 241652 -800 241764 480 0 FreeSans 1120 90 0 0 la_oenb[32]
port 473 nsew signal input
flabel metal2 s 245198 -800 245310 480 0 FreeSans 1120 90 0 0 la_oenb[33]
port 474 nsew signal input
flabel metal2 s 248744 -800 248856 480 0 FreeSans 1120 90 0 0 la_oenb[34]
port 475 nsew signal input
flabel metal2 s 252290 -800 252402 480 0 FreeSans 1120 90 0 0 la_oenb[35]
port 476 nsew signal input
flabel metal2 s 255836 -800 255948 480 0 FreeSans 1120 90 0 0 la_oenb[36]
port 477 nsew signal input
flabel metal2 s 259382 -800 259494 480 0 FreeSans 1120 90 0 0 la_oenb[37]
port 478 nsew signal input
flabel metal2 s 262928 -800 263040 480 0 FreeSans 1120 90 0 0 la_oenb[38]
port 479 nsew signal input
flabel metal2 s 266474 -800 266586 480 0 FreeSans 1120 90 0 0 la_oenb[39]
port 480 nsew signal input
flabel metal2 s 138818 -800 138930 480 0 FreeSans 1120 90 0 0 la_oenb[3]
port 481 nsew signal input
flabel metal2 s 270020 -800 270132 480 0 FreeSans 1120 90 0 0 la_oenb[40]
port 482 nsew signal input
flabel metal2 s 273566 -800 273678 480 0 FreeSans 1120 90 0 0 la_oenb[41]
port 483 nsew signal input
flabel metal2 s 277112 -800 277224 480 0 FreeSans 1120 90 0 0 la_oenb[42]
port 484 nsew signal input
flabel metal2 s 280658 -800 280770 480 0 FreeSans 1120 90 0 0 la_oenb[43]
port 485 nsew signal input
flabel metal2 s 284204 -800 284316 480 0 FreeSans 1120 90 0 0 la_oenb[44]
port 486 nsew signal input
flabel metal2 s 287750 -800 287862 480 0 FreeSans 1120 90 0 0 la_oenb[45]
port 487 nsew signal input
flabel metal2 s 291296 -800 291408 480 0 FreeSans 1120 90 0 0 la_oenb[46]
port 488 nsew signal input
flabel metal2 s 294842 -800 294954 480 0 FreeSans 1120 90 0 0 la_oenb[47]
port 489 nsew signal input
flabel metal2 s 298388 -800 298500 480 0 FreeSans 1120 90 0 0 la_oenb[48]
port 490 nsew signal input
flabel metal2 s 301934 -800 302046 480 0 FreeSans 1120 90 0 0 la_oenb[49]
port 491 nsew signal input
flabel metal2 s 142364 -800 142476 480 0 FreeSans 1120 90 0 0 la_oenb[4]
port 492 nsew signal input
flabel metal2 s 305480 -800 305592 480 0 FreeSans 1120 90 0 0 la_oenb[50]
port 493 nsew signal input
flabel metal2 s 309026 -800 309138 480 0 FreeSans 1120 90 0 0 la_oenb[51]
port 494 nsew signal input
flabel metal2 s 312572 -800 312684 480 0 FreeSans 1120 90 0 0 la_oenb[52]
port 495 nsew signal input
flabel metal2 s 316118 -800 316230 480 0 FreeSans 1120 90 0 0 la_oenb[53]
port 496 nsew signal input
flabel metal2 s 319664 -800 319776 480 0 FreeSans 1120 90 0 0 la_oenb[54]
port 497 nsew signal input
flabel metal2 s 323210 -800 323322 480 0 FreeSans 1120 90 0 0 la_oenb[55]
port 498 nsew signal input
flabel metal2 s 326756 -800 326868 480 0 FreeSans 1120 90 0 0 la_oenb[56]
port 499 nsew signal input
flabel metal2 s 330302 -800 330414 480 0 FreeSans 1120 90 0 0 la_oenb[57]
port 500 nsew signal input
flabel metal2 s 333848 -800 333960 480 0 FreeSans 1120 90 0 0 la_oenb[58]
port 501 nsew signal input
flabel metal2 s 337394 -800 337506 480 0 FreeSans 1120 90 0 0 la_oenb[59]
port 502 nsew signal input
flabel metal2 s 145910 -800 146022 480 0 FreeSans 1120 90 0 0 la_oenb[5]
port 503 nsew signal input
flabel metal2 s 340940 -800 341052 480 0 FreeSans 1120 90 0 0 la_oenb[60]
port 504 nsew signal input
flabel metal2 s 344486 -800 344598 480 0 FreeSans 1120 90 0 0 la_oenb[61]
port 505 nsew signal input
flabel metal2 s 348032 -800 348144 480 0 FreeSans 1120 90 0 0 la_oenb[62]
port 506 nsew signal input
flabel metal2 s 351578 -800 351690 480 0 FreeSans 1120 90 0 0 la_oenb[63]
port 507 nsew signal input
flabel metal2 s 355124 -800 355236 480 0 FreeSans 1120 90 0 0 la_oenb[64]
port 508 nsew signal input
flabel metal2 s 358670 -800 358782 480 0 FreeSans 1120 90 0 0 la_oenb[65]
port 509 nsew signal input
flabel metal2 s 362216 -800 362328 480 0 FreeSans 1120 90 0 0 la_oenb[66]
port 510 nsew signal input
flabel metal2 s 365762 -800 365874 480 0 FreeSans 1120 90 0 0 la_oenb[67]
port 511 nsew signal input
flabel metal2 s 369308 -800 369420 480 0 FreeSans 1120 90 0 0 la_oenb[68]
port 512 nsew signal input
flabel metal2 s 372854 -800 372966 480 0 FreeSans 1120 90 0 0 la_oenb[69]
port 513 nsew signal input
flabel metal2 s 149456 -800 149568 480 0 FreeSans 1120 90 0 0 la_oenb[6]
port 514 nsew signal input
flabel metal2 s 376400 -800 376512 480 0 FreeSans 1120 90 0 0 la_oenb[70]
port 515 nsew signal input
flabel metal2 s 379946 -800 380058 480 0 FreeSans 1120 90 0 0 la_oenb[71]
port 516 nsew signal input
flabel metal2 s 383492 -800 383604 480 0 FreeSans 1120 90 0 0 la_oenb[72]
port 517 nsew signal input
flabel metal2 s 387038 -800 387150 480 0 FreeSans 1120 90 0 0 la_oenb[73]
port 518 nsew signal input
flabel metal2 s 390584 -800 390696 480 0 FreeSans 1120 90 0 0 la_oenb[74]
port 519 nsew signal input
flabel metal2 s 394130 -800 394242 480 0 FreeSans 1120 90 0 0 la_oenb[75]
port 520 nsew signal input
flabel metal2 s 397676 -800 397788 480 0 FreeSans 1120 90 0 0 la_oenb[76]
port 521 nsew signal input
flabel metal2 s 401222 -800 401334 480 0 FreeSans 1120 90 0 0 la_oenb[77]
port 522 nsew signal input
flabel metal2 s 404768 -800 404880 480 0 FreeSans 1120 90 0 0 la_oenb[78]
port 523 nsew signal input
flabel metal2 s 408314 -800 408426 480 0 FreeSans 1120 90 0 0 la_oenb[79]
port 524 nsew signal input
flabel metal2 s 153002 -800 153114 480 0 FreeSans 1120 90 0 0 la_oenb[7]
port 525 nsew signal input
flabel metal2 s 411860 -800 411972 480 0 FreeSans 1120 90 0 0 la_oenb[80]
port 526 nsew signal input
flabel metal2 s 415406 -800 415518 480 0 FreeSans 1120 90 0 0 la_oenb[81]
port 527 nsew signal input
flabel metal2 s 418952 -800 419064 480 0 FreeSans 1120 90 0 0 la_oenb[82]
port 528 nsew signal input
flabel metal2 s 422498 -800 422610 480 0 FreeSans 1120 90 0 0 la_oenb[83]
port 529 nsew signal input
flabel metal2 s 426044 -800 426156 480 0 FreeSans 1120 90 0 0 la_oenb[84]
port 530 nsew signal input
flabel metal2 s 429590 -800 429702 480 0 FreeSans 1120 90 0 0 la_oenb[85]
port 531 nsew signal input
flabel metal2 s 433136 -800 433248 480 0 FreeSans 1120 90 0 0 la_oenb[86]
port 532 nsew signal input
flabel metal2 s 436682 -800 436794 480 0 FreeSans 1120 90 0 0 la_oenb[87]
port 533 nsew signal input
flabel metal2 s 440228 -800 440340 480 0 FreeSans 1120 90 0 0 la_oenb[88]
port 534 nsew signal input
flabel metal2 s 443774 -800 443886 480 0 FreeSans 1120 90 0 0 la_oenb[89]
port 535 nsew signal input
flabel metal2 s 156548 -800 156660 480 0 FreeSans 1120 90 0 0 la_oenb[8]
port 536 nsew signal input
flabel metal2 s 447320 -800 447432 480 0 FreeSans 1120 90 0 0 la_oenb[90]
port 537 nsew signal input
flabel metal2 s 450866 -800 450978 480 0 FreeSans 1120 90 0 0 la_oenb[91]
port 538 nsew signal input
flabel metal2 s 454412 -800 454524 480 0 FreeSans 1120 90 0 0 la_oenb[92]
port 539 nsew signal input
flabel metal2 s 457958 -800 458070 480 0 FreeSans 1120 90 0 0 la_oenb[93]
port 540 nsew signal input
flabel metal2 s 461504 -800 461616 480 0 FreeSans 1120 90 0 0 la_oenb[94]
port 541 nsew signal input
flabel metal2 s 465050 -800 465162 480 0 FreeSans 1120 90 0 0 la_oenb[95]
port 542 nsew signal input
flabel metal2 s 468596 -800 468708 480 0 FreeSans 1120 90 0 0 la_oenb[96]
port 543 nsew signal input
flabel metal2 s 472142 -800 472254 480 0 FreeSans 1120 90 0 0 la_oenb[97]
port 544 nsew signal input
flabel metal2 s 475688 -800 475800 480 0 FreeSans 1120 90 0 0 la_oenb[98]
port 545 nsew signal input
flabel metal2 s 479234 -800 479346 480 0 FreeSans 1120 90 0 0 la_oenb[99]
port 546 nsew signal input
flabel metal2 s 160094 -800 160206 480 0 FreeSans 1120 90 0 0 la_oenb[9]
port 547 nsew signal input
flabel metal2 s 579704 -800 579816 480 0 FreeSans 1120 90 0 0 user_clock2
port 548 nsew signal input
flabel metal2 s 580886 -800 580998 480 0 FreeSans 1120 90 0 0 user_irq[0]
port 549 nsew signal tristate
flabel metal2 s 582068 -800 582180 480 0 FreeSans 1120 90 0 0 user_irq[1]
port 550 nsew signal tristate
flabel metal2 s 583250 -800 583362 480 0 FreeSans 1120 90 0 0 user_irq[2]
port 551 nsew signal tristate
flabel metal3 s 582340 639784 584800 644584 0 FreeSans 1120 0 0 0 vccd1
port 552 nsew signal bidirectional
flabel metal3 s 582340 629784 584800 634584 0 FreeSans 1120 0 0 0 vccd1
port 553 nsew signal bidirectional
flabel metal3 s 0 643842 1660 648642 0 FreeSans 1120 0 0 0 vccd2
port 554 nsew signal bidirectional
flabel metal3 s 0 633842 1660 638642 0 FreeSans 1120 0 0 0 vccd2
port 555 nsew signal bidirectional
flabel metal3 s 582340 540562 584800 545362 0 FreeSans 1120 0 0 0 vdda1
port 556 nsew signal bidirectional
flabel metal3 s 582340 550562 584800 555362 0 FreeSans 1120 0 0 0 vdda1
port 557 nsew signal bidirectional
flabel metal3 s 582340 235230 584800 240030 0 FreeSans 1120 0 0 0 vdda1
port 558 nsew signal bidirectional
flabel metal3 s 582340 225230 584800 230030 0 FreeSans 1120 0 0 0 vdda1
port 559 nsew signal bidirectional
flabel metal3 s 0 204888 1660 209688 0 FreeSans 1120 0 0 0 vdda2
port 560 nsew signal bidirectional
flabel metal3 s 0 214888 1660 219688 0 FreeSans 1120 0 0 0 vdda2
port 561 nsew signal bidirectional
flabel metal3 s 520594 702340 525394 704800 0 FreeSans 1920 180 0 0 vssa1
port 562 nsew signal bidirectional
flabel metal3 s 510594 702340 515394 704800 0 FreeSans 1920 180 0 0 vssa1
port 563 nsew signal bidirectional
flabel metal3 s 582340 146830 584800 151630 0 FreeSans 1120 0 0 0 vssa1
port 564 nsew signal bidirectional
flabel metal3 s 582340 136830 584800 141630 0 FreeSans 1120 0 0 0 vssa1
port 565 nsew signal bidirectional
flabel metal3 s 0 559442 1660 564242 0 FreeSans 1120 0 0 0 vssa2
port 566 nsew signal bidirectional
flabel metal3 s 0 549442 1660 554242 0 FreeSans 1120 0 0 0 vssa2
port 567 nsew signal bidirectional
flabel metal3 s 582340 191430 584800 196230 0 FreeSans 1120 0 0 0 vssd1
port 568 nsew signal bidirectional
flabel metal3 s 582340 181430 584800 186230 0 FreeSans 1120 0 0 0 vssd1
port 569 nsew signal bidirectional
flabel metal3 s 0 172888 1660 177688 0 FreeSans 1120 0 0 0 vssd2
port 570 nsew signal bidirectional
flabel metal3 s 0 162888 1660 167688 0 FreeSans 1120 0 0 0 vssd2
port 571 nsew signal bidirectional
flabel metal2 s 524 -800 636 480 0 FreeSans 1120 90 0 0 wb_clk_i
port 572 nsew signal input
flabel metal2 s 1706 -800 1818 480 0 FreeSans 1120 90 0 0 wb_rst_i
port 573 nsew signal input
flabel metal2 s 2888 -800 3000 480 0 FreeSans 1120 90 0 0 wbs_ack_o
port 574 nsew signal tristate
flabel metal2 s 7616 -800 7728 480 0 FreeSans 1120 90 0 0 wbs_adr_i[0]
port 575 nsew signal input
flabel metal2 s 47804 -800 47916 480 0 FreeSans 1120 90 0 0 wbs_adr_i[10]
port 576 nsew signal input
flabel metal2 s 51350 -800 51462 480 0 FreeSans 1120 90 0 0 wbs_adr_i[11]
port 577 nsew signal input
flabel metal2 s 54896 -800 55008 480 0 FreeSans 1120 90 0 0 wbs_adr_i[12]
port 578 nsew signal input
flabel metal2 s 58442 -800 58554 480 0 FreeSans 1120 90 0 0 wbs_adr_i[13]
port 579 nsew signal input
flabel metal2 s 61988 -800 62100 480 0 FreeSans 1120 90 0 0 wbs_adr_i[14]
port 580 nsew signal input
flabel metal2 s 65534 -800 65646 480 0 FreeSans 1120 90 0 0 wbs_adr_i[15]
port 581 nsew signal input
flabel metal2 s 69080 -800 69192 480 0 FreeSans 1120 90 0 0 wbs_adr_i[16]
port 582 nsew signal input
flabel metal2 s 72626 -800 72738 480 0 FreeSans 1120 90 0 0 wbs_adr_i[17]
port 583 nsew signal input
flabel metal2 s 76172 -800 76284 480 0 FreeSans 1120 90 0 0 wbs_adr_i[18]
port 584 nsew signal input
flabel metal2 s 79718 -800 79830 480 0 FreeSans 1120 90 0 0 wbs_adr_i[19]
port 585 nsew signal input
flabel metal2 s 12344 -800 12456 480 0 FreeSans 1120 90 0 0 wbs_adr_i[1]
port 586 nsew signal input
flabel metal2 s 83264 -800 83376 480 0 FreeSans 1120 90 0 0 wbs_adr_i[20]
port 587 nsew signal input
flabel metal2 s 86810 -800 86922 480 0 FreeSans 1120 90 0 0 wbs_adr_i[21]
port 588 nsew signal input
flabel metal2 s 90356 -800 90468 480 0 FreeSans 1120 90 0 0 wbs_adr_i[22]
port 589 nsew signal input
flabel metal2 s 93902 -800 94014 480 0 FreeSans 1120 90 0 0 wbs_adr_i[23]
port 590 nsew signal input
flabel metal2 s 97448 -800 97560 480 0 FreeSans 1120 90 0 0 wbs_adr_i[24]
port 591 nsew signal input
flabel metal2 s 100994 -800 101106 480 0 FreeSans 1120 90 0 0 wbs_adr_i[25]
port 592 nsew signal input
flabel metal2 s 104540 -800 104652 480 0 FreeSans 1120 90 0 0 wbs_adr_i[26]
port 593 nsew signal input
flabel metal2 s 108086 -800 108198 480 0 FreeSans 1120 90 0 0 wbs_adr_i[27]
port 594 nsew signal input
flabel metal2 s 111632 -800 111744 480 0 FreeSans 1120 90 0 0 wbs_adr_i[28]
port 595 nsew signal input
flabel metal2 s 115178 -800 115290 480 0 FreeSans 1120 90 0 0 wbs_adr_i[29]
port 596 nsew signal input
flabel metal2 s 17072 -800 17184 480 0 FreeSans 1120 90 0 0 wbs_adr_i[2]
port 597 nsew signal input
flabel metal2 s 118724 -800 118836 480 0 FreeSans 1120 90 0 0 wbs_adr_i[30]
port 598 nsew signal input
flabel metal2 s 122270 -800 122382 480 0 FreeSans 1120 90 0 0 wbs_adr_i[31]
port 599 nsew signal input
flabel metal2 s 21800 -800 21912 480 0 FreeSans 1120 90 0 0 wbs_adr_i[3]
port 600 nsew signal input
flabel metal2 s 26528 -800 26640 480 0 FreeSans 1120 90 0 0 wbs_adr_i[4]
port 601 nsew signal input
flabel metal2 s 30074 -800 30186 480 0 FreeSans 1120 90 0 0 wbs_adr_i[5]
port 602 nsew signal input
flabel metal2 s 33620 -800 33732 480 0 FreeSans 1120 90 0 0 wbs_adr_i[6]
port 603 nsew signal input
flabel metal2 s 37166 -800 37278 480 0 FreeSans 1120 90 0 0 wbs_adr_i[7]
port 604 nsew signal input
flabel metal2 s 40712 -800 40824 480 0 FreeSans 1120 90 0 0 wbs_adr_i[8]
port 605 nsew signal input
flabel metal2 s 44258 -800 44370 480 0 FreeSans 1120 90 0 0 wbs_adr_i[9]
port 606 nsew signal input
flabel metal2 s 4070 -800 4182 480 0 FreeSans 1120 90 0 0 wbs_cyc_i
port 607 nsew signal input
flabel metal2 s 8798 -800 8910 480 0 FreeSans 1120 90 0 0 wbs_dat_i[0]
port 608 nsew signal input
flabel metal2 s 48986 -800 49098 480 0 FreeSans 1120 90 0 0 wbs_dat_i[10]
port 609 nsew signal input
flabel metal2 s 52532 -800 52644 480 0 FreeSans 1120 90 0 0 wbs_dat_i[11]
port 610 nsew signal input
flabel metal2 s 56078 -800 56190 480 0 FreeSans 1120 90 0 0 wbs_dat_i[12]
port 611 nsew signal input
flabel metal2 s 59624 -800 59736 480 0 FreeSans 1120 90 0 0 wbs_dat_i[13]
port 612 nsew signal input
flabel metal2 s 63170 -800 63282 480 0 FreeSans 1120 90 0 0 wbs_dat_i[14]
port 613 nsew signal input
flabel metal2 s 66716 -800 66828 480 0 FreeSans 1120 90 0 0 wbs_dat_i[15]
port 614 nsew signal input
flabel metal2 s 70262 -800 70374 480 0 FreeSans 1120 90 0 0 wbs_dat_i[16]
port 615 nsew signal input
flabel metal2 s 73808 -800 73920 480 0 FreeSans 1120 90 0 0 wbs_dat_i[17]
port 616 nsew signal input
flabel metal2 s 77354 -800 77466 480 0 FreeSans 1120 90 0 0 wbs_dat_i[18]
port 617 nsew signal input
flabel metal2 s 80900 -800 81012 480 0 FreeSans 1120 90 0 0 wbs_dat_i[19]
port 618 nsew signal input
flabel metal2 s 13526 -800 13638 480 0 FreeSans 1120 90 0 0 wbs_dat_i[1]
port 619 nsew signal input
flabel metal2 s 84446 -800 84558 480 0 FreeSans 1120 90 0 0 wbs_dat_i[20]
port 620 nsew signal input
flabel metal2 s 87992 -800 88104 480 0 FreeSans 1120 90 0 0 wbs_dat_i[21]
port 621 nsew signal input
flabel metal2 s 91538 -800 91650 480 0 FreeSans 1120 90 0 0 wbs_dat_i[22]
port 622 nsew signal input
flabel metal2 s 95084 -800 95196 480 0 FreeSans 1120 90 0 0 wbs_dat_i[23]
port 623 nsew signal input
flabel metal2 s 98630 -800 98742 480 0 FreeSans 1120 90 0 0 wbs_dat_i[24]
port 624 nsew signal input
flabel metal2 s 102176 -800 102288 480 0 FreeSans 1120 90 0 0 wbs_dat_i[25]
port 625 nsew signal input
flabel metal2 s 105722 -800 105834 480 0 FreeSans 1120 90 0 0 wbs_dat_i[26]
port 626 nsew signal input
flabel metal2 s 109268 -800 109380 480 0 FreeSans 1120 90 0 0 wbs_dat_i[27]
port 627 nsew signal input
flabel metal2 s 112814 -800 112926 480 0 FreeSans 1120 90 0 0 wbs_dat_i[28]
port 628 nsew signal input
flabel metal2 s 116360 -800 116472 480 0 FreeSans 1120 90 0 0 wbs_dat_i[29]
port 629 nsew signal input
flabel metal2 s 18254 -800 18366 480 0 FreeSans 1120 90 0 0 wbs_dat_i[2]
port 630 nsew signal input
flabel metal2 s 119906 -800 120018 480 0 FreeSans 1120 90 0 0 wbs_dat_i[30]
port 631 nsew signal input
flabel metal2 s 123452 -800 123564 480 0 FreeSans 1120 90 0 0 wbs_dat_i[31]
port 632 nsew signal input
flabel metal2 s 22982 -800 23094 480 0 FreeSans 1120 90 0 0 wbs_dat_i[3]
port 633 nsew signal input
flabel metal2 s 27710 -800 27822 480 0 FreeSans 1120 90 0 0 wbs_dat_i[4]
port 634 nsew signal input
flabel metal2 s 31256 -800 31368 480 0 FreeSans 1120 90 0 0 wbs_dat_i[5]
port 635 nsew signal input
flabel metal2 s 34802 -800 34914 480 0 FreeSans 1120 90 0 0 wbs_dat_i[6]
port 636 nsew signal input
flabel metal2 s 38348 -800 38460 480 0 FreeSans 1120 90 0 0 wbs_dat_i[7]
port 637 nsew signal input
flabel metal2 s 41894 -800 42006 480 0 FreeSans 1120 90 0 0 wbs_dat_i[8]
port 638 nsew signal input
flabel metal2 s 45440 -800 45552 480 0 FreeSans 1120 90 0 0 wbs_dat_i[9]
port 639 nsew signal input
flabel metal2 s 9980 -800 10092 480 0 FreeSans 1120 90 0 0 wbs_dat_o[0]
port 640 nsew signal tristate
flabel metal2 s 50168 -800 50280 480 0 FreeSans 1120 90 0 0 wbs_dat_o[10]
port 641 nsew signal tristate
flabel metal2 s 53714 -800 53826 480 0 FreeSans 1120 90 0 0 wbs_dat_o[11]
port 642 nsew signal tristate
flabel metal2 s 57260 -800 57372 480 0 FreeSans 1120 90 0 0 wbs_dat_o[12]
port 643 nsew signal tristate
flabel metal2 s 60806 -800 60918 480 0 FreeSans 1120 90 0 0 wbs_dat_o[13]
port 644 nsew signal tristate
flabel metal2 s 64352 -800 64464 480 0 FreeSans 1120 90 0 0 wbs_dat_o[14]
port 645 nsew signal tristate
flabel metal2 s 67898 -800 68010 480 0 FreeSans 1120 90 0 0 wbs_dat_o[15]
port 646 nsew signal tristate
flabel metal2 s 71444 -800 71556 480 0 FreeSans 1120 90 0 0 wbs_dat_o[16]
port 647 nsew signal tristate
flabel metal2 s 74990 -800 75102 480 0 FreeSans 1120 90 0 0 wbs_dat_o[17]
port 648 nsew signal tristate
flabel metal2 s 78536 -800 78648 480 0 FreeSans 1120 90 0 0 wbs_dat_o[18]
port 649 nsew signal tristate
flabel metal2 s 82082 -800 82194 480 0 FreeSans 1120 90 0 0 wbs_dat_o[19]
port 650 nsew signal tristate
flabel metal2 s 14708 -800 14820 480 0 FreeSans 1120 90 0 0 wbs_dat_o[1]
port 651 nsew signal tristate
flabel metal2 s 85628 -800 85740 480 0 FreeSans 1120 90 0 0 wbs_dat_o[20]
port 652 nsew signal tristate
flabel metal2 s 89174 -800 89286 480 0 FreeSans 1120 90 0 0 wbs_dat_o[21]
port 653 nsew signal tristate
flabel metal2 s 92720 -800 92832 480 0 FreeSans 1120 90 0 0 wbs_dat_o[22]
port 654 nsew signal tristate
flabel metal2 s 96266 -800 96378 480 0 FreeSans 1120 90 0 0 wbs_dat_o[23]
port 655 nsew signal tristate
flabel metal2 s 99812 -800 99924 480 0 FreeSans 1120 90 0 0 wbs_dat_o[24]
port 656 nsew signal tristate
flabel metal2 s 103358 -800 103470 480 0 FreeSans 1120 90 0 0 wbs_dat_o[25]
port 657 nsew signal tristate
flabel metal2 s 106904 -800 107016 480 0 FreeSans 1120 90 0 0 wbs_dat_o[26]
port 658 nsew signal tristate
flabel metal2 s 110450 -800 110562 480 0 FreeSans 1120 90 0 0 wbs_dat_o[27]
port 659 nsew signal tristate
flabel metal2 s 113996 -800 114108 480 0 FreeSans 1120 90 0 0 wbs_dat_o[28]
port 660 nsew signal tristate
flabel metal2 s 117542 -800 117654 480 0 FreeSans 1120 90 0 0 wbs_dat_o[29]
port 661 nsew signal tristate
flabel metal2 s 19436 -800 19548 480 0 FreeSans 1120 90 0 0 wbs_dat_o[2]
port 662 nsew signal tristate
flabel metal2 s 121088 -800 121200 480 0 FreeSans 1120 90 0 0 wbs_dat_o[30]
port 663 nsew signal tristate
flabel metal2 s 124634 -800 124746 480 0 FreeSans 1120 90 0 0 wbs_dat_o[31]
port 664 nsew signal tristate
flabel metal2 s 24164 -800 24276 480 0 FreeSans 1120 90 0 0 wbs_dat_o[3]
port 665 nsew signal tristate
flabel metal2 s 28892 -800 29004 480 0 FreeSans 1120 90 0 0 wbs_dat_o[4]
port 666 nsew signal tristate
flabel metal2 s 32438 -800 32550 480 0 FreeSans 1120 90 0 0 wbs_dat_o[5]
port 667 nsew signal tristate
flabel metal2 s 35984 -800 36096 480 0 FreeSans 1120 90 0 0 wbs_dat_o[6]
port 668 nsew signal tristate
flabel metal2 s 39530 -800 39642 480 0 FreeSans 1120 90 0 0 wbs_dat_o[7]
port 669 nsew signal tristate
flabel metal2 s 43076 -800 43188 480 0 FreeSans 1120 90 0 0 wbs_dat_o[8]
port 670 nsew signal tristate
flabel metal2 s 46622 -800 46734 480 0 FreeSans 1120 90 0 0 wbs_dat_o[9]
port 671 nsew signal tristate
flabel metal2 s 11162 -800 11274 480 0 FreeSans 1120 90 0 0 wbs_sel_i[0]
port 672 nsew signal input
flabel metal2 s 15890 -800 16002 480 0 FreeSans 1120 90 0 0 wbs_sel_i[1]
port 673 nsew signal input
flabel metal2 s 20618 -800 20730 480 0 FreeSans 1120 90 0 0 wbs_sel_i[2]
port 674 nsew signal input
flabel metal2 s 25346 -800 25458 480 0 FreeSans 1120 90 0 0 wbs_sel_i[3]
port 675 nsew signal input
flabel metal2 s 5252 -800 5364 480 0 FreeSans 1120 90 0 0 wbs_stb_i
port 676 nsew signal input
flabel metal2 s 6434 -800 6546 480 0 FreeSans 1120 90 0 0 wbs_we_i
port 677 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
