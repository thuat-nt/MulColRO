magic
tech sky130A
timestamp 1695195202
<< pwell >>
rect -6716 -1248 6716 1248
<< nmoslvt >>
rect -6618 -1143 -6268 1143
rect -6239 -1143 -5889 1143
rect -5860 -1143 -5510 1143
rect -5481 -1143 -5131 1143
rect -5102 -1143 -4752 1143
rect -4723 -1143 -4373 1143
rect -4344 -1143 -3994 1143
rect -3965 -1143 -3615 1143
rect -3586 -1143 -3236 1143
rect -3207 -1143 -2857 1143
rect -2828 -1143 -2478 1143
rect -2449 -1143 -2099 1143
rect -2070 -1143 -1720 1143
rect -1691 -1143 -1341 1143
rect -1312 -1143 -962 1143
rect -933 -1143 -583 1143
rect -554 -1143 -204 1143
rect -175 -1143 175 1143
rect 204 -1143 554 1143
rect 583 -1143 933 1143
rect 962 -1143 1312 1143
rect 1341 -1143 1691 1143
rect 1720 -1143 2070 1143
rect 2099 -1143 2449 1143
rect 2478 -1143 2828 1143
rect 2857 -1143 3207 1143
rect 3236 -1143 3586 1143
rect 3615 -1143 3965 1143
rect 3994 -1143 4344 1143
rect 4373 -1143 4723 1143
rect 4752 -1143 5102 1143
rect 5131 -1143 5481 1143
rect 5510 -1143 5860 1143
rect 5889 -1143 6239 1143
rect 6268 -1143 6618 1143
<< ndiff >>
rect -6647 1137 -6618 1143
rect -6647 -1137 -6641 1137
rect -6624 -1137 -6618 1137
rect -6647 -1143 -6618 -1137
rect -6268 1137 -6239 1143
rect -6268 -1137 -6262 1137
rect -6245 -1137 -6239 1137
rect -6268 -1143 -6239 -1137
rect -5889 1137 -5860 1143
rect -5889 -1137 -5883 1137
rect -5866 -1137 -5860 1137
rect -5889 -1143 -5860 -1137
rect -5510 1137 -5481 1143
rect -5510 -1137 -5504 1137
rect -5487 -1137 -5481 1137
rect -5510 -1143 -5481 -1137
rect -5131 1137 -5102 1143
rect -5131 -1137 -5125 1137
rect -5108 -1137 -5102 1137
rect -5131 -1143 -5102 -1137
rect -4752 1137 -4723 1143
rect -4752 -1137 -4746 1137
rect -4729 -1137 -4723 1137
rect -4752 -1143 -4723 -1137
rect -4373 1137 -4344 1143
rect -4373 -1137 -4367 1137
rect -4350 -1137 -4344 1137
rect -4373 -1143 -4344 -1137
rect -3994 1137 -3965 1143
rect -3994 -1137 -3988 1137
rect -3971 -1137 -3965 1137
rect -3994 -1143 -3965 -1137
rect -3615 1137 -3586 1143
rect -3615 -1137 -3609 1137
rect -3592 -1137 -3586 1137
rect -3615 -1143 -3586 -1137
rect -3236 1137 -3207 1143
rect -3236 -1137 -3230 1137
rect -3213 -1137 -3207 1137
rect -3236 -1143 -3207 -1137
rect -2857 1137 -2828 1143
rect -2857 -1137 -2851 1137
rect -2834 -1137 -2828 1137
rect -2857 -1143 -2828 -1137
rect -2478 1137 -2449 1143
rect -2478 -1137 -2472 1137
rect -2455 -1137 -2449 1137
rect -2478 -1143 -2449 -1137
rect -2099 1137 -2070 1143
rect -2099 -1137 -2093 1137
rect -2076 -1137 -2070 1137
rect -2099 -1143 -2070 -1137
rect -1720 1137 -1691 1143
rect -1720 -1137 -1714 1137
rect -1697 -1137 -1691 1137
rect -1720 -1143 -1691 -1137
rect -1341 1137 -1312 1143
rect -1341 -1137 -1335 1137
rect -1318 -1137 -1312 1137
rect -1341 -1143 -1312 -1137
rect -962 1137 -933 1143
rect -962 -1137 -956 1137
rect -939 -1137 -933 1137
rect -962 -1143 -933 -1137
rect -583 1137 -554 1143
rect -583 -1137 -577 1137
rect -560 -1137 -554 1137
rect -583 -1143 -554 -1137
rect -204 1137 -175 1143
rect -204 -1137 -198 1137
rect -181 -1137 -175 1137
rect -204 -1143 -175 -1137
rect 175 1137 204 1143
rect 175 -1137 181 1137
rect 198 -1137 204 1137
rect 175 -1143 204 -1137
rect 554 1137 583 1143
rect 554 -1137 560 1137
rect 577 -1137 583 1137
rect 554 -1143 583 -1137
rect 933 1137 962 1143
rect 933 -1137 939 1137
rect 956 -1137 962 1137
rect 933 -1143 962 -1137
rect 1312 1137 1341 1143
rect 1312 -1137 1318 1137
rect 1335 -1137 1341 1137
rect 1312 -1143 1341 -1137
rect 1691 1137 1720 1143
rect 1691 -1137 1697 1137
rect 1714 -1137 1720 1137
rect 1691 -1143 1720 -1137
rect 2070 1137 2099 1143
rect 2070 -1137 2076 1137
rect 2093 -1137 2099 1137
rect 2070 -1143 2099 -1137
rect 2449 1137 2478 1143
rect 2449 -1137 2455 1137
rect 2472 -1137 2478 1137
rect 2449 -1143 2478 -1137
rect 2828 1137 2857 1143
rect 2828 -1137 2834 1137
rect 2851 -1137 2857 1137
rect 2828 -1143 2857 -1137
rect 3207 1137 3236 1143
rect 3207 -1137 3213 1137
rect 3230 -1137 3236 1137
rect 3207 -1143 3236 -1137
rect 3586 1137 3615 1143
rect 3586 -1137 3592 1137
rect 3609 -1137 3615 1137
rect 3586 -1143 3615 -1137
rect 3965 1137 3994 1143
rect 3965 -1137 3971 1137
rect 3988 -1137 3994 1137
rect 3965 -1143 3994 -1137
rect 4344 1137 4373 1143
rect 4344 -1137 4350 1137
rect 4367 -1137 4373 1137
rect 4344 -1143 4373 -1137
rect 4723 1137 4752 1143
rect 4723 -1137 4729 1137
rect 4746 -1137 4752 1137
rect 4723 -1143 4752 -1137
rect 5102 1137 5131 1143
rect 5102 -1137 5108 1137
rect 5125 -1137 5131 1137
rect 5102 -1143 5131 -1137
rect 5481 1137 5510 1143
rect 5481 -1137 5487 1137
rect 5504 -1137 5510 1137
rect 5481 -1143 5510 -1137
rect 5860 1137 5889 1143
rect 5860 -1137 5866 1137
rect 5883 -1137 5889 1137
rect 5860 -1143 5889 -1137
rect 6239 1137 6268 1143
rect 6239 -1137 6245 1137
rect 6262 -1137 6268 1137
rect 6239 -1143 6268 -1137
rect 6618 1137 6647 1143
rect 6618 -1137 6624 1137
rect 6641 -1137 6647 1137
rect 6618 -1143 6647 -1137
<< ndiffc >>
rect -6641 -1137 -6624 1137
rect -6262 -1137 -6245 1137
rect -5883 -1137 -5866 1137
rect -5504 -1137 -5487 1137
rect -5125 -1137 -5108 1137
rect -4746 -1137 -4729 1137
rect -4367 -1137 -4350 1137
rect -3988 -1137 -3971 1137
rect -3609 -1137 -3592 1137
rect -3230 -1137 -3213 1137
rect -2851 -1137 -2834 1137
rect -2472 -1137 -2455 1137
rect -2093 -1137 -2076 1137
rect -1714 -1137 -1697 1137
rect -1335 -1137 -1318 1137
rect -956 -1137 -939 1137
rect -577 -1137 -560 1137
rect -198 -1137 -181 1137
rect 181 -1137 198 1137
rect 560 -1137 577 1137
rect 939 -1137 956 1137
rect 1318 -1137 1335 1137
rect 1697 -1137 1714 1137
rect 2076 -1137 2093 1137
rect 2455 -1137 2472 1137
rect 2834 -1137 2851 1137
rect 3213 -1137 3230 1137
rect 3592 -1137 3609 1137
rect 3971 -1137 3988 1137
rect 4350 -1137 4367 1137
rect 4729 -1137 4746 1137
rect 5108 -1137 5125 1137
rect 5487 -1137 5504 1137
rect 5866 -1137 5883 1137
rect 6245 -1137 6262 1137
rect 6624 -1137 6641 1137
<< psubdiff >>
rect -6698 1213 -6650 1230
rect 6650 1213 6698 1230
rect -6698 1182 -6681 1213
rect 6681 1182 6698 1213
rect -6698 -1213 -6681 -1182
rect 6681 -1213 6698 -1182
rect -6698 -1230 -6650 -1213
rect 6650 -1230 6698 -1213
<< psubdiffcont >>
rect -6650 1213 6650 1230
rect -6698 -1182 -6681 1182
rect 6681 -1182 6698 1182
rect -6650 -1230 6650 -1213
<< poly >>
rect -6618 1179 -6268 1187
rect -6618 1162 -6610 1179
rect -6276 1162 -6268 1179
rect -6618 1143 -6268 1162
rect -6239 1179 -5889 1187
rect -6239 1162 -6231 1179
rect -5897 1162 -5889 1179
rect -6239 1143 -5889 1162
rect -5860 1179 -5510 1187
rect -5860 1162 -5852 1179
rect -5518 1162 -5510 1179
rect -5860 1143 -5510 1162
rect -5481 1179 -5131 1187
rect -5481 1162 -5473 1179
rect -5139 1162 -5131 1179
rect -5481 1143 -5131 1162
rect -5102 1179 -4752 1187
rect -5102 1162 -5094 1179
rect -4760 1162 -4752 1179
rect -5102 1143 -4752 1162
rect -4723 1179 -4373 1187
rect -4723 1162 -4715 1179
rect -4381 1162 -4373 1179
rect -4723 1143 -4373 1162
rect -4344 1179 -3994 1187
rect -4344 1162 -4336 1179
rect -4002 1162 -3994 1179
rect -4344 1143 -3994 1162
rect -3965 1179 -3615 1187
rect -3965 1162 -3957 1179
rect -3623 1162 -3615 1179
rect -3965 1143 -3615 1162
rect -3586 1179 -3236 1187
rect -3586 1162 -3578 1179
rect -3244 1162 -3236 1179
rect -3586 1143 -3236 1162
rect -3207 1179 -2857 1187
rect -3207 1162 -3199 1179
rect -2865 1162 -2857 1179
rect -3207 1143 -2857 1162
rect -2828 1179 -2478 1187
rect -2828 1162 -2820 1179
rect -2486 1162 -2478 1179
rect -2828 1143 -2478 1162
rect -2449 1179 -2099 1187
rect -2449 1162 -2441 1179
rect -2107 1162 -2099 1179
rect -2449 1143 -2099 1162
rect -2070 1179 -1720 1187
rect -2070 1162 -2062 1179
rect -1728 1162 -1720 1179
rect -2070 1143 -1720 1162
rect -1691 1179 -1341 1187
rect -1691 1162 -1683 1179
rect -1349 1162 -1341 1179
rect -1691 1143 -1341 1162
rect -1312 1179 -962 1187
rect -1312 1162 -1304 1179
rect -970 1162 -962 1179
rect -1312 1143 -962 1162
rect -933 1179 -583 1187
rect -933 1162 -925 1179
rect -591 1162 -583 1179
rect -933 1143 -583 1162
rect -554 1179 -204 1187
rect -554 1162 -546 1179
rect -212 1162 -204 1179
rect -554 1143 -204 1162
rect -175 1179 175 1187
rect -175 1162 -167 1179
rect 167 1162 175 1179
rect -175 1143 175 1162
rect 204 1179 554 1187
rect 204 1162 212 1179
rect 546 1162 554 1179
rect 204 1143 554 1162
rect 583 1179 933 1187
rect 583 1162 591 1179
rect 925 1162 933 1179
rect 583 1143 933 1162
rect 962 1179 1312 1187
rect 962 1162 970 1179
rect 1304 1162 1312 1179
rect 962 1143 1312 1162
rect 1341 1179 1691 1187
rect 1341 1162 1349 1179
rect 1683 1162 1691 1179
rect 1341 1143 1691 1162
rect 1720 1179 2070 1187
rect 1720 1162 1728 1179
rect 2062 1162 2070 1179
rect 1720 1143 2070 1162
rect 2099 1179 2449 1187
rect 2099 1162 2107 1179
rect 2441 1162 2449 1179
rect 2099 1143 2449 1162
rect 2478 1179 2828 1187
rect 2478 1162 2486 1179
rect 2820 1162 2828 1179
rect 2478 1143 2828 1162
rect 2857 1179 3207 1187
rect 2857 1162 2865 1179
rect 3199 1162 3207 1179
rect 2857 1143 3207 1162
rect 3236 1179 3586 1187
rect 3236 1162 3244 1179
rect 3578 1162 3586 1179
rect 3236 1143 3586 1162
rect 3615 1179 3965 1187
rect 3615 1162 3623 1179
rect 3957 1162 3965 1179
rect 3615 1143 3965 1162
rect 3994 1179 4344 1187
rect 3994 1162 4002 1179
rect 4336 1162 4344 1179
rect 3994 1143 4344 1162
rect 4373 1179 4723 1187
rect 4373 1162 4381 1179
rect 4715 1162 4723 1179
rect 4373 1143 4723 1162
rect 4752 1179 5102 1187
rect 4752 1162 4760 1179
rect 5094 1162 5102 1179
rect 4752 1143 5102 1162
rect 5131 1179 5481 1187
rect 5131 1162 5139 1179
rect 5473 1162 5481 1179
rect 5131 1143 5481 1162
rect 5510 1179 5860 1187
rect 5510 1162 5518 1179
rect 5852 1162 5860 1179
rect 5510 1143 5860 1162
rect 5889 1179 6239 1187
rect 5889 1162 5897 1179
rect 6231 1162 6239 1179
rect 5889 1143 6239 1162
rect 6268 1179 6618 1187
rect 6268 1162 6276 1179
rect 6610 1162 6618 1179
rect 6268 1143 6618 1162
rect -6618 -1162 -6268 -1143
rect -6618 -1179 -6610 -1162
rect -6276 -1179 -6268 -1162
rect -6618 -1187 -6268 -1179
rect -6239 -1162 -5889 -1143
rect -6239 -1179 -6231 -1162
rect -5897 -1179 -5889 -1162
rect -6239 -1187 -5889 -1179
rect -5860 -1162 -5510 -1143
rect -5860 -1179 -5852 -1162
rect -5518 -1179 -5510 -1162
rect -5860 -1187 -5510 -1179
rect -5481 -1162 -5131 -1143
rect -5481 -1179 -5473 -1162
rect -5139 -1179 -5131 -1162
rect -5481 -1187 -5131 -1179
rect -5102 -1162 -4752 -1143
rect -5102 -1179 -5094 -1162
rect -4760 -1179 -4752 -1162
rect -5102 -1187 -4752 -1179
rect -4723 -1162 -4373 -1143
rect -4723 -1179 -4715 -1162
rect -4381 -1179 -4373 -1162
rect -4723 -1187 -4373 -1179
rect -4344 -1162 -3994 -1143
rect -4344 -1179 -4336 -1162
rect -4002 -1179 -3994 -1162
rect -4344 -1187 -3994 -1179
rect -3965 -1162 -3615 -1143
rect -3965 -1179 -3957 -1162
rect -3623 -1179 -3615 -1162
rect -3965 -1187 -3615 -1179
rect -3586 -1162 -3236 -1143
rect -3586 -1179 -3578 -1162
rect -3244 -1179 -3236 -1162
rect -3586 -1187 -3236 -1179
rect -3207 -1162 -2857 -1143
rect -3207 -1179 -3199 -1162
rect -2865 -1179 -2857 -1162
rect -3207 -1187 -2857 -1179
rect -2828 -1162 -2478 -1143
rect -2828 -1179 -2820 -1162
rect -2486 -1179 -2478 -1162
rect -2828 -1187 -2478 -1179
rect -2449 -1162 -2099 -1143
rect -2449 -1179 -2441 -1162
rect -2107 -1179 -2099 -1162
rect -2449 -1187 -2099 -1179
rect -2070 -1162 -1720 -1143
rect -2070 -1179 -2062 -1162
rect -1728 -1179 -1720 -1162
rect -2070 -1187 -1720 -1179
rect -1691 -1162 -1341 -1143
rect -1691 -1179 -1683 -1162
rect -1349 -1179 -1341 -1162
rect -1691 -1187 -1341 -1179
rect -1312 -1162 -962 -1143
rect -1312 -1179 -1304 -1162
rect -970 -1179 -962 -1162
rect -1312 -1187 -962 -1179
rect -933 -1162 -583 -1143
rect -933 -1179 -925 -1162
rect -591 -1179 -583 -1162
rect -933 -1187 -583 -1179
rect -554 -1162 -204 -1143
rect -554 -1179 -546 -1162
rect -212 -1179 -204 -1162
rect -554 -1187 -204 -1179
rect -175 -1162 175 -1143
rect -175 -1179 -167 -1162
rect 167 -1179 175 -1162
rect -175 -1187 175 -1179
rect 204 -1162 554 -1143
rect 204 -1179 212 -1162
rect 546 -1179 554 -1162
rect 204 -1187 554 -1179
rect 583 -1162 933 -1143
rect 583 -1179 591 -1162
rect 925 -1179 933 -1162
rect 583 -1187 933 -1179
rect 962 -1162 1312 -1143
rect 962 -1179 970 -1162
rect 1304 -1179 1312 -1162
rect 962 -1187 1312 -1179
rect 1341 -1162 1691 -1143
rect 1341 -1179 1349 -1162
rect 1683 -1179 1691 -1162
rect 1341 -1187 1691 -1179
rect 1720 -1162 2070 -1143
rect 1720 -1179 1728 -1162
rect 2062 -1179 2070 -1162
rect 1720 -1187 2070 -1179
rect 2099 -1162 2449 -1143
rect 2099 -1179 2107 -1162
rect 2441 -1179 2449 -1162
rect 2099 -1187 2449 -1179
rect 2478 -1162 2828 -1143
rect 2478 -1179 2486 -1162
rect 2820 -1179 2828 -1162
rect 2478 -1187 2828 -1179
rect 2857 -1162 3207 -1143
rect 2857 -1179 2865 -1162
rect 3199 -1179 3207 -1162
rect 2857 -1187 3207 -1179
rect 3236 -1162 3586 -1143
rect 3236 -1179 3244 -1162
rect 3578 -1179 3586 -1162
rect 3236 -1187 3586 -1179
rect 3615 -1162 3965 -1143
rect 3615 -1179 3623 -1162
rect 3957 -1179 3965 -1162
rect 3615 -1187 3965 -1179
rect 3994 -1162 4344 -1143
rect 3994 -1179 4002 -1162
rect 4336 -1179 4344 -1162
rect 3994 -1187 4344 -1179
rect 4373 -1162 4723 -1143
rect 4373 -1179 4381 -1162
rect 4715 -1179 4723 -1162
rect 4373 -1187 4723 -1179
rect 4752 -1162 5102 -1143
rect 4752 -1179 4760 -1162
rect 5094 -1179 5102 -1162
rect 4752 -1187 5102 -1179
rect 5131 -1162 5481 -1143
rect 5131 -1179 5139 -1162
rect 5473 -1179 5481 -1162
rect 5131 -1187 5481 -1179
rect 5510 -1162 5860 -1143
rect 5510 -1179 5518 -1162
rect 5852 -1179 5860 -1162
rect 5510 -1187 5860 -1179
rect 5889 -1162 6239 -1143
rect 5889 -1179 5897 -1162
rect 6231 -1179 6239 -1162
rect 5889 -1187 6239 -1179
rect 6268 -1162 6618 -1143
rect 6268 -1179 6276 -1162
rect 6610 -1179 6618 -1162
rect 6268 -1187 6618 -1179
<< polycont >>
rect -6610 1162 -6276 1179
rect -6231 1162 -5897 1179
rect -5852 1162 -5518 1179
rect -5473 1162 -5139 1179
rect -5094 1162 -4760 1179
rect -4715 1162 -4381 1179
rect -4336 1162 -4002 1179
rect -3957 1162 -3623 1179
rect -3578 1162 -3244 1179
rect -3199 1162 -2865 1179
rect -2820 1162 -2486 1179
rect -2441 1162 -2107 1179
rect -2062 1162 -1728 1179
rect -1683 1162 -1349 1179
rect -1304 1162 -970 1179
rect -925 1162 -591 1179
rect -546 1162 -212 1179
rect -167 1162 167 1179
rect 212 1162 546 1179
rect 591 1162 925 1179
rect 970 1162 1304 1179
rect 1349 1162 1683 1179
rect 1728 1162 2062 1179
rect 2107 1162 2441 1179
rect 2486 1162 2820 1179
rect 2865 1162 3199 1179
rect 3244 1162 3578 1179
rect 3623 1162 3957 1179
rect 4002 1162 4336 1179
rect 4381 1162 4715 1179
rect 4760 1162 5094 1179
rect 5139 1162 5473 1179
rect 5518 1162 5852 1179
rect 5897 1162 6231 1179
rect 6276 1162 6610 1179
rect -6610 -1179 -6276 -1162
rect -6231 -1179 -5897 -1162
rect -5852 -1179 -5518 -1162
rect -5473 -1179 -5139 -1162
rect -5094 -1179 -4760 -1162
rect -4715 -1179 -4381 -1162
rect -4336 -1179 -4002 -1162
rect -3957 -1179 -3623 -1162
rect -3578 -1179 -3244 -1162
rect -3199 -1179 -2865 -1162
rect -2820 -1179 -2486 -1162
rect -2441 -1179 -2107 -1162
rect -2062 -1179 -1728 -1162
rect -1683 -1179 -1349 -1162
rect -1304 -1179 -970 -1162
rect -925 -1179 -591 -1162
rect -546 -1179 -212 -1162
rect -167 -1179 167 -1162
rect 212 -1179 546 -1162
rect 591 -1179 925 -1162
rect 970 -1179 1304 -1162
rect 1349 -1179 1683 -1162
rect 1728 -1179 2062 -1162
rect 2107 -1179 2441 -1162
rect 2486 -1179 2820 -1162
rect 2865 -1179 3199 -1162
rect 3244 -1179 3578 -1162
rect 3623 -1179 3957 -1162
rect 4002 -1179 4336 -1162
rect 4381 -1179 4715 -1162
rect 4760 -1179 5094 -1162
rect 5139 -1179 5473 -1162
rect 5518 -1179 5852 -1162
rect 5897 -1179 6231 -1162
rect 6276 -1179 6610 -1162
<< locali >>
rect -6698 1213 -6650 1230
rect 6650 1213 6698 1230
rect -6698 1182 -6681 1213
rect 6681 1182 6698 1213
rect -6618 1162 -6610 1179
rect -6276 1162 -6268 1179
rect -6239 1162 -6231 1179
rect -5897 1162 -5889 1179
rect -5860 1162 -5852 1179
rect -5518 1162 -5510 1179
rect -5481 1162 -5473 1179
rect -5139 1162 -5131 1179
rect -5102 1162 -5094 1179
rect -4760 1162 -4752 1179
rect -4723 1162 -4715 1179
rect -4381 1162 -4373 1179
rect -4344 1162 -4336 1179
rect -4002 1162 -3994 1179
rect -3965 1162 -3957 1179
rect -3623 1162 -3615 1179
rect -3586 1162 -3578 1179
rect -3244 1162 -3236 1179
rect -3207 1162 -3199 1179
rect -2865 1162 -2857 1179
rect -2828 1162 -2820 1179
rect -2486 1162 -2478 1179
rect -2449 1162 -2441 1179
rect -2107 1162 -2099 1179
rect -2070 1162 -2062 1179
rect -1728 1162 -1720 1179
rect -1691 1162 -1683 1179
rect -1349 1162 -1341 1179
rect -1312 1162 -1304 1179
rect -970 1162 -962 1179
rect -933 1162 -925 1179
rect -591 1162 -583 1179
rect -554 1162 -546 1179
rect -212 1162 -204 1179
rect -175 1162 -167 1179
rect 167 1162 175 1179
rect 204 1162 212 1179
rect 546 1162 554 1179
rect 583 1162 591 1179
rect 925 1162 933 1179
rect 962 1162 970 1179
rect 1304 1162 1312 1179
rect 1341 1162 1349 1179
rect 1683 1162 1691 1179
rect 1720 1162 1728 1179
rect 2062 1162 2070 1179
rect 2099 1162 2107 1179
rect 2441 1162 2449 1179
rect 2478 1162 2486 1179
rect 2820 1162 2828 1179
rect 2857 1162 2865 1179
rect 3199 1162 3207 1179
rect 3236 1162 3244 1179
rect 3578 1162 3586 1179
rect 3615 1162 3623 1179
rect 3957 1162 3965 1179
rect 3994 1162 4002 1179
rect 4336 1162 4344 1179
rect 4373 1162 4381 1179
rect 4715 1162 4723 1179
rect 4752 1162 4760 1179
rect 5094 1162 5102 1179
rect 5131 1162 5139 1179
rect 5473 1162 5481 1179
rect 5510 1162 5518 1179
rect 5852 1162 5860 1179
rect 5889 1162 5897 1179
rect 6231 1162 6239 1179
rect 6268 1162 6276 1179
rect 6610 1162 6618 1179
rect -6641 1137 -6624 1145
rect -6641 -1145 -6624 -1137
rect -6262 1137 -6245 1145
rect -6262 -1145 -6245 -1137
rect -5883 1137 -5866 1145
rect -5883 -1145 -5866 -1137
rect -5504 1137 -5487 1145
rect -5504 -1145 -5487 -1137
rect -5125 1137 -5108 1145
rect -5125 -1145 -5108 -1137
rect -4746 1137 -4729 1145
rect -4746 -1145 -4729 -1137
rect -4367 1137 -4350 1145
rect -4367 -1145 -4350 -1137
rect -3988 1137 -3971 1145
rect -3988 -1145 -3971 -1137
rect -3609 1137 -3592 1145
rect -3609 -1145 -3592 -1137
rect -3230 1137 -3213 1145
rect -3230 -1145 -3213 -1137
rect -2851 1137 -2834 1145
rect -2851 -1145 -2834 -1137
rect -2472 1137 -2455 1145
rect -2472 -1145 -2455 -1137
rect -2093 1137 -2076 1145
rect -2093 -1145 -2076 -1137
rect -1714 1137 -1697 1145
rect -1714 -1145 -1697 -1137
rect -1335 1137 -1318 1145
rect -1335 -1145 -1318 -1137
rect -956 1137 -939 1145
rect -956 -1145 -939 -1137
rect -577 1137 -560 1145
rect -577 -1145 -560 -1137
rect -198 1137 -181 1145
rect -198 -1145 -181 -1137
rect 181 1137 198 1145
rect 181 -1145 198 -1137
rect 560 1137 577 1145
rect 560 -1145 577 -1137
rect 939 1137 956 1145
rect 939 -1145 956 -1137
rect 1318 1137 1335 1145
rect 1318 -1145 1335 -1137
rect 1697 1137 1714 1145
rect 1697 -1145 1714 -1137
rect 2076 1137 2093 1145
rect 2076 -1145 2093 -1137
rect 2455 1137 2472 1145
rect 2455 -1145 2472 -1137
rect 2834 1137 2851 1145
rect 2834 -1145 2851 -1137
rect 3213 1137 3230 1145
rect 3213 -1145 3230 -1137
rect 3592 1137 3609 1145
rect 3592 -1145 3609 -1137
rect 3971 1137 3988 1145
rect 3971 -1145 3988 -1137
rect 4350 1137 4367 1145
rect 4350 -1145 4367 -1137
rect 4729 1137 4746 1145
rect 4729 -1145 4746 -1137
rect 5108 1137 5125 1145
rect 5108 -1145 5125 -1137
rect 5487 1137 5504 1145
rect 5487 -1145 5504 -1137
rect 5866 1137 5883 1145
rect 5866 -1145 5883 -1137
rect 6245 1137 6262 1145
rect 6245 -1145 6262 -1137
rect 6624 1137 6641 1145
rect 6624 -1145 6641 -1137
rect -6618 -1179 -6610 -1162
rect -6276 -1179 -6268 -1162
rect -6239 -1179 -6231 -1162
rect -5897 -1179 -5889 -1162
rect -5860 -1179 -5852 -1162
rect -5518 -1179 -5510 -1162
rect -5481 -1179 -5473 -1162
rect -5139 -1179 -5131 -1162
rect -5102 -1179 -5094 -1162
rect -4760 -1179 -4752 -1162
rect -4723 -1179 -4715 -1162
rect -4381 -1179 -4373 -1162
rect -4344 -1179 -4336 -1162
rect -4002 -1179 -3994 -1162
rect -3965 -1179 -3957 -1162
rect -3623 -1179 -3615 -1162
rect -3586 -1179 -3578 -1162
rect -3244 -1179 -3236 -1162
rect -3207 -1179 -3199 -1162
rect -2865 -1179 -2857 -1162
rect -2828 -1179 -2820 -1162
rect -2486 -1179 -2478 -1162
rect -2449 -1179 -2441 -1162
rect -2107 -1179 -2099 -1162
rect -2070 -1179 -2062 -1162
rect -1728 -1179 -1720 -1162
rect -1691 -1179 -1683 -1162
rect -1349 -1179 -1341 -1162
rect -1312 -1179 -1304 -1162
rect -970 -1179 -962 -1162
rect -933 -1179 -925 -1162
rect -591 -1179 -583 -1162
rect -554 -1179 -546 -1162
rect -212 -1179 -204 -1162
rect -175 -1179 -167 -1162
rect 167 -1179 175 -1162
rect 204 -1179 212 -1162
rect 546 -1179 554 -1162
rect 583 -1179 591 -1162
rect 925 -1179 933 -1162
rect 962 -1179 970 -1162
rect 1304 -1179 1312 -1162
rect 1341 -1179 1349 -1162
rect 1683 -1179 1691 -1162
rect 1720 -1179 1728 -1162
rect 2062 -1179 2070 -1162
rect 2099 -1179 2107 -1162
rect 2441 -1179 2449 -1162
rect 2478 -1179 2486 -1162
rect 2820 -1179 2828 -1162
rect 2857 -1179 2865 -1162
rect 3199 -1179 3207 -1162
rect 3236 -1179 3244 -1162
rect 3578 -1179 3586 -1162
rect 3615 -1179 3623 -1162
rect 3957 -1179 3965 -1162
rect 3994 -1179 4002 -1162
rect 4336 -1179 4344 -1162
rect 4373 -1179 4381 -1162
rect 4715 -1179 4723 -1162
rect 4752 -1179 4760 -1162
rect 5094 -1179 5102 -1162
rect 5131 -1179 5139 -1162
rect 5473 -1179 5481 -1162
rect 5510 -1179 5518 -1162
rect 5852 -1179 5860 -1162
rect 5889 -1179 5897 -1162
rect 6231 -1179 6239 -1162
rect 6268 -1179 6276 -1162
rect 6610 -1179 6618 -1162
rect -6698 -1213 -6681 -1182
rect 6681 -1213 6698 -1182
rect -6698 -1230 -6650 -1213
rect 6650 -1230 6698 -1213
<< viali >>
rect -6610 1162 -6276 1179
rect -6231 1162 -5897 1179
rect -5852 1162 -5518 1179
rect -5473 1162 -5139 1179
rect -5094 1162 -4760 1179
rect -4715 1162 -4381 1179
rect -4336 1162 -4002 1179
rect -3957 1162 -3623 1179
rect -3578 1162 -3244 1179
rect -3199 1162 -2865 1179
rect -2820 1162 -2486 1179
rect -2441 1162 -2107 1179
rect -2062 1162 -1728 1179
rect -1683 1162 -1349 1179
rect -1304 1162 -970 1179
rect -925 1162 -591 1179
rect -546 1162 -212 1179
rect -167 1162 167 1179
rect 212 1162 546 1179
rect 591 1162 925 1179
rect 970 1162 1304 1179
rect 1349 1162 1683 1179
rect 1728 1162 2062 1179
rect 2107 1162 2441 1179
rect 2486 1162 2820 1179
rect 2865 1162 3199 1179
rect 3244 1162 3578 1179
rect 3623 1162 3957 1179
rect 4002 1162 4336 1179
rect 4381 1162 4715 1179
rect 4760 1162 5094 1179
rect 5139 1162 5473 1179
rect 5518 1162 5852 1179
rect 5897 1162 6231 1179
rect 6276 1162 6610 1179
rect -6641 -1137 -6624 1137
rect -6262 -1137 -6245 1137
rect -5883 -1137 -5866 1137
rect -5504 -1137 -5487 1137
rect -5125 -1137 -5108 1137
rect -4746 -1137 -4729 1137
rect -4367 -1137 -4350 1137
rect -3988 -1137 -3971 1137
rect -3609 -1137 -3592 1137
rect -3230 -1137 -3213 1137
rect -2851 -1137 -2834 1137
rect -2472 -1137 -2455 1137
rect -2093 -1137 -2076 1137
rect -1714 -1137 -1697 1137
rect -1335 -1137 -1318 1137
rect -956 -1137 -939 1137
rect -577 -1137 -560 1137
rect -198 -1137 -181 1137
rect 181 -1137 198 1137
rect 560 -1137 577 1137
rect 939 -1137 956 1137
rect 1318 -1137 1335 1137
rect 1697 -1137 1714 1137
rect 2076 -1137 2093 1137
rect 2455 -1137 2472 1137
rect 2834 -1137 2851 1137
rect 3213 -1137 3230 1137
rect 3592 -1137 3609 1137
rect 3971 -1137 3988 1137
rect 4350 -1137 4367 1137
rect 4729 -1137 4746 1137
rect 5108 -1137 5125 1137
rect 5487 -1137 5504 1137
rect 5866 -1137 5883 1137
rect 6245 -1137 6262 1137
rect 6624 -1137 6641 1137
rect -6610 -1179 -6276 -1162
rect -6231 -1179 -5897 -1162
rect -5852 -1179 -5518 -1162
rect -5473 -1179 -5139 -1162
rect -5094 -1179 -4760 -1162
rect -4715 -1179 -4381 -1162
rect -4336 -1179 -4002 -1162
rect -3957 -1179 -3623 -1162
rect -3578 -1179 -3244 -1162
rect -3199 -1179 -2865 -1162
rect -2820 -1179 -2486 -1162
rect -2441 -1179 -2107 -1162
rect -2062 -1179 -1728 -1162
rect -1683 -1179 -1349 -1162
rect -1304 -1179 -970 -1162
rect -925 -1179 -591 -1162
rect -546 -1179 -212 -1162
rect -167 -1179 167 -1162
rect 212 -1179 546 -1162
rect 591 -1179 925 -1162
rect 970 -1179 1304 -1162
rect 1349 -1179 1683 -1162
rect 1728 -1179 2062 -1162
rect 2107 -1179 2441 -1162
rect 2486 -1179 2820 -1162
rect 2865 -1179 3199 -1162
rect 3244 -1179 3578 -1162
rect 3623 -1179 3957 -1162
rect 4002 -1179 4336 -1162
rect 4381 -1179 4715 -1162
rect 4760 -1179 5094 -1162
rect 5139 -1179 5473 -1162
rect 5518 -1179 5852 -1162
rect 5897 -1179 6231 -1162
rect 6276 -1179 6610 -1162
<< metal1 >>
rect -6616 1179 -6270 1182
rect -6616 1162 -6610 1179
rect -6276 1162 -6270 1179
rect -6616 1159 -6270 1162
rect -6237 1179 -5891 1182
rect -6237 1162 -6231 1179
rect -5897 1162 -5891 1179
rect -6237 1159 -5891 1162
rect -5858 1179 -5512 1182
rect -5858 1162 -5852 1179
rect -5518 1162 -5512 1179
rect -5858 1159 -5512 1162
rect -5479 1179 -5133 1182
rect -5479 1162 -5473 1179
rect -5139 1162 -5133 1179
rect -5479 1159 -5133 1162
rect -5100 1179 -4754 1182
rect -5100 1162 -5094 1179
rect -4760 1162 -4754 1179
rect -5100 1159 -4754 1162
rect -4721 1179 -4375 1182
rect -4721 1162 -4715 1179
rect -4381 1162 -4375 1179
rect -4721 1159 -4375 1162
rect -4342 1179 -3996 1182
rect -4342 1162 -4336 1179
rect -4002 1162 -3996 1179
rect -4342 1159 -3996 1162
rect -3963 1179 -3617 1182
rect -3963 1162 -3957 1179
rect -3623 1162 -3617 1179
rect -3963 1159 -3617 1162
rect -3584 1179 -3238 1182
rect -3584 1162 -3578 1179
rect -3244 1162 -3238 1179
rect -3584 1159 -3238 1162
rect -3205 1179 -2859 1182
rect -3205 1162 -3199 1179
rect -2865 1162 -2859 1179
rect -3205 1159 -2859 1162
rect -2826 1179 -2480 1182
rect -2826 1162 -2820 1179
rect -2486 1162 -2480 1179
rect -2826 1159 -2480 1162
rect -2447 1179 -2101 1182
rect -2447 1162 -2441 1179
rect -2107 1162 -2101 1179
rect -2447 1159 -2101 1162
rect -2068 1179 -1722 1182
rect -2068 1162 -2062 1179
rect -1728 1162 -1722 1179
rect -2068 1159 -1722 1162
rect -1689 1179 -1343 1182
rect -1689 1162 -1683 1179
rect -1349 1162 -1343 1179
rect -1689 1159 -1343 1162
rect -1310 1179 -964 1182
rect -1310 1162 -1304 1179
rect -970 1162 -964 1179
rect -1310 1159 -964 1162
rect -931 1179 -585 1182
rect -931 1162 -925 1179
rect -591 1162 -585 1179
rect -931 1159 -585 1162
rect -552 1179 -206 1182
rect -552 1162 -546 1179
rect -212 1162 -206 1179
rect -552 1159 -206 1162
rect -173 1179 173 1182
rect -173 1162 -167 1179
rect 167 1162 173 1179
rect -173 1159 173 1162
rect 206 1179 552 1182
rect 206 1162 212 1179
rect 546 1162 552 1179
rect 206 1159 552 1162
rect 585 1179 931 1182
rect 585 1162 591 1179
rect 925 1162 931 1179
rect 585 1159 931 1162
rect 964 1179 1310 1182
rect 964 1162 970 1179
rect 1304 1162 1310 1179
rect 964 1159 1310 1162
rect 1343 1179 1689 1182
rect 1343 1162 1349 1179
rect 1683 1162 1689 1179
rect 1343 1159 1689 1162
rect 1722 1179 2068 1182
rect 1722 1162 1728 1179
rect 2062 1162 2068 1179
rect 1722 1159 2068 1162
rect 2101 1179 2447 1182
rect 2101 1162 2107 1179
rect 2441 1162 2447 1179
rect 2101 1159 2447 1162
rect 2480 1179 2826 1182
rect 2480 1162 2486 1179
rect 2820 1162 2826 1179
rect 2480 1159 2826 1162
rect 2859 1179 3205 1182
rect 2859 1162 2865 1179
rect 3199 1162 3205 1179
rect 2859 1159 3205 1162
rect 3238 1179 3584 1182
rect 3238 1162 3244 1179
rect 3578 1162 3584 1179
rect 3238 1159 3584 1162
rect 3617 1179 3963 1182
rect 3617 1162 3623 1179
rect 3957 1162 3963 1179
rect 3617 1159 3963 1162
rect 3996 1179 4342 1182
rect 3996 1162 4002 1179
rect 4336 1162 4342 1179
rect 3996 1159 4342 1162
rect 4375 1179 4721 1182
rect 4375 1162 4381 1179
rect 4715 1162 4721 1179
rect 4375 1159 4721 1162
rect 4754 1179 5100 1182
rect 4754 1162 4760 1179
rect 5094 1162 5100 1179
rect 4754 1159 5100 1162
rect 5133 1179 5479 1182
rect 5133 1162 5139 1179
rect 5473 1162 5479 1179
rect 5133 1159 5479 1162
rect 5512 1179 5858 1182
rect 5512 1162 5518 1179
rect 5852 1162 5858 1179
rect 5512 1159 5858 1162
rect 5891 1179 6237 1182
rect 5891 1162 5897 1179
rect 6231 1162 6237 1179
rect 5891 1159 6237 1162
rect 6270 1179 6616 1182
rect 6270 1162 6276 1179
rect 6610 1162 6616 1179
rect 6270 1159 6616 1162
rect -6644 1137 -6621 1143
rect -6644 -1137 -6641 1137
rect -6624 -1137 -6621 1137
rect -6644 -1143 -6621 -1137
rect -6265 1137 -6242 1143
rect -6265 -1137 -6262 1137
rect -6245 -1137 -6242 1137
rect -6265 -1143 -6242 -1137
rect -5886 1137 -5863 1143
rect -5886 -1137 -5883 1137
rect -5866 -1137 -5863 1137
rect -5886 -1143 -5863 -1137
rect -5507 1137 -5484 1143
rect -5507 -1137 -5504 1137
rect -5487 -1137 -5484 1137
rect -5507 -1143 -5484 -1137
rect -5128 1137 -5105 1143
rect -5128 -1137 -5125 1137
rect -5108 -1137 -5105 1137
rect -5128 -1143 -5105 -1137
rect -4749 1137 -4726 1143
rect -4749 -1137 -4746 1137
rect -4729 -1137 -4726 1137
rect -4749 -1143 -4726 -1137
rect -4370 1137 -4347 1143
rect -4370 -1137 -4367 1137
rect -4350 -1137 -4347 1137
rect -4370 -1143 -4347 -1137
rect -3991 1137 -3968 1143
rect -3991 -1137 -3988 1137
rect -3971 -1137 -3968 1137
rect -3991 -1143 -3968 -1137
rect -3612 1137 -3589 1143
rect -3612 -1137 -3609 1137
rect -3592 -1137 -3589 1137
rect -3612 -1143 -3589 -1137
rect -3233 1137 -3210 1143
rect -3233 -1137 -3230 1137
rect -3213 -1137 -3210 1137
rect -3233 -1143 -3210 -1137
rect -2854 1137 -2831 1143
rect -2854 -1137 -2851 1137
rect -2834 -1137 -2831 1137
rect -2854 -1143 -2831 -1137
rect -2475 1137 -2452 1143
rect -2475 -1137 -2472 1137
rect -2455 -1137 -2452 1137
rect -2475 -1143 -2452 -1137
rect -2096 1137 -2073 1143
rect -2096 -1137 -2093 1137
rect -2076 -1137 -2073 1137
rect -2096 -1143 -2073 -1137
rect -1717 1137 -1694 1143
rect -1717 -1137 -1714 1137
rect -1697 -1137 -1694 1137
rect -1717 -1143 -1694 -1137
rect -1338 1137 -1315 1143
rect -1338 -1137 -1335 1137
rect -1318 -1137 -1315 1137
rect -1338 -1143 -1315 -1137
rect -959 1137 -936 1143
rect -959 -1137 -956 1137
rect -939 -1137 -936 1137
rect -959 -1143 -936 -1137
rect -580 1137 -557 1143
rect -580 -1137 -577 1137
rect -560 -1137 -557 1137
rect -580 -1143 -557 -1137
rect -201 1137 -178 1143
rect -201 -1137 -198 1137
rect -181 -1137 -178 1137
rect -201 -1143 -178 -1137
rect 178 1137 201 1143
rect 178 -1137 181 1137
rect 198 -1137 201 1137
rect 178 -1143 201 -1137
rect 557 1137 580 1143
rect 557 -1137 560 1137
rect 577 -1137 580 1137
rect 557 -1143 580 -1137
rect 936 1137 959 1143
rect 936 -1137 939 1137
rect 956 -1137 959 1137
rect 936 -1143 959 -1137
rect 1315 1137 1338 1143
rect 1315 -1137 1318 1137
rect 1335 -1137 1338 1137
rect 1315 -1143 1338 -1137
rect 1694 1137 1717 1143
rect 1694 -1137 1697 1137
rect 1714 -1137 1717 1137
rect 1694 -1143 1717 -1137
rect 2073 1137 2096 1143
rect 2073 -1137 2076 1137
rect 2093 -1137 2096 1137
rect 2073 -1143 2096 -1137
rect 2452 1137 2475 1143
rect 2452 -1137 2455 1137
rect 2472 -1137 2475 1137
rect 2452 -1143 2475 -1137
rect 2831 1137 2854 1143
rect 2831 -1137 2834 1137
rect 2851 -1137 2854 1137
rect 2831 -1143 2854 -1137
rect 3210 1137 3233 1143
rect 3210 -1137 3213 1137
rect 3230 -1137 3233 1137
rect 3210 -1143 3233 -1137
rect 3589 1137 3612 1143
rect 3589 -1137 3592 1137
rect 3609 -1137 3612 1137
rect 3589 -1143 3612 -1137
rect 3968 1137 3991 1143
rect 3968 -1137 3971 1137
rect 3988 -1137 3991 1137
rect 3968 -1143 3991 -1137
rect 4347 1137 4370 1143
rect 4347 -1137 4350 1137
rect 4367 -1137 4370 1137
rect 4347 -1143 4370 -1137
rect 4726 1137 4749 1143
rect 4726 -1137 4729 1137
rect 4746 -1137 4749 1137
rect 4726 -1143 4749 -1137
rect 5105 1137 5128 1143
rect 5105 -1137 5108 1137
rect 5125 -1137 5128 1137
rect 5105 -1143 5128 -1137
rect 5484 1137 5507 1143
rect 5484 -1137 5487 1137
rect 5504 -1137 5507 1137
rect 5484 -1143 5507 -1137
rect 5863 1137 5886 1143
rect 5863 -1137 5866 1137
rect 5883 -1137 5886 1137
rect 5863 -1143 5886 -1137
rect 6242 1137 6265 1143
rect 6242 -1137 6245 1137
rect 6262 -1137 6265 1137
rect 6242 -1143 6265 -1137
rect 6621 1137 6644 1143
rect 6621 -1137 6624 1137
rect 6641 -1137 6644 1137
rect 6621 -1143 6644 -1137
rect -6616 -1162 -6270 -1159
rect -6616 -1179 -6610 -1162
rect -6276 -1179 -6270 -1162
rect -6616 -1182 -6270 -1179
rect -6237 -1162 -5891 -1159
rect -6237 -1179 -6231 -1162
rect -5897 -1179 -5891 -1162
rect -6237 -1182 -5891 -1179
rect -5858 -1162 -5512 -1159
rect -5858 -1179 -5852 -1162
rect -5518 -1179 -5512 -1162
rect -5858 -1182 -5512 -1179
rect -5479 -1162 -5133 -1159
rect -5479 -1179 -5473 -1162
rect -5139 -1179 -5133 -1162
rect -5479 -1182 -5133 -1179
rect -5100 -1162 -4754 -1159
rect -5100 -1179 -5094 -1162
rect -4760 -1179 -4754 -1162
rect -5100 -1182 -4754 -1179
rect -4721 -1162 -4375 -1159
rect -4721 -1179 -4715 -1162
rect -4381 -1179 -4375 -1162
rect -4721 -1182 -4375 -1179
rect -4342 -1162 -3996 -1159
rect -4342 -1179 -4336 -1162
rect -4002 -1179 -3996 -1162
rect -4342 -1182 -3996 -1179
rect -3963 -1162 -3617 -1159
rect -3963 -1179 -3957 -1162
rect -3623 -1179 -3617 -1162
rect -3963 -1182 -3617 -1179
rect -3584 -1162 -3238 -1159
rect -3584 -1179 -3578 -1162
rect -3244 -1179 -3238 -1162
rect -3584 -1182 -3238 -1179
rect -3205 -1162 -2859 -1159
rect -3205 -1179 -3199 -1162
rect -2865 -1179 -2859 -1162
rect -3205 -1182 -2859 -1179
rect -2826 -1162 -2480 -1159
rect -2826 -1179 -2820 -1162
rect -2486 -1179 -2480 -1162
rect -2826 -1182 -2480 -1179
rect -2447 -1162 -2101 -1159
rect -2447 -1179 -2441 -1162
rect -2107 -1179 -2101 -1162
rect -2447 -1182 -2101 -1179
rect -2068 -1162 -1722 -1159
rect -2068 -1179 -2062 -1162
rect -1728 -1179 -1722 -1162
rect -2068 -1182 -1722 -1179
rect -1689 -1162 -1343 -1159
rect -1689 -1179 -1683 -1162
rect -1349 -1179 -1343 -1162
rect -1689 -1182 -1343 -1179
rect -1310 -1162 -964 -1159
rect -1310 -1179 -1304 -1162
rect -970 -1179 -964 -1162
rect -1310 -1182 -964 -1179
rect -931 -1162 -585 -1159
rect -931 -1179 -925 -1162
rect -591 -1179 -585 -1162
rect -931 -1182 -585 -1179
rect -552 -1162 -206 -1159
rect -552 -1179 -546 -1162
rect -212 -1179 -206 -1162
rect -552 -1182 -206 -1179
rect -173 -1162 173 -1159
rect -173 -1179 -167 -1162
rect 167 -1179 173 -1162
rect -173 -1182 173 -1179
rect 206 -1162 552 -1159
rect 206 -1179 212 -1162
rect 546 -1179 552 -1162
rect 206 -1182 552 -1179
rect 585 -1162 931 -1159
rect 585 -1179 591 -1162
rect 925 -1179 931 -1162
rect 585 -1182 931 -1179
rect 964 -1162 1310 -1159
rect 964 -1179 970 -1162
rect 1304 -1179 1310 -1162
rect 964 -1182 1310 -1179
rect 1343 -1162 1689 -1159
rect 1343 -1179 1349 -1162
rect 1683 -1179 1689 -1162
rect 1343 -1182 1689 -1179
rect 1722 -1162 2068 -1159
rect 1722 -1179 1728 -1162
rect 2062 -1179 2068 -1162
rect 1722 -1182 2068 -1179
rect 2101 -1162 2447 -1159
rect 2101 -1179 2107 -1162
rect 2441 -1179 2447 -1162
rect 2101 -1182 2447 -1179
rect 2480 -1162 2826 -1159
rect 2480 -1179 2486 -1162
rect 2820 -1179 2826 -1162
rect 2480 -1182 2826 -1179
rect 2859 -1162 3205 -1159
rect 2859 -1179 2865 -1162
rect 3199 -1179 3205 -1162
rect 2859 -1182 3205 -1179
rect 3238 -1162 3584 -1159
rect 3238 -1179 3244 -1162
rect 3578 -1179 3584 -1162
rect 3238 -1182 3584 -1179
rect 3617 -1162 3963 -1159
rect 3617 -1179 3623 -1162
rect 3957 -1179 3963 -1162
rect 3617 -1182 3963 -1179
rect 3996 -1162 4342 -1159
rect 3996 -1179 4002 -1162
rect 4336 -1179 4342 -1162
rect 3996 -1182 4342 -1179
rect 4375 -1162 4721 -1159
rect 4375 -1179 4381 -1162
rect 4715 -1179 4721 -1162
rect 4375 -1182 4721 -1179
rect 4754 -1162 5100 -1159
rect 4754 -1179 4760 -1162
rect 5094 -1179 5100 -1162
rect 4754 -1182 5100 -1179
rect 5133 -1162 5479 -1159
rect 5133 -1179 5139 -1162
rect 5473 -1179 5479 -1162
rect 5133 -1182 5479 -1179
rect 5512 -1162 5858 -1159
rect 5512 -1179 5518 -1162
rect 5852 -1179 5858 -1162
rect 5512 -1182 5858 -1179
rect 5891 -1162 6237 -1159
rect 5891 -1179 5897 -1162
rect 6231 -1179 6237 -1162
rect 5891 -1182 6237 -1179
rect 6270 -1162 6616 -1159
rect 6270 -1179 6276 -1162
rect 6610 -1179 6616 -1162
rect 6270 -1182 6616 -1179
<< properties >>
string FIXED_BBOX -6689 -1221 6689 1221
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 22.857142857142858 l 3.5 m 1 nf 35 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
