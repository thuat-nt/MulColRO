* NGSPICE file created from user_analog_project_wrapper.ext - technology: sky130A

.subckt sky130_fd_pr__res_generic_m1_SAT4UL m1_n1000_n1057# m1_n1000_1000#
R0 m1_n1000_n1057# m1_n1000_1000# sky130_fd_pr__res_generic_m1 w=10 l=10
.ends

.subckt R_0_125 R1/m1_n1000_n1057# R1/m1_n1000_1000#
XR1 R1/m1_n1000_n1057# R1/m1_n1000_1000# sky130_fd_pr__res_generic_m1_SAT4UL
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_79GNHJ a_4558_n3000# a_n1500_n3097# a_n4616_n3000#
+ a_1558_n3097# a_1500_n3000# w_n4754_n3219# a_n4558_n3097# a_n1558_n3000#
X0 a_1500_n3000# a_n1500_n3097# a_n1558_n3000# w_n4754_n3219# sky130_fd_pr__pfet_01v8_lvt ad=4.35 pd=30.3 as=4.35 ps=30.3 w=30 l=15
X1 a_4558_n3000# a_1558_n3097# a_1500_n3000# w_n4754_n3219# sky130_fd_pr__pfet_01v8_lvt ad=8.7 pd=60.6 as=4.35 ps=30.3 w=30 l=15
X2 a_n1558_n3000# a_n4558_n3097# a_n4616_n3000# w_n4754_n3219# sky130_fd_pr__pfet_01v8_lvt ad=4.35 pd=30.3 as=8.7 ps=60.6 w=30 l=15
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_RM6ABE a_300_n3000# w_n1154_n3219# a_n958_n3097#
+ a_n358_n3000# a_958_n3000# a_n1016_n3000# a_n300_n3097# a_358_n3097#
X0 a_n358_n3000# a_n958_n3097# a_n1016_n3000# w_n1154_n3219# sky130_fd_pr__pfet_01v8_lvt ad=4.35 pd=30.3 as=8.7 ps=60.6 w=30 l=3
X1 a_300_n3000# a_n300_n3097# a_n358_n3000# w_n1154_n3219# sky130_fd_pr__pfet_01v8_lvt ad=4.35 pd=30.3 as=4.35 ps=30.3 w=30 l=3
X2 a_958_n3000# a_358_n3097# a_300_n3000# w_n1154_n3219# sky130_fd_pr__pfet_01v8_lvt ad=8.7 pd=60.6 as=4.35 ps=30.3 w=30 l=3
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_9U978C a_n3087_n1000# a_3029_n1000# a_29_n1088#
+ a_n3189_n1174# a_n3029_n1088# a_n29_n1000#
X0 a_n29_n1000# a_n3029_n1088# a_n3087_n1000# a_n3189_n1174# sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.3 as=2.9 ps=20.6 w=10 l=15
X1 a_3029_n1000# a_29_n1088# a_n29_n1000# a_n3189_n1174# sky130_fd_pr__nfet_01v8_lvt ad=2.9 pd=20.6 as=1.45 ps=10.3 w=10 l=15
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_RM3WAQ a_12536_n2374# a_n1108_n2374# a_11778_n2374#
+ a_1924_n2374# a_n7930_n2374# a_n408_n2286# a_11020_n2374# a_n6414_n2374# a_10262_n2374#
+ a_n5656_n2374# a_11720_n2286# a_10962_n2286# a_n4898_n2374# a_10204_n2286# a_5714_n2374#
+ a_4956_n2374# a_n4140_n2374# a_n3382_n2374# a_n8688_n2374# a_n9446_n2374# a_9504_n2374#
+ a_3440_n2374# a_2682_n2374# a_13236_n2286# a_8746_n2374# a_12478_n2286# a_2624_n2286#
+ a_7988_n2374# a_1166_n2374# a_n7172_n2374# a_1866_n2286# a_1108_n2286# a_7230_n2374#
+ a_6472_n2374# a_7930_n2286# a_6414_n2286# a_5656_n2286# a_4198_n2374# a_4898_n2286#
+ a_408_n2374# a_4140_n2286# a_n1924_n2286# a_n12536_n2286# a_n350_n2374# a_9446_n2286#
+ a_3382_n2286# a_n11778_n2286# a_8688_n2286# a_n11020_n2286# a_n10262_n2286# a_7172_n2286#
+ a_n5714_n2286# a_n4956_n2286# a_n3440_n2286# a_n13294_n2286# a_n11720_n2374# a_n2682_n2286#
+ a_n9504_n2286# a_n10204_n2374# a_n10962_n2374# a_n13396_n2460# a_n1166_n2286# a_n7988_n2286#
+ a_n8746_n2286# a_350_n2286# a_n7230_n2286# a_n6472_n2286# a_n2624_n2374# a_n13236_n2374#
+ a_n4198_n2286# a_n1866_n2374# a_n12478_n2374#
X0 a_n11778_n2286# a_n12478_n2374# a_n12536_n2286# a_n13396_n2460# sky130_fd_pr__nfet_01v8_lvt ad=3.31 pd=23.1 as=3.31 ps=23.1 w=22.9 l=3.5
X1 a_n8746_n2286# a_n9446_n2374# a_n9504_n2286# a_n13396_n2460# sky130_fd_pr__nfet_01v8_lvt ad=3.31 pd=23.1 as=3.31 ps=23.1 w=22.9 l=3.5
X2 a_350_n2286# a_n350_n2374# a_n408_n2286# a_n13396_n2460# sky130_fd_pr__nfet_01v8_lvt ad=3.31 pd=23.1 as=3.31 ps=23.1 w=22.9 l=3.5
X3 a_10204_n2286# a_9504_n2374# a_9446_n2286# a_n13396_n2460# sky130_fd_pr__nfet_01v8_lvt ad=3.31 pd=23.1 as=3.31 ps=23.1 w=22.9 l=3.5
X4 a_n1924_n2286# a_n2624_n2374# a_n2682_n2286# a_n13396_n2460# sky130_fd_pr__nfet_01v8_lvt ad=3.31 pd=23.1 as=3.31 ps=23.1 w=22.9 l=3.5
X5 a_7172_n2286# a_6472_n2374# a_6414_n2286# a_n13396_n2460# sky130_fd_pr__nfet_01v8_lvt ad=3.31 pd=23.1 as=3.31 ps=23.1 w=22.9 l=3.5
X6 a_4898_n2286# a_4198_n2374# a_4140_n2286# a_n13396_n2460# sky130_fd_pr__nfet_01v8_lvt ad=3.31 pd=23.1 as=3.31 ps=23.1 w=22.9 l=3.5
X7 a_12478_n2286# a_11778_n2374# a_11720_n2286# a_n13396_n2460# sky130_fd_pr__nfet_01v8_lvt ad=3.31 pd=23.1 as=3.31 ps=23.1 w=22.9 l=3.5
X8 a_n9504_n2286# a_n10204_n2374# a_n10262_n2286# a_n13396_n2460# sky130_fd_pr__nfet_01v8_lvt ad=3.31 pd=23.1 as=3.31 ps=23.1 w=22.9 l=3.5
X9 a_1108_n2286# a_408_n2374# a_350_n2286# a_n13396_n2460# sky130_fd_pr__nfet_01v8_lvt ad=3.31 pd=23.1 as=3.31 ps=23.1 w=22.9 l=3.5
X10 a_n7988_n2286# a_n8688_n2374# a_n8746_n2286# a_n13396_n2460# sky130_fd_pr__nfet_01v8_lvt ad=3.31 pd=23.1 as=3.31 ps=23.1 w=22.9 l=3.5
X11 a_9446_n2286# a_8746_n2374# a_8688_n2286# a_n13396_n2460# sky130_fd_pr__nfet_01v8_lvt ad=3.31 pd=23.1 as=3.31 ps=23.1 w=22.9 l=3.5
X12 a_n1166_n2286# a_n1866_n2374# a_n1924_n2286# a_n13396_n2460# sky130_fd_pr__nfet_01v8_lvt ad=3.31 pd=23.1 as=3.31 ps=23.1 w=22.9 l=3.5
X13 a_11720_n2286# a_11020_n2374# a_10962_n2286# a_n13396_n2460# sky130_fd_pr__nfet_01v8_lvt ad=3.31 pd=23.1 as=3.31 ps=23.1 w=22.9 l=3.5
X14 a_2624_n2286# a_1924_n2374# a_1866_n2286# a_n13396_n2460# sky130_fd_pr__nfet_01v8_lvt ad=3.31 pd=23.1 as=3.31 ps=23.1 w=22.9 l=3.5
X15 a_n5714_n2286# a_n6414_n2374# a_n6472_n2286# a_n13396_n2460# sky130_fd_pr__nfet_01v8_lvt ad=3.31 pd=23.1 as=3.31 ps=23.1 w=22.9 l=3.5
X16 a_n3440_n2286# a_n4140_n2374# a_n4198_n2286# a_n13396_n2460# sky130_fd_pr__nfet_01v8_lvt ad=3.31 pd=23.1 as=3.31 ps=23.1 w=22.9 l=3.5
X17 a_n2682_n2286# a_n3382_n2374# a_n3440_n2286# a_n13396_n2460# sky130_fd_pr__nfet_01v8_lvt ad=3.31 pd=23.1 as=3.31 ps=23.1 w=22.9 l=3.5
X18 a_4140_n2286# a_3440_n2374# a_3382_n2286# a_n13396_n2460# sky130_fd_pr__nfet_01v8_lvt ad=3.31 pd=23.1 as=3.31 ps=23.1 w=22.9 l=3.5
X19 a_1866_n2286# a_1166_n2374# a_1108_n2286# a_n13396_n2460# sky130_fd_pr__nfet_01v8_lvt ad=3.31 pd=23.1 as=3.31 ps=23.1 w=22.9 l=3.5
X20 a_8688_n2286# a_7988_n2374# a_7930_n2286# a_n13396_n2460# sky130_fd_pr__nfet_01v8_lvt ad=3.31 pd=23.1 as=3.31 ps=23.1 w=22.9 l=3.5
X21 a_10962_n2286# a_10262_n2374# a_10204_n2286# a_n13396_n2460# sky130_fd_pr__nfet_01v8_lvt ad=3.31 pd=23.1 as=3.31 ps=23.1 w=22.9 l=3.5
X22 a_n11020_n2286# a_n11720_n2374# a_n11778_n2286# a_n13396_n2460# sky130_fd_pr__nfet_01v8_lvt ad=3.31 pd=23.1 as=3.31 ps=23.1 w=22.9 l=3.5
X23 a_n10262_n2286# a_n10962_n2374# a_n11020_n2286# a_n13396_n2460# sky130_fd_pr__nfet_01v8_lvt ad=3.31 pd=23.1 as=3.31 ps=23.1 w=22.9 l=3.5
X24 a_n4956_n2286# a_n5656_n2374# a_n5714_n2286# a_n13396_n2460# sky130_fd_pr__nfet_01v8_lvt ad=3.31 pd=23.1 as=3.31 ps=23.1 w=22.9 l=3.5
X25 a_6414_n2286# a_5714_n2374# a_5656_n2286# a_n13396_n2460# sky130_fd_pr__nfet_01v8_lvt ad=3.31 pd=23.1 as=3.31 ps=23.1 w=22.9 l=3.5
X26 a_n12536_n2286# a_n13236_n2374# a_n13294_n2286# a_n13396_n2460# sky130_fd_pr__nfet_01v8_lvt ad=3.31 pd=23.1 as=6.63 ps=46.3 w=22.9 l=3.5
X27 a_3382_n2286# a_2682_n2374# a_2624_n2286# a_n13396_n2460# sky130_fd_pr__nfet_01v8_lvt ad=3.31 pd=23.1 as=3.31 ps=23.1 w=22.9 l=3.5
X28 a_n6472_n2286# a_n7172_n2374# a_n7230_n2286# a_n13396_n2460# sky130_fd_pr__nfet_01v8_lvt ad=3.31 pd=23.1 as=3.31 ps=23.1 w=22.9 l=3.5
X29 a_7930_n2286# a_7230_n2374# a_7172_n2286# a_n13396_n2460# sky130_fd_pr__nfet_01v8_lvt ad=3.31 pd=23.1 as=3.31 ps=23.1 w=22.9 l=3.5
X30 a_n408_n2286# a_n1108_n2374# a_n1166_n2286# a_n13396_n2460# sky130_fd_pr__nfet_01v8_lvt ad=3.31 pd=23.1 as=3.31 ps=23.1 w=22.9 l=3.5
X31 a_13236_n2286# a_12536_n2374# a_12478_n2286# a_n13396_n2460# sky130_fd_pr__nfet_01v8_lvt ad=6.63 pd=46.3 as=3.31 ps=23.1 w=22.9 l=3.5
X32 a_n7230_n2286# a_n7930_n2374# a_n7988_n2286# a_n13396_n2460# sky130_fd_pr__nfet_01v8_lvt ad=3.31 pd=23.1 as=3.31 ps=23.1 w=22.9 l=3.5
X33 a_n4198_n2286# a_n4898_n2374# a_n4956_n2286# a_n13396_n2460# sky130_fd_pr__nfet_01v8_lvt ad=3.31 pd=23.1 as=3.31 ps=23.1 w=22.9 l=3.5
X34 a_5656_n2286# a_4956_n2374# a_4898_n2286# a_n13396_n2460# sky130_fd_pr__nfet_01v8_lvt ad=3.31 pd=23.1 as=3.31 ps=23.1 w=22.9 l=3.5
.ends

.subckt diffamp PCAS REF PIX GM_BIAS VDD VSS OUT
XXM1 m1_35096_n15744# m1_32048_n23188# VDD m1_32048_n23188# VDD VDD m1_32048_n23188#
+ m1_35096_n15744# sky130_fd_pr__pfet_01v8_lvt_79GNHJ
XXM2 OUT VDD PCAS m1_32020_n12120# m1_32020_n12120# OUT PCAS PCAS sky130_fd_pr__pfet_01v8_lvt_RM6ABE
XXM3 m1_31296_n26048# m1_31296_n26048# GM_BIAS VSS GM_BIAS VSS sky130_fd_pr__nfet_01v8_lvt_9U978C
XXM4 m1_32048_n23188# VDD PCAS m1_35096_n15744# m1_35096_n15744# m1_32048_n23188#
+ PCAS PCAS sky130_fd_pr__pfet_01v8_lvt_RM6ABE
XXM5 PIX PIX PIX PIX PIX m1_31296_n26048# PIX PIX PIX PIX m1_31296_n26048# OUT PIX
+ m1_31296_n26048# PIX PIX PIX PIX PIX PIX PIX PIX PIX m1_31296_n26048# PIX OUT m1_31296_n26048#
+ PIX PIX PIX OUT m1_31296_n26048# PIX PIX OUT OUT m1_31296_n26048# PIX OUT PIX m1_31296_n26048#
+ m1_31296_n26048# m1_31296_n26048# PIX OUT OUT OUT m1_31296_n26048# m1_31296_n26048#
+ OUT m1_31296_n26048# OUT m1_31296_n26048# m1_31296_n26048# OUT PIX OUT m1_31296_n26048#
+ PIX PIX VSS OUT m1_31296_n26048# OUT OUT OUT m1_31296_n26048# PIX PIX OUT PIX PIX
+ sky130_fd_pr__nfet_01v8_lvt_RM3WAQ
XXM6 REF REF REF REF REF m1_32048_n23188# REF REF REF REF m1_32048_n23188# m1_31296_n26048#
+ REF m1_32048_n23188# REF REF REF REF REF REF REF REF REF m1_32048_n23188# REF m1_31296_n26048#
+ m1_32048_n23188# REF REF REF m1_31296_n26048# m1_32048_n23188# REF REF m1_31296_n26048#
+ m1_31296_n26048# m1_32048_n23188# REF m1_31296_n26048# REF m1_32048_n23188# m1_32048_n23188#
+ m1_32048_n23188# REF m1_31296_n26048# m1_31296_n26048# m1_31296_n26048# m1_32048_n23188#
+ m1_32048_n23188# m1_31296_n26048# m1_32048_n23188# m1_31296_n26048# m1_32048_n23188#
+ m1_32048_n23188# m1_31296_n26048# REF m1_31296_n26048# m1_32048_n23188# REF REF
+ VSS m1_31296_n26048# m1_32048_n23188# m1_31296_n26048# m1_31296_n26048# m1_31296_n26048#
+ m1_32048_n23188# REF REF m1_31296_n26048# REF REF sky130_fd_pr__nfet_01v8_lvt_RM3WAQ
XXM8 VDD m1_32048_n23188# m1_32020_n12120# m1_32048_n23188# m1_32020_n12120# VDD m1_32048_n23188#
+ VDD sky130_fd_pr__pfet_01v8_lvt_79GNHJ
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_6LX62X a_35_n100# a_n35_n188# a_n195_n274# a_n93_n100#
X0 a_35_n100# a_n35_n188# a_n93_n100# a_n195_n274# sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.35
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_4QFWD3 a_n93_n200# a_n35_n297# a_35_n200# w_n231_n419#
X0 a_35_n200# a_n35_n297# a_n93_n200# w_n231_n419# sky130_fd_pr__pfet_01v8_lvt ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.35
.ends

.subckt not out in VDD VSS
XXM1 out in VSS VSS sky130_fd_pr__nfet_01v8_lvt_6LX62X
XXM10 VDD in out VDD sky130_fd_pr__pfet_01v8_lvt_4QFWD3
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_ER7S26 a_n221_n4000# a_93_n4097# a_35_n4000# a_291_n4000#
+ a_n349_n4000# a_221_n4097# a_n163_n4097# w_n487_n4219# a_163_n4000# a_n93_n4000#
+ a_n291_n4097# a_n35_n4097#
X0 a_163_n4000# a_93_n4097# a_35_n4000# w_n487_n4219# sky130_fd_pr__pfet_01v8_lvt ad=5.8 pd=40.3 as=5.8 ps=40.3 w=40 l=0.35
X1 a_35_n4000# a_n35_n4097# a_n93_n4000# w_n487_n4219# sky130_fd_pr__pfet_01v8_lvt ad=5.8 pd=40.3 as=5.8 ps=40.3 w=40 l=0.35
X2 a_n221_n4000# a_n291_n4097# a_n349_n4000# w_n487_n4219# sky130_fd_pr__pfet_01v8_lvt ad=5.8 pd=40.3 as=11.6 ps=80.6 w=40 l=0.35
X3 a_n93_n4000# a_n163_n4097# a_n221_n4000# w_n487_n4219# sky130_fd_pr__pfet_01v8_lvt ad=5.8 pd=40.3 as=5.8 ps=40.3 w=40 l=0.35
X4 a_291_n4000# a_221_n4097# a_163_n4000# w_n487_n4219# sky130_fd_pr__pfet_01v8_lvt ad=11.6 pd=80.6 as=5.8 ps=40.3 w=40 l=0.35
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_4833E6 a_n1016_n4000# a_1016_n4088# G D B a_n958_n4088#
+ a_300_n4000# a_n1616_n4088# S a_358_n4088# a_n358_n4000# a_958_n4000#
X0 a_n1016_n4000# a_n1616_n4088# D B sky130_fd_pr__nfet_01v8_lvt ad=5.8 pd=40.3 as=11.6 ps=80.6 w=40 l=3
X1 a_n358_n4000# a_n958_n4088# a_n1016_n4000# B sky130_fd_pr__nfet_01v8_lvt ad=5.8 pd=40.3 as=5.8 ps=40.3 w=40 l=3
X2 S a_1016_n4088# a_958_n4000# B sky130_fd_pr__nfet_01v8_lvt ad=11.6 pd=80.6 as=5.8 ps=40.3 w=40 l=3
X3 a_300_n4000# G a_n358_n4000# B sky130_fd_pr__nfet_01v8_lvt ad=5.8 pd=40.3 as=5.8 ps=40.3 w=40 l=3
X4 a_958_n4000# a_358_n4088# a_300_n4000# B sky130_fd_pr__nfet_01v8_lvt ad=5.8 pd=40.3 as=5.8 ps=40.3 w=40 l=3
.ends

.subckt switch in out toggle VSS VDD
Xx1 x1/out toggle VDD VSS not
XXM26 in x1/out in in out x1/out x1/out out out out x1/out x1/out sky130_fd_pr__pfet_01v8_lvt_ER7S26
XXM1 out toggle toggle in VSS toggle out toggle out toggle in in sky130_fd_pr__nfet_01v8_lvt_4833E6
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_T4BG7Y a_200_n5000# a_n360_n5174# a_n200_n5088#
+ a_n258_n5000#
X0 a_200_n5000# a_n200_n5088# a_n258_n5000# a_n360_n5174# sky130_fd_pr__nfet_01v8_lvt ad=14.5 pd=101 as=14.5 ps=101 w=50 l=2
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_B5Z988 a_n1000_n1097# w_n1196_n1219# a_1000_n1000#
+ a_n1058_n1000#
X0 a_1000_n1000# a_n1000_n1097# a_n1058_n1000# w_n1196_n1219# sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.6 as=2.9 ps=20.6 w=10 l=10
.ends

.subckt curr_mir Vtune VDD Ib VSS
XXM1 VSS VSS m1_1036_6332# m1_1036_6332# sky130_fd_pr__nfet_01v8_lvt_T4BG7Y
XXM2 VSS VSS m1_1036_6332# Ib sky130_fd_pr__nfet_01v8_lvt_T4BG7Y
XXM10 Vtune VDD VDD m1_1036_6332# sky130_fd_pr__pfet_01v8_lvt_B5Z988
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_CEE7V5 G D B a_358_n597# a_n300_n597# a_958_n500#
+ S a_300_n500#
X0 S G D B sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.29 as=1.45 ps=10.6 w=5 l=3
X1 a_300_n500# a_n300_n597# S B sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=3
X2 a_958_n500# a_358_n597# a_300_n500# B sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.6 as=0.725 ps=5.29 w=5 l=3
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_8WRJS5 a_29_n347# G D B a_629_n250# a_n629_n347#
+ a_687_n347# a_n29_n250# a_1287_n250# S
X0 a_1287_n250# a_687_n347# a_629_n250# B sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.363 ps=2.79 w=2.5 l=3
X1 a_629_n250# a_29_n347# a_n29_n250# B sky130_fd_pr__pfet_01v8_lvt ad=0.363 pd=2.79 as=0.363 ps=2.79 w=2.5 l=3
X2 a_n29_n250# a_n629_n347# S B sky130_fd_pr__pfet_01v8_lvt ad=0.363 pd=2.79 as=0.363 ps=2.79 w=2.5 l=3
X3 S G D B sky130_fd_pr__pfet_01v8_lvt ad=0.363 pd=2.79 as=0.725 ps=5.58 w=2.5 l=3
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_HZEGLD a_958_n1600# G a_1016_n1688# D B a_n958_n1688#
+ a_1616_n1600# a_300_n1600# a_n300_n1688# S a_358_n1688# a_n358_n1600#
X0 a_300_n1600# a_n300_n1688# a_n358_n1600# B sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.3 as=2.32 ps=16.3 w=16 l=3
X1 a_958_n1600# a_358_n1688# a_300_n1600# B sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.3 as=2.32 ps=16.3 w=16 l=3
X2 S G D B sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.3 as=4.64 ps=32.6 w=16 l=3
X3 a_n358_n1600# a_n958_n1688# S B sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.3 as=2.32 ps=16.3 w=16 l=3
X4 a_1616_n1600# a_1016_n1688# a_958_n1600# B sky130_fd_pr__nfet_01v8_lvt ad=4.64 pd=32.6 as=2.32 ps=16.3 w=16 l=3
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_RFVHWA G D B S
X0 S G D B sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=3
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_7233E2 G D B S
X0 S G D B sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.6 as=2.32 ps=16.6 w=8 l=3
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_CEAZV5 G a_29_n597# D B a_629_n500# S
X0 a_629_n500# a_29_n597# S B sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.6 as=0.725 ps=5.29 w=5 l=3
X1 S G D B sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.29 as=1.45 ps=10.6 w=5 l=3
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_ZYFHHD c0 c1
X0 c0 c1 sky130_fd_pr__cap_mim_m3_1 l=4 w=2
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_LEXMNV G D a_n958_n2097# w_n1812_n2219# a_n358_n2000#
+ a_958_n2000# a_n300_n2097# a_1616_n2000# a_358_n2097# S a_300_n2000# a_1016_n2097#
X0 S G D w_n1812_n2219# sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.3 as=5.8 ps=40.6 w=20 l=3
X1 a_n358_n2000# a_n958_n2097# S w_n1812_n2219# sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=3
X2 a_1616_n2000# a_1016_n2097# a_958_n2000# w_n1812_n2219# sky130_fd_pr__pfet_01v8_lvt ad=5.8 pd=40.6 as=2.9 ps=20.3 w=20 l=3
X3 a_300_n2000# a_n300_n2097# a_n358_n2000# w_n1812_n2219# sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=3
X4 a_958_n2000# a_358_n2097# a_300_n2000# w_n1812_n2219# sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.3 as=2.9 ps=20.3 w=20 l=3
.ends

.subckt opamp opbias inp inn VDD out VSS
XXM14 inn XM5/G VDD inn inn XM26/D XM26/D XM5/G sky130_fd_pr__pfet_01v8_lvt_CEE7V5
XXM15 inp XM2/G VDD inp inp XM26/D XM26/D XM2/G sky130_fd_pr__pfet_01v8_lvt_CEE7V5
XXM26 opbias opbias XM26/D VDD VDD opbias opbias XM26/D XM26/D VDD sky130_fd_pr__pfet_01v8_lvt_8WRJS5
XXM17 out XM2/G XM2/G out VSS XM2/G VSS VSS XM2/G VSS XM2/G out sky130_fd_pr__nfet_01v8_lvt_HZEGLD
XXM19 XM5/G XM5/G VSS VSS sky130_fd_pr__nfet_01v8_lvt_RFVHWA
XXM2 XM2/G XM4/G VSS VSS sky130_fd_pr__nfet_01v8_lvt_7233E2
XXM3 XM4/G XM4/G XM4/G VDD XM4/G VDD sky130_fd_pr__pfet_01v8_lvt_CEAZV5
XXM4 XM4/G XM4/G XM5/D VDD XM5/D VDD sky130_fd_pr__pfet_01v8_lvt_CEAZV5
XXM5 XM5/G XM5/D VSS VSS sky130_fd_pr__nfet_01v8_lvt_7233E2
XXC1 XM5/D out sky130_fd_pr__cap_mim_m3_1_ZYFHHD
XXC2 out XM2/G sky130_fd_pr__cap_mim_m3_1_ZYFHHD
XXM20 XM5/G XM2/G VSS VSS sky130_fd_pr__nfet_01v8_lvt_RFVHWA
XXM10 XM5/D out XM5/D VDD out out XM5/D VDD XM5/D VDD VDD XM5/D sky130_fd_pr__pfet_01v8_lvt_LEXMNV
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_3HBNLG c0 c1
X0 c0 c1 sky130_fd_pr__cap_mim_m3_1 l=30 w=30
.ends

.subckt integrator sw4 sw3 rst sw2 sw1 opbias en Vtune intin VDD intout VSS
Xx1 x9/in x1/out sw1 VSS VDD switch
Xx3 Vtune VDD intin VSS curr_mir
Xx2 intin x9/in x7/out VSS VDD switch
Xx4 opbias VSS x9/in VDD intout VSS opamp
Xx5 x9/in intout rst VSS VDD switch
Xx6 intin VSS en VSS VDD switch
Xx7 x7/out en VDD VSS not
Xx8 x9/in x8/out sw4 VSS VDD switch
Xx9 x9/in x9/out sw2 VSS VDD switch
XXC1 x1/out intout sky130_fd_pr__cap_mim_m3_1_3HBNLG
XXC2 x9/out intout sky130_fd_pr__cap_mim_m3_1_3HBNLG
XXC3 XC3/c0 intout sky130_fd_pr__cap_mim_m3_1_3HBNLG
Xx10 x9/in XC3/c0 sw3 VSS VDD switch
XXC4 x8/out intout sky130_fd_pr__cap_mim_m3_1_3HBNLG
.ends

.subckt mux2_1 SEL0 IN1 IN0 VDD OUT VSS
Xx1 x1/out SEL0 VDD VSS not
Xx5 IN0 OUT x1/out VSS VDD switch
Xx6 IN1 OUT SEL0 VSS VDD switch
.ends

.subckt buffer opbias in out VDD VSS
Xx1 opbias in out VDD out VSS opamp
.ends

.subckt ColROs VDD AIn0 AIn1 AIn2 AIn3 AIn4 AIn5 REG0 REG1 REG2 REG3 REG4 REG5 REG6
+ AOut VSS
Xx1 AIn3 AIn0 AIn1 AIn2 VDD VSS x3/IN0 diffamp
Xx2 REG5 REG4 REG1 REG3 REG2 AIn4 REG0 AIn5 x3/IN0 VDD x3/IN1 VSS integrator
Xx3 REG6 x3/IN1 x3/IN0 VDD x7/in VSS mux2_1
Xx7 AIn4 x7/in AOut VDD VSS buffer
.ends

.subckt MulColROs VDD AOut[3] AOut[2] AOut[1] AOut[0] REG6 REG5 REG4 REG3 REG2 REG1
+ REG0 AIn5 AIn4 AIn3 AIn2 AIn0 AIn[3] AIn[2] AIn[1] AIn[0] VSS
XxMulColROs[3] VDD AIn0 AIn[3] AIn2 AIn3 AIn4 AIn5 REG0 REG1 REG2 REG3 REG4 REG5 REG6
+ AOut[3] VSS ColROs
XxMulColROs[2] VDD AIn0 AIn[2] AIn2 AIn3 AIn4 AIn5 REG0 REG1 REG2 REG3 REG4 REG5 REG6
+ AOut[2] VSS ColROs
XxMulColROs[1] VDD AIn0 AIn[1] AIn2 AIn3 AIn4 AIn5 REG0 REG1 REG2 REG3 REG4 REG5 REG6
+ AOut[1] VSS ColROs
XxMulColROs[0] VDD AIn0 AIn[0] AIn2 AIn3 AIn4 AIn5 REG0 REG1 REG2 REG3 REG4 REG5 REG6
+ AOut[0] VSS ColROs
.ends

.subckt sky130_fd_pr__res_generic_m3_DPAT6Q m3_n1100_n87# m3_n1100_30#
R0 m3_n1100_n87# m3_n1100_30# sky130_fd_pr__res_generic_m3 w=11 l=0.3
.ends

.subckt user_analog_project_wrapper gpio_analog[0] gpio_analog[10] gpio_analog[11]
+ gpio_analog[12] gpio_analog[13] gpio_analog[14] gpio_analog[15] gpio_analog[16]
+ gpio_analog[17] gpio_analog[1] gpio_analog[2] gpio_analog[3] gpio_analog[4] gpio_analog[5]
+ gpio_analog[6] gpio_analog[7] gpio_analog[8] gpio_analog[9] gpio_noesd[0] gpio_noesd[10]
+ gpio_noesd[11] gpio_noesd[12] gpio_noesd[13] gpio_noesd[14] gpio_noesd[15] gpio_noesd[16]
+ gpio_noesd[17] gpio_noesd[1] gpio_noesd[2] gpio_noesd[3] gpio_noesd[4] gpio_noesd[5]
+ gpio_noesd[6] gpio_noesd[7] gpio_noesd[8] gpio_noesd[9] io_analog[0] io_analog[10]
+ io_analog[1] io_analog[2] io_analog[3] io_analog[7] io_analog[8] io_analog[9] io_analog[4]
+ io_analog[5] io_analog[6] io_clamp_high[0] io_clamp_high[1] io_clamp_high[2] io_clamp_low[0]
+ io_clamp_low[1] io_clamp_low[2] io_in[0] io_in[10] io_in[11] io_in[12] io_in[13]
+ io_in[14] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21]
+ io_in[22] io_in[23] io_in[24] io_in[25] io_in[26] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_in[8] io_in[9] io_in_3v3[0] io_in_3v3[10] io_in_3v3[11] io_in_3v3[12]
+ io_in_3v3[13] io_in_3v3[14] io_in_3v3[15] io_in_3v3[16] io_in_3v3[17] io_in_3v3[18]
+ io_in_3v3[19] io_in_3v3[1] io_in_3v3[20] io_in_3v3[21] io_in_3v3[22] io_in_3v3[23]
+ io_in_3v3[24] io_in_3v3[25] io_in_3v3[26] io_in_3v3[2] io_in_3v3[3] io_in_3v3[4]
+ io_in_3v3[5] io_in_3v3[6] io_in_3v3[7] io_in_3v3[8] io_in_3v3[9] io_oeb[0] io_oeb[10]
+ io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18]
+ io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25]
+ io_oeb[26] io_oeb[2] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8]
+ io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15]
+ io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22]
+ io_out[23] io_out[24] io_out[25] io_out[26] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] io_out[8] io_out[9] la_data_in[0] la_data_in[100] la_data_in[101]
+ la_data_in[102] la_data_in[103] la_data_in[104] la_data_in[105] la_data_in[106]
+ la_data_in[107] la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110] la_data_in[111]
+ la_data_in[112] la_data_in[113] la_data_in[114] la_data_in[115] la_data_in[116]
+ la_data_in[117] la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120] la_data_in[121]
+ la_data_in[122] la_data_in[123] la_data_in[124] la_data_in[125] la_data_in[126]
+ la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15] la_data_in[16]
+ la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20] la_data_in[21]
+ la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26] la_data_in[27]
+ la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31] la_data_in[32]
+ la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37] la_data_in[38]
+ la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42] la_data_in[43]
+ la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48] la_data_in[49]
+ la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53] la_data_in[54]
+ la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59] la_data_in[5]
+ la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64] la_data_in[65]
+ la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6] la_data_in[70]
+ la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75] la_data_in[76]
+ la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80] la_data_in[81]
+ la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86] la_data_in[87]
+ la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91] la_data_in[92]
+ la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97] la_data_in[98]
+ la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101] la_data_out[102]
+ la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106] la_data_out[107]
+ la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110] la_data_out[111]
+ la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115] la_data_out[116]
+ la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11] la_data_out[120]
+ la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124] la_data_out[125]
+ la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13] la_data_out[14]
+ la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19]
+ la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24]
+ la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29]
+ la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34]
+ la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39]
+ la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44]
+ la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49]
+ la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54]
+ la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59]
+ la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[64]
+ la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68] la_data_out[69]
+ la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73] la_data_out[74]
+ la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78] la_data_out[79]
+ la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83] la_data_out[84]
+ la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88] la_data_out[89]
+ la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93] la_data_out[94]
+ la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98] la_data_out[99]
+ la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102] la_oenb[103] la_oenb[104]
+ la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109] la_oenb[10] la_oenb[110]
+ la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115] la_oenb[116] la_oenb[117]
+ la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121] la_oenb[122] la_oenb[123]
+ la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33]
+ la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3]
+ la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46]
+ la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52]
+ la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59]
+ la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[64] la_oenb[65]
+ la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6] la_oenb[70] la_oenb[71]
+ la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76] la_oenb[77] la_oenb[78]
+ la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82] la_oenb[83] la_oenb[84]
+ la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89] la_oenb[8] la_oenb[90]
+ la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95] la_oenb[96] la_oenb[97]
+ la_oenb[98] la_oenb[99] la_oenb[9] user_clock2 user_irq[0] user_irq[1] user_irq[2]
+ vccd1 vccd2 vdda1 vdda2 vssa1 vssa2 vssd1 vssd2 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0]
+ wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15]
+ wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20]
+ wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26]
+ wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31]
+ wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9]
+ wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14]
+ wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1]
+ wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25]
+ wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30]
+ wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8]
+ wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13]
+ wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19]
+ wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24]
+ wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2]
+ wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6]
+ wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3]
+ wbs_stb_i wbs_we_i
XXR[15] vccd1 io_oeb[15] R_0_125
Xx1 vccd1 io_analog[3] io_analog[2] io_analog[1] io_analog[0] io_in[0] io_in[1] io_in[2]
+ io_in[3] io_in[4] io_in[5] io_in[6] gpio_analog[8] gpio_analog[7] gpio_analog[6]
+ gpio_analog[5] gpio_analog[0] gpio_analog[4] gpio_analog[3] gpio_analog[2] gpio_analog[1]
+ vssd1 MulColROs
XXR[14] vccd1 io_oeb[14] R_0_125
XR1 vssd1 io_clamp_low[2] sky130_fd_pr__res_generic_m3_DPAT6Q
XXR[13] vccd1 io_oeb[13] R_0_125
XR2 vssd1 io_clamp_high[2] sky130_fd_pr__res_generic_m3_DPAT6Q
XXR[12] vccd1 io_oeb[12] R_0_125
XXR[11] vccd1 io_oeb[11] R_0_125
XR4 vssd1 io_clamp_low[1] sky130_fd_pr__res_generic_m3_DPAT6Q
XXR[10] vccd1 io_oeb[10] R_0_125
XR5 vssd1 io_clamp_high[1] sky130_fd_pr__res_generic_m3_DPAT6Q
XR6 vssd1 io_clamp_low[0] sky130_fd_pr__res_generic_m3_DPAT6Q
XR7 vssd1 io_clamp_high[0] sky130_fd_pr__res_generic_m3_DPAT6Q
XXR[9] vccd1 io_oeb[9] R_0_125
XXR[8] vccd1 io_oeb[8] R_0_125
XXR[7] vccd1 io_oeb[7] R_0_125
XXR[6] vccd1 io_oeb[6] R_0_125
XXR[5] vccd1 io_oeb[5] R_0_125
XXR[4] vccd1 io_oeb[4] R_0_125
XXR[3] vccd1 io_oeb[3] R_0_125
XXR[2] vccd1 io_oeb[2] R_0_125
XXR[1] vccd1 io_oeb[1] R_0_125
XXR[0] vccd1 io_oeb[0] R_0_125
.ends

