magic
tech sky130A
magscale 1 2
timestamp 1698123815
<< error_p >>
rect -287 4081 -225 4087
rect -159 4081 -97 4087
rect -31 4081 31 4087
rect 97 4081 159 4087
rect 225 4081 287 4087
rect -287 4047 -275 4081
rect -159 4047 -147 4081
rect -31 4047 -19 4081
rect 97 4047 109 4081
rect 225 4047 237 4081
rect -287 4041 -225 4047
rect -159 4041 -97 4047
rect -31 4041 31 4047
rect 97 4041 159 4047
rect 225 4041 287 4047
rect -287 -4047 -225 -4041
rect -159 -4047 -97 -4041
rect -31 -4047 31 -4041
rect 97 -4047 159 -4041
rect 225 -4047 287 -4041
rect -287 -4081 -275 -4047
rect -159 -4081 -147 -4047
rect -31 -4081 -19 -4047
rect 97 -4081 109 -4047
rect 225 -4081 237 -4047
rect -287 -4087 -225 -4081
rect -159 -4087 -97 -4081
rect -31 -4087 31 -4081
rect 97 -4087 159 -4081
rect 225 -4087 287 -4081
<< nwell >>
rect -487 -4219 487 4219
<< pmoslvt >>
rect -291 -4000 -221 4000
rect -163 -4000 -93 4000
rect -35 -4000 35 4000
rect 93 -4000 163 4000
rect 221 -4000 291 4000
<< pdiff >>
rect -349 3988 -291 4000
rect -349 -3988 -337 3988
rect -303 -3988 -291 3988
rect -349 -4000 -291 -3988
rect -221 3988 -163 4000
rect -221 -3988 -209 3988
rect -175 -3988 -163 3988
rect -221 -4000 -163 -3988
rect -93 3988 -35 4000
rect -93 -3988 -81 3988
rect -47 -3988 -35 3988
rect -93 -4000 -35 -3988
rect 35 3988 93 4000
rect 35 -3988 47 3988
rect 81 -3988 93 3988
rect 35 -4000 93 -3988
rect 163 3988 221 4000
rect 163 -3988 175 3988
rect 209 -3988 221 3988
rect 163 -4000 221 -3988
rect 291 3988 349 4000
rect 291 -3988 303 3988
rect 337 -3988 349 3988
rect 291 -4000 349 -3988
<< pdiffc >>
rect -337 -3988 -303 3988
rect -209 -3988 -175 3988
rect -81 -3988 -47 3988
rect 47 -3988 81 3988
rect 175 -3988 209 3988
rect 303 -3988 337 3988
<< nsubdiff >>
rect -451 4149 -355 4183
rect 355 4149 451 4183
rect -451 4087 -417 4149
rect 417 4087 451 4149
rect -451 -4149 -417 -4087
rect 417 -4149 451 -4087
rect -451 -4183 -355 -4149
rect 355 -4183 451 -4149
<< nsubdiffcont >>
rect -355 4149 355 4183
rect -451 -4087 -417 4087
rect 417 -4087 451 4087
rect -355 -4183 355 -4149
<< poly >>
rect -291 4081 -221 4097
rect -291 4047 -275 4081
rect -237 4047 -221 4081
rect -291 4000 -221 4047
rect -163 4081 -93 4097
rect -163 4047 -147 4081
rect -109 4047 -93 4081
rect -163 4000 -93 4047
rect -35 4081 35 4097
rect -35 4047 -19 4081
rect 19 4047 35 4081
rect -35 4000 35 4047
rect 93 4081 163 4097
rect 93 4047 109 4081
rect 147 4047 163 4081
rect 93 4000 163 4047
rect 221 4081 291 4097
rect 221 4047 237 4081
rect 275 4047 291 4081
rect 221 4000 291 4047
rect -291 -4047 -221 -4000
rect -291 -4081 -275 -4047
rect -237 -4081 -221 -4047
rect -291 -4097 -221 -4081
rect -163 -4047 -93 -4000
rect -163 -4081 -147 -4047
rect -109 -4081 -93 -4047
rect -163 -4097 -93 -4081
rect -35 -4047 35 -4000
rect -35 -4081 -19 -4047
rect 19 -4081 35 -4047
rect -35 -4097 35 -4081
rect 93 -4047 163 -4000
rect 93 -4081 109 -4047
rect 147 -4081 163 -4047
rect 93 -4097 163 -4081
rect 221 -4047 291 -4000
rect 221 -4081 237 -4047
rect 275 -4081 291 -4047
rect 221 -4097 291 -4081
<< polycont >>
rect -275 4047 -237 4081
rect -147 4047 -109 4081
rect -19 4047 19 4081
rect 109 4047 147 4081
rect 237 4047 275 4081
rect -275 -4081 -237 -4047
rect -147 -4081 -109 -4047
rect -19 -4081 19 -4047
rect 109 -4081 147 -4047
rect 237 -4081 275 -4047
<< locali >>
rect -451 4149 -355 4183
rect 355 4149 451 4183
rect -451 4087 -417 4149
rect 417 4087 451 4149
rect -291 4047 -275 4081
rect -237 4047 -221 4081
rect -163 4047 -147 4081
rect -109 4047 -93 4081
rect -35 4047 -19 4081
rect 19 4047 35 4081
rect 93 4047 109 4081
rect 147 4047 163 4081
rect 221 4047 237 4081
rect 275 4047 291 4081
rect -337 3988 -303 4004
rect -337 -4004 -303 -3988
rect -209 3988 -175 4004
rect -209 -4004 -175 -3988
rect -81 3988 -47 4004
rect -81 -4004 -47 -3988
rect 47 3988 81 4004
rect 47 -4004 81 -3988
rect 175 3988 209 4004
rect 175 -4004 209 -3988
rect 303 3988 337 4004
rect 303 -4004 337 -3988
rect -291 -4081 -275 -4047
rect -237 -4081 -221 -4047
rect -163 -4081 -147 -4047
rect -109 -4081 -93 -4047
rect -35 -4081 -19 -4047
rect 19 -4081 35 -4047
rect 93 -4081 109 -4047
rect 147 -4081 163 -4047
rect 221 -4081 237 -4047
rect 275 -4081 291 -4047
rect -451 -4149 -417 -4087
rect 417 -4149 451 -4087
rect -451 -4183 -355 -4149
rect 355 -4183 451 -4149
<< viali >>
rect -275 4047 -237 4081
rect -147 4047 -109 4081
rect -19 4047 19 4081
rect 109 4047 147 4081
rect 237 4047 275 4081
rect -337 -3988 -303 3988
rect -209 -3988 -175 3988
rect -81 -3988 -47 3988
rect 47 -3988 81 3988
rect 175 -3988 209 3988
rect 303 -3988 337 3988
rect -275 -4081 -237 -4047
rect -147 -4081 -109 -4047
rect -19 -4081 19 -4047
rect 109 -4081 147 -4047
rect 237 -4081 275 -4047
<< metal1 >>
rect -287 4081 -225 4087
rect -287 4047 -275 4081
rect -237 4047 -225 4081
rect -287 4041 -225 4047
rect -159 4081 -97 4087
rect -159 4047 -147 4081
rect -109 4047 -97 4081
rect -159 4041 -97 4047
rect -31 4081 31 4087
rect -31 4047 -19 4081
rect 19 4047 31 4081
rect -31 4041 31 4047
rect 97 4081 159 4087
rect 97 4047 109 4081
rect 147 4047 159 4081
rect 97 4041 159 4047
rect 225 4081 287 4087
rect 225 4047 237 4081
rect 275 4047 287 4081
rect 225 4041 287 4047
rect -343 3988 -297 4000
rect -343 -3988 -337 3988
rect -303 -3988 -297 3988
rect -343 -4000 -297 -3988
rect -215 3988 -169 4000
rect -215 -3988 -209 3988
rect -175 -3988 -169 3988
rect -215 -4000 -169 -3988
rect -87 3988 -41 4000
rect -87 -3988 -81 3988
rect -47 -3988 -41 3988
rect -87 -4000 -41 -3988
rect 41 3988 87 4000
rect 41 -3988 47 3988
rect 81 -3988 87 3988
rect 41 -4000 87 -3988
rect 169 3988 215 4000
rect 169 -3988 175 3988
rect 209 -3988 215 3988
rect 169 -4000 215 -3988
rect 297 3988 343 4000
rect 297 -3988 303 3988
rect 337 -3988 343 3988
rect 297 -4000 343 -3988
rect -287 -4047 -225 -4041
rect -287 -4081 -275 -4047
rect -237 -4081 -225 -4047
rect -287 -4087 -225 -4081
rect -159 -4047 -97 -4041
rect -159 -4081 -147 -4047
rect -109 -4081 -97 -4047
rect -159 -4087 -97 -4081
rect -31 -4047 31 -4041
rect -31 -4081 -19 -4047
rect 19 -4081 31 -4047
rect -31 -4087 31 -4081
rect 97 -4047 159 -4041
rect 97 -4081 109 -4047
rect 147 -4081 159 -4047
rect 97 -4087 159 -4081
rect 225 -4047 287 -4041
rect 225 -4081 237 -4047
rect 275 -4081 287 -4047
rect 225 -4087 287 -4081
<< properties >>
string FIXED_BBOX -434 -4166 434 4166
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 40.0 l 0.35 m 1 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
