magic
tech sky130A
magscale 1 2
timestamp 1695908076
<< nwell >>
rect -1812 -4219 1812 4219
<< pmoslvt >>
rect -1616 -4000 -1016 4000
rect -958 -4000 -358 4000
rect -300 -4000 300 4000
rect 358 -4000 958 4000
rect 1016 -4000 1616 4000
<< pdiff >>
rect -1674 3988 -1616 4000
rect -1674 -3988 -1662 3988
rect -1628 -3988 -1616 3988
rect -1674 -4000 -1616 -3988
rect -1016 3988 -958 4000
rect -1016 -3988 -1004 3988
rect -970 -3988 -958 3988
rect -1016 -4000 -958 -3988
rect -358 3988 -300 4000
rect -358 -3988 -346 3988
rect -312 -3988 -300 3988
rect -358 -4000 -300 -3988
rect 300 3988 358 4000
rect 300 -3988 312 3988
rect 346 -3988 358 3988
rect 300 -4000 358 -3988
rect 958 3988 1016 4000
rect 958 -3988 970 3988
rect 1004 -3988 1016 3988
rect 958 -4000 1016 -3988
rect 1616 3988 1674 4000
rect 1616 -3988 1628 3988
rect 1662 -3988 1674 3988
rect 1616 -4000 1674 -3988
<< pdiffc >>
rect -1662 -3988 -1628 3988
rect -1004 -3988 -970 3988
rect -346 -3988 -312 3988
rect 312 -3988 346 3988
rect 970 -3988 1004 3988
rect 1628 -3988 1662 3988
<< nsubdiff >>
rect -1776 4149 -1680 4183
rect 1680 4149 1776 4183
rect -1776 4087 -1742 4149
rect 1742 4087 1776 4149
rect -1776 -4149 -1742 -4087
rect 1742 -4149 1776 -4087
rect -1776 -4183 -1680 -4149
rect 1680 -4183 1776 -4149
<< nsubdiffcont >>
rect -1680 4149 1680 4183
rect -1776 -4087 -1742 4087
rect 1742 -4087 1776 4087
rect -1680 -4183 1680 -4149
<< poly >>
rect -1616 4081 -1016 4097
rect -1616 4047 -1600 4081
rect -1032 4047 -1016 4081
rect -1616 4000 -1016 4047
rect -958 4081 -358 4097
rect -958 4047 -942 4081
rect -374 4047 -358 4081
rect -958 4000 -358 4047
rect -300 4081 300 4097
rect -300 4047 -284 4081
rect 284 4047 300 4081
rect -300 4000 300 4047
rect 358 4081 958 4097
rect 358 4047 374 4081
rect 942 4047 958 4081
rect 358 4000 958 4047
rect 1016 4081 1616 4097
rect 1016 4047 1032 4081
rect 1600 4047 1616 4081
rect 1016 4000 1616 4047
rect -1616 -4047 -1016 -4000
rect -1616 -4081 -1600 -4047
rect -1032 -4081 -1016 -4047
rect -1616 -4097 -1016 -4081
rect -958 -4047 -358 -4000
rect -958 -4081 -942 -4047
rect -374 -4081 -358 -4047
rect -958 -4097 -358 -4081
rect -300 -4047 300 -4000
rect -300 -4081 -284 -4047
rect 284 -4081 300 -4047
rect -300 -4097 300 -4081
rect 358 -4047 958 -4000
rect 358 -4081 374 -4047
rect 942 -4081 958 -4047
rect 358 -4097 958 -4081
rect 1016 -4047 1616 -4000
rect 1016 -4081 1032 -4047
rect 1600 -4081 1616 -4047
rect 1016 -4097 1616 -4081
<< polycont >>
rect -1600 4047 -1032 4081
rect -942 4047 -374 4081
rect -284 4047 284 4081
rect 374 4047 942 4081
rect 1032 4047 1600 4081
rect -1600 -4081 -1032 -4047
rect -942 -4081 -374 -4047
rect -284 -4081 284 -4047
rect 374 -4081 942 -4047
rect 1032 -4081 1600 -4047
<< locali >>
rect -1776 4149 -1680 4183
rect 1680 4149 1776 4183
rect -1776 4087 -1742 4149
rect 1742 4087 1776 4149
rect -1616 4047 -1600 4081
rect -1032 4047 -1016 4081
rect -958 4047 -942 4081
rect -374 4047 -358 4081
rect -300 4047 -284 4081
rect 284 4047 300 4081
rect 358 4047 374 4081
rect 942 4047 958 4081
rect 1016 4047 1032 4081
rect 1600 4047 1616 4081
rect -1662 3988 -1628 4004
rect -1662 -4004 -1628 -3988
rect -1004 3988 -970 4004
rect -1004 -4004 -970 -3988
rect -346 3988 -312 4004
rect -346 -4004 -312 -3988
rect 312 3988 346 4004
rect 312 -4004 346 -3988
rect 970 3988 1004 4004
rect 970 -4004 1004 -3988
rect 1628 3988 1662 4004
rect 1628 -4004 1662 -3988
rect -1616 -4081 -1600 -4047
rect -1032 -4081 -1016 -4047
rect -958 -4081 -942 -4047
rect -374 -4081 -358 -4047
rect -300 -4081 -284 -4047
rect 284 -4081 300 -4047
rect 358 -4081 374 -4047
rect 942 -4081 958 -4047
rect 1016 -4081 1032 -4047
rect 1600 -4081 1616 -4047
rect -1776 -4149 -1742 -4087
rect 1742 -4149 1776 -4087
rect -1776 -4183 -1680 -4149
rect 1680 -4183 1776 -4149
<< viali >>
rect -1600 4047 -1032 4081
rect -942 4047 -374 4081
rect -284 4047 284 4081
rect 374 4047 942 4081
rect 1032 4047 1600 4081
rect -1662 -3988 -1628 3988
rect -1004 -3988 -970 3988
rect -346 -3988 -312 3988
rect 312 -3988 346 3988
rect 970 -3988 1004 3988
rect 1628 -3988 1662 3988
rect -1600 -4081 -1032 -4047
rect -942 -4081 -374 -4047
rect -284 -4081 284 -4047
rect 374 -4081 942 -4047
rect 1032 -4081 1600 -4047
<< metal1 >>
rect -1612 4081 -1020 4087
rect -1612 4047 -1600 4081
rect -1032 4047 -1020 4081
rect -1612 4041 -1020 4047
rect -954 4081 -362 4087
rect -954 4047 -942 4081
rect -374 4047 -362 4081
rect -954 4041 -362 4047
rect -296 4081 296 4087
rect -296 4047 -284 4081
rect 284 4047 296 4081
rect -296 4041 296 4047
rect 362 4081 954 4087
rect 362 4047 374 4081
rect 942 4047 954 4081
rect 362 4041 954 4047
rect 1020 4081 1612 4087
rect 1020 4047 1032 4081
rect 1600 4047 1612 4081
rect 1020 4041 1612 4047
rect -1668 3988 -1622 4000
rect -1668 -3988 -1662 3988
rect -1628 -3988 -1622 3988
rect -1668 -4000 -1622 -3988
rect -1010 3988 -964 4000
rect -1010 -3988 -1004 3988
rect -970 -3988 -964 3988
rect -1010 -4000 -964 -3988
rect -352 3988 -306 4000
rect -352 -3988 -346 3988
rect -312 -3988 -306 3988
rect -352 -4000 -306 -3988
rect 306 3988 352 4000
rect 306 -3988 312 3988
rect 346 -3988 352 3988
rect 306 -4000 352 -3988
rect 964 3988 1010 4000
rect 964 -3988 970 3988
rect 1004 -3988 1010 3988
rect 964 -4000 1010 -3988
rect 1622 3988 1668 4000
rect 1622 -3988 1628 3988
rect 1662 -3988 1668 3988
rect 1622 -4000 1668 -3988
rect -1612 -4047 -1020 -4041
rect -1612 -4081 -1600 -4047
rect -1032 -4081 -1020 -4047
rect -1612 -4087 -1020 -4081
rect -954 -4047 -362 -4041
rect -954 -4081 -942 -4047
rect -374 -4081 -362 -4047
rect -954 -4087 -362 -4081
rect -296 -4047 296 -4041
rect -296 -4081 -284 -4047
rect 284 -4081 296 -4047
rect -296 -4087 296 -4081
rect 362 -4047 954 -4041
rect 362 -4081 374 -4047
rect 942 -4081 954 -4047
rect 362 -4087 954 -4081
rect 1020 -4047 1612 -4041
rect 1020 -4081 1032 -4047
rect 1600 -4081 1612 -4047
rect 1020 -4087 1612 -4081
<< labels >>
rlabel poly -300 4000 300 4047 1 G
rlabel locali -1662 3988 -1628 4004 1 D
rlabel locali 1628 3988 1662 4004 1 S
rlabel nsubdiffcont -1680 4149 1680 4183 1 B
<< properties >>
string FIXED_BBOX -1759 -4166 1759 4166
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 40.0 l 3.0 m 1 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
