magic
tech sky130A
timestamp 1695377223
<< metal1 >>
rect 14251 11814 25323 13960
rect 12183 9432 12283 9442
rect 12183 9353 12192 9432
rect 12272 9353 12283 9432
rect 12183 9342 12283 9353
rect 12789 9434 12910 9460
rect 12789 9341 12804 9434
rect 12886 9341 12910 9434
rect 11876 4931 11994 4942
rect 11876 4903 12576 4931
rect 11876 4805 12460 4903
rect 12561 4805 12576 4903
rect 11876 4773 12576 4805
rect 11876 -2302 11994 4773
rect 12789 359 12910 9341
rect 12256 342 12356 355
rect 12256 266 12269 342
rect 12340 266 12356 342
rect 12256 255 12356 266
rect 12789 283 12806 359
rect 12883 283 12910 359
rect 12789 -2315 12910 283
rect 19232 -1874 20091 11814
rect 26202 9402 26453 9432
rect 26202 9323 26294 9402
rect 26367 9323 26453 9402
rect 26202 357 26453 9323
rect 27043 9396 27143 9408
rect 27043 9321 27053 9396
rect 27130 9321 27143 9396
rect 27043 9308 27143 9321
rect 26202 274 26292 357
rect 26374 274 26453 357
rect 11898 -3347 11980 -2793
rect 12793 -3051 12875 -2794
rect 26202 -3051 26453 274
rect 26663 4885 26886 4914
rect 26663 4805 26723 4885
rect 26806 4805 26886 4885
rect 12793 -3203 26461 -3051
rect 12793 -3346 12875 -3203
rect 11894 -3506 11983 -3347
rect 12785 -3446 12885 -3346
rect 26663 -3506 26886 4805
rect 27098 4895 27198 4902
rect 27098 4809 27104 4895
rect 27190 4809 27198 4895
rect 27098 4802 27198 4809
rect 27114 368 27214 380
rect 27114 296 27125 368
rect 27201 296 27214 368
rect 27114 280 27214 296
rect 11885 -3625 26888 -3506
<< via1 >>
rect 12192 9353 12272 9432
rect 12804 9341 12886 9434
rect 12460 4805 12561 4903
rect 12269 266 12340 342
rect 12806 283 12883 359
rect 26294 9323 26367 9402
rect 27053 9321 27130 9396
rect 26292 274 26374 357
rect 26723 4805 26806 4885
rect 27104 4809 27190 4895
rect 27125 296 27201 368
<< metal2 >>
rect 12158 9450 12316 9461
rect 12158 9324 12174 9450
rect 12303 9324 12316 9450
rect 12158 9313 12316 9324
rect 12790 9434 12907 9451
rect 12790 9341 12804 9434
rect 12886 9341 12907 9434
rect 12790 9318 12907 9341
rect 17281 7183 22125 11438
rect 27006 9425 27173 9444
rect 26271 9402 26384 9425
rect 26271 9323 26294 9402
rect 26367 9323 26384 9402
rect 26271 9302 26384 9323
rect 27006 9296 27017 9425
rect 27154 9296 27173 9425
rect 27006 9281 27173 9296
rect 21117 6597 22076 7183
rect 27055 4925 27241 4944
rect 12448 4903 12570 4916
rect 12448 4805 12460 4903
rect 12561 4805 12570 4903
rect 26700 4885 26830 4908
rect 12448 4783 12570 4805
rect 26700 4805 26723 4885
rect 26806 4805 26830 4885
rect 26700 4782 26830 4805
rect 27055 4782 27078 4925
rect 27217 4782 27241 4925
rect 27055 4767 27241 4782
rect 17183 2445 18138 3127
rect 12245 358 12369 374
rect 12245 248 12253 358
rect 12361 248 12369 358
rect 12788 359 12906 379
rect 12788 283 12806 359
rect 12883 283 12906 359
rect 12788 264 12906 283
rect 12245 230 12369 248
rect 17183 -1701 22027 2445
rect 27085 398 27241 422
rect 26272 357 26400 375
rect 26272 274 26292 357
rect 26374 274 26400 357
rect 26272 254 26400 274
rect 27085 271 27093 398
rect 27232 271 27241 398
rect 27085 235 27241 271
rect 17271 -1810 22027 -1701
<< via2 >>
rect 12174 9432 12303 9450
rect 12174 9353 12192 9432
rect 12192 9353 12272 9432
rect 12272 9353 12303 9432
rect 12174 9324 12303 9353
rect 12804 9341 12886 9434
rect 14592 9045 14790 9238
rect 26294 9323 26367 9402
rect 27017 9396 27154 9425
rect 27017 9321 27053 9396
rect 27053 9321 27130 9396
rect 27130 9321 27154 9396
rect 27017 9296 27154 9321
rect 24573 9017 24772 9209
rect 12460 4805 12561 4903
rect 15483 4823 15544 4882
rect 26723 4805 26806 4885
rect 27078 4895 27217 4925
rect 27078 4809 27104 4895
rect 27104 4809 27190 4895
rect 27190 4809 27217 4895
rect 27078 4782 27217 4809
rect 14650 4542 14767 4674
rect 21574 4499 21768 4688
rect 12253 342 12361 358
rect 12253 266 12269 342
rect 12269 266 12340 342
rect 12340 266 12361 342
rect 12253 248 12361 266
rect 12806 283 12883 359
rect 14538 -42 14784 196
rect 26292 274 26374 357
rect 27093 368 27232 398
rect 27093 296 27125 368
rect 27125 296 27201 368
rect 27201 296 27232 368
rect 27093 271 27232 296
rect 24553 -43 24784 186
<< metal3 >>
rect 12073 9512 12393 9557
rect 12073 9251 12100 9512
rect 12364 9251 12393 9512
rect 26945 9467 27247 9489
rect 12783 9434 15588 9453
rect 12783 9341 12804 9434
rect 12886 9341 15588 9434
rect 12783 9312 15588 9341
rect 23775 9402 26464 9429
rect 23775 9323 26294 9402
rect 26367 9323 26464 9402
rect 23775 9288 26464 9323
rect 12073 9200 12393 9251
rect 14553 9238 14830 9267
rect 26945 9253 26971 9467
rect 27225 9253 27247 9467
rect 14553 9045 14592 9238
rect 14790 9045 14830 9238
rect 14553 8979 14830 9045
rect 24531 9209 24816 9243
rect 26945 9229 27247 9253
rect 24531 9017 24573 9209
rect 24772 9017 24816 9209
rect 24531 8983 24816 9017
rect 26993 4961 27296 4978
rect 12443 4908 15569 4921
rect 12443 4903 15573 4908
rect 12443 4805 12460 4903
rect 12561 4882 15573 4903
rect 12561 4823 15483 4882
rect 15544 4823 15573 4882
rect 12561 4805 15573 4823
rect 12443 4797 15573 4805
rect 23747 4885 26873 4911
rect 23747 4805 26723 4885
rect 26806 4805 26873 4885
rect 12443 4780 15569 4797
rect 23747 4770 26873 4805
rect 26993 4746 27017 4961
rect 27274 4746 27296 4961
rect 26993 4732 27296 4746
rect 14616 4674 14797 4708
rect 14616 4542 14650 4674
rect 14767 4542 14797 4674
rect 14616 4515 14797 4542
rect 21542 4688 21800 4721
rect 21542 4499 21574 4688
rect 21768 4499 21800 4688
rect 21542 4468 21800 4499
rect 27026 457 27299 511
rect 12171 400 12433 437
rect 12171 216 12212 400
rect 12397 216 12433 400
rect 12774 359 15521 393
rect 12774 283 12806 359
rect 12883 283 15521 359
rect 12774 252 15521 283
rect 23750 357 26464 386
rect 23750 274 26292 357
rect 26374 274 26464 357
rect 23750 245 26464 274
rect 12171 186 12433 216
rect 14508 196 14809 220
rect 27026 209 27066 457
rect 27267 209 27299 457
rect 14508 -42 14538 196
rect 14784 -42 14809 196
rect 14508 -62 14809 -42
rect 24521 186 24818 201
rect 24521 -43 24553 186
rect 24784 -43 24818 186
rect 27026 162 27299 209
rect 24521 -65 24818 -43
<< via3 >>
rect 12100 9450 12364 9512
rect 12100 9324 12174 9450
rect 12174 9324 12303 9450
rect 12303 9324 12364 9450
rect 12100 9251 12364 9324
rect 26971 9425 27225 9467
rect 26971 9296 27017 9425
rect 27017 9296 27154 9425
rect 27154 9296 27225 9425
rect 26971 9253 27225 9296
rect 14592 9045 14790 9238
rect 24573 9017 24772 9209
rect 27017 4925 27274 4961
rect 27017 4782 27078 4925
rect 27078 4782 27217 4925
rect 27217 4782 27274 4925
rect 27017 4746 27274 4782
rect 14650 4542 14767 4674
rect 21574 4499 21768 4688
rect 12212 358 12397 400
rect 12212 248 12253 358
rect 12253 248 12361 358
rect 12361 248 12397 358
rect 12212 216 12397 248
rect 27066 398 27267 457
rect 27066 271 27093 398
rect 27093 271 27232 398
rect 27232 271 27267 398
rect 27066 209 27267 271
rect 14538 -42 14784 196
rect 24553 -43 24784 186
<< metal4 >>
rect 11877 9512 14922 10126
rect 11877 9251 12100 9512
rect 12364 9251 14922 9512
rect 11877 9238 14922 9251
rect 11877 9045 14592 9238
rect 14790 9045 14922 9238
rect 11877 8575 14922 9045
rect 24476 9467 27521 10108
rect 24476 9253 26971 9467
rect 27225 9253 27521 9467
rect 24476 9209 27521 9253
rect 24476 9017 24573 9209
rect 24772 9017 27521 9209
rect 24476 8557 27521 9017
rect 23209 6450 27397 6473
rect 14256 4961 27397 6450
rect 14256 4746 27017 4961
rect 27274 4746 27397 4961
rect 14256 4688 27397 4746
rect 14256 4674 21574 4688
rect 14256 4542 14650 4674
rect 14767 4542 21574 4674
rect 14256 4499 21574 4542
rect 21768 4499 27397 4688
rect 14256 3257 27397 4499
rect 14256 3230 25097 3257
rect 11896 400 14941 1066
rect 11896 216 12212 400
rect 12397 216 14941 400
rect 11896 196 14941 216
rect 11896 -42 14538 196
rect 14784 -42 14941 196
rect 11896 -485 14941 -42
rect 24423 457 27468 1060
rect 24423 209 27066 457
rect 27267 209 27468 457
rect 24423 186 27468 209
rect 24423 -43 24553 186
rect 24784 -43 27468 186
rect 24423 -491 27468 -43
use not  x1
timestamp 1695377178
transform 0 1 11852 1 0 -3137
box 238 -289 934 495
use not  x2
timestamp 1695377178
transform 0 -1 12929 1 0 -3139
box 238 -289 934 495
use switch  x3
timestamp 1695377223
transform 0 1 13842 1 0 2681
box -57 -475 4321 5709
use switch  x4
timestamp 1695377223
transform 0 -1 25493 1 0 -1857
box -57 -475 4321 5709
use switch  x5
timestamp 1695377223
transform 0 1 13793 1 0 -1857
box -57 -475 4321 5709
use switch  x6
timestamp 1695377223
transform 0 -1 25482 1 0 2663
box -57 -475 4321 5709
use switch  x7
timestamp 1695377223
transform 0 -1 25519 1 0 7181
box -57 -475 4321 5709
use switch  x8
timestamp 1695377223
transform 0 1 13868 1 0 7205
box -57 -475 4321 5709
<< labels >>
flabel metal1 12785 -3446 12885 -3346 0 FreeSans 128 0 0 0 SEL0
port 0 nsew
flabel metal1 11886 -3609 11986 -3509 0 FreeSans 128 0 0 0 SEL1
port 1 nsew
flabel metal1 12256 255 12356 355 0 FreeSans 128 0 0 0 IN0
port 2 nsew
flabel metal1 27114 280 27214 380 0 FreeSans 128 0 0 0 IN1
port 3 nsew
flabel metal1 12183 9342 12283 9442 0 FreeSans 128 0 0 0 IN2
port 5 nsew
flabel metal1 27043 9308 27143 9408 0 FreeSans 128 0 0 0 IN3
port 6 nsew
flabel metal1 27098 4802 27198 4902 0 FreeSans 128 0 0 0 OUT
port 4 nsew
rlabel metal1 14251 11814 25323 13960 1 VDD
<< end >>
