magic
tech sky130A
timestamp 1695432261
<< metal1 >>
rect 9308 15285 9872 15369
rect 2597 15169 2704 15195
rect 2597 15063 2621 15169
rect 2673 15063 2704 15169
rect 2201 8252 2335 8281
rect 2201 8193 2237 8252
rect 2298 8193 2335 8252
rect 2201 6239 2335 8193
rect 2597 6273 2704 15063
rect 9308 15108 9438 15285
rect 9748 15108 9872 15285
rect 3208 13018 3308 13030
rect 3208 12938 3214 13018
rect 3297 12938 3308 13018
rect 3208 12930 3308 12938
rect 2962 6869 3071 12775
rect 3232 8489 3332 8497
rect 3232 8403 3238 8489
rect 3324 8403 3332 8489
rect 3232 8397 3332 8403
rect 2957 6239 3054 6391
rect 2201 6232 3054 6239
rect 2201 6134 3057 6232
rect 2957 6132 3057 6134
rect 3272 5872 3377 6397
rect 3272 5766 3295 5872
rect 3347 5766 3377 5872
rect 3272 5740 3377 5766
rect 3707 5869 4268 11002
rect 9308 6110 9872 15108
rect 10261 10497 10361 10506
rect 10261 10416 10269 10497
rect 10353 10416 10361 10497
rect 10261 10406 10361 10416
rect 3707 5631 3821 5869
rect 4160 5631 4268 5869
rect 3707 5588 4268 5631
<< via1 >>
rect 2621 15063 2673 15169
rect 2237 8193 2298 8252
rect 9438 15108 9748 15285
rect 3214 12938 3297 13018
rect 3238 8403 3324 8489
rect 3295 5766 3347 5872
rect 10269 10416 10353 10497
rect 3821 5631 4160 5869
<< metal2 >>
rect 2120 15285 10436 16746
rect 2120 15169 9438 15285
rect 2120 15063 2621 15169
rect 2673 15108 9438 15169
rect 9748 15108 10436 15285
rect 2673 15063 10436 15108
rect 2120 15037 10436 15063
rect 3057 13018 5270 14366
rect 3057 12938 3214 13018
rect 3297 12938 5270 13018
rect 3057 12816 5270 12938
rect 2947 12742 3094 12769
rect 2947 12682 2988 12742
rect 3045 12682 3094 12742
rect 2947 12659 3094 12682
rect 5773 12758 5891 12775
rect 5773 12679 5790 12758
rect 5880 12679 5891 12758
rect 5773 12667 5891 12679
rect 7877 10497 10395 14832
rect 7877 10416 10269 10497
rect 10353 10416 10395 10497
rect 3065 8489 5278 9868
rect 3065 8403 3238 8489
rect 3324 8403 5278 8489
rect 3065 8318 5278 8403
rect 2192 8252 2351 8275
rect 2192 8193 2237 8252
rect 2298 8193 2351 8252
rect 2192 8165 2351 8193
rect 5789 8245 5889 8269
rect 5789 8179 5805 8245
rect 5876 8179 5889 8245
rect 5789 8144 5889 8179
rect 7877 6134 10395 10416
rect 2100 5872 10416 5920
rect 2100 5766 3295 5872
rect 3347 5869 10416 5872
rect 3347 5766 3821 5869
rect 2100 5631 3821 5766
rect 4160 5631 10416 5869
rect 2100 4211 10416 5631
<< via2 >>
rect 2988 12682 3045 12742
rect 5790 12679 5880 12758
rect 2237 8193 2298 8252
rect 5805 8179 5876 8245
<< metal3 >>
rect 2947 12758 5902 12781
rect 2947 12742 5790 12758
rect 2947 12682 2988 12742
rect 3045 12682 5790 12742
rect 2947 12679 5790 12682
rect 5880 12679 5902 12758
rect 2947 12656 5902 12679
rect 5775 8279 5905 8283
rect 2180 8252 5905 8279
rect 2180 8193 2237 8252
rect 2298 8245 5905 8252
rect 2298 8193 5805 8245
rect 2180 8179 5805 8193
rect 5876 8179 5905 8245
rect 2180 8154 5905 8179
rect 5775 8141 5905 8154
use not  x1
timestamp 1695395215
transform 0 -1 3093 1 0 6035
box 238 -289 934 495
use switch  x5
timestamp 1695432073
transform 0 1 4161 -1 0 14889
box -57 -475 4321 5709
use switch  x6
timestamp 1695432073
transform 0 1 4170 -1 0 10392
box -57 -475 4321 5709
<< labels >>
flabel metal1 2957 6132 3057 6232 0 FreeSans 128 0 0 0 SEL0
port 0 nsew
flabel metal1 3208 12930 3308 13030 0 FreeSans 128 0 0 0 IN0
port 3 nsew
flabel metal1 3232 8397 3332 8497 0 FreeSans 128 0 0 0 IN1
port 1 nsew
flabel metal1 10261 10406 10361 10506 0 FreeSans 128 0 0 0 OUT
port 2 nsew
rlabel metal2 2100 4211 10416 5920 1 GROUND
port 4 nsew
rlabel metal2 2120 15037 10436 16746 1 VDD
port 5 nsew
rlabel metal2 5244 4612 6614 5395 1 GROUND
rlabel metal2 5494 15495 6864 16278 1 VDD
<< end >>
