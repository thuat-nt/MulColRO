magic
tech sky130A
magscale 1 2
timestamp 1695365668
<< error_p >>
rect 18727 3662 18762 3696
rect 18728 3643 18762 3662
rect 17150 2383 17165 3249
rect 17184 2383 17218 3303
rect 17184 2349 17199 2383
rect 18747 2330 18762 3643
rect 18781 3609 18816 3643
rect 18781 2330 18815 3609
rect 26150 3503 26185 3537
rect 28459 3520 28493 3538
rect 26151 3484 26185 3503
rect 18781 2296 18796 2330
rect 26170 2171 26185 3484
rect 26204 3450 26239 3484
rect 26204 2171 26238 3450
rect 26204 2137 26219 2171
rect 28423 2118 28493 3520
rect 31977 3360 32011 3414
rect 28423 2082 28476 2118
rect 31996 2065 32011 3360
rect 32030 3326 32065 3360
rect 32915 3326 32950 3360
rect 32030 2065 32064 3326
rect 32916 3307 32950 3326
rect 32030 2031 32045 2065
rect 32935 2012 32950 3307
rect 32969 3273 33004 3307
rect 32969 2012 33003 3273
rect 32969 1978 32984 2012
rect 33874 1959 33889 3307
rect 33908 1959 33942 3361
rect 33908 1925 33923 1959
<< error_s >>
rect 34793 3820 34828 3854
rect 34794 3801 34828 3820
rect 34813 1906 34828 3801
rect 34847 3767 34882 3801
rect 34847 1906 34881 3767
rect 43726 2446 43728 3848
rect 43829 1970 44498 10385
rect 44594 8508 44600 9860
rect 51752 2446 51754 3848
rect 51855 1970 52524 10385
rect 52620 8508 52626 9860
rect 59778 2446 59780 3848
rect 59881 1970 60550 10385
rect 60646 8508 60652 9860
rect 34847 1872 34862 1906
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
use opamp  x1
timestamp 1695307921
transform 1 0 12744 0 1 1800
box 0 -1200 23059 8696
use switch  x2
timestamp 1695359377
transform 1 0 35856 0 1 1400
box -114 -950 8642 11418
use switch  x3
timestamp 1695359377
transform 1 0 43882 0 1 1400
box -114 -950 8642 11418
use switch  x4
timestamp 1695359377
transform 1 0 51908 0 1 1400
box -114 -950 8642 11418
use switch  x5
timestamp 1695359377
transform 1 0 59934 0 1 1400
box -114 -950 8642 11418
use sky130_fd_pr__cap_mim_m3_1_3HBNLG  XC1
timestamp 1695196838
transform 1 0 3186 0 1 3640
box -3186 -3040 3186 3040
use sky130_fd_pr__cap_mim_m3_1_3HBNLG  XC2
timestamp 1695196838
transform 1 0 9558 0 1 3640
box -3186 -3040 3186 3040
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 opbias
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 cdsin
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 cdsout
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 sw1
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 sw2
port 4 nsew
<< end >>
