magic
tech sky130A
magscale 1 2
timestamp 1695365668
<< error_p >>
rect 12355 3662 12390 3696
rect 12356 3643 12390 3662
rect 10778 2383 10793 3249
rect 10812 2383 10846 3303
rect 10812 2349 10827 2383
rect 12375 2330 12390 3643
rect 12409 3609 12444 3643
rect 12409 2330 12443 3609
rect 19778 3503 19813 3537
rect 22087 3520 22121 3538
rect 19779 3484 19813 3503
rect 12409 2296 12424 2330
rect 19798 2171 19813 3484
rect 19832 3450 19867 3484
rect 19832 2171 19866 3450
rect 19832 2137 19847 2171
rect 22051 2118 22121 3520
rect 25605 3360 25639 3414
rect 22051 2082 22104 2118
rect 25624 2065 25639 3360
rect 25658 3326 25693 3360
rect 26543 3326 26578 3360
rect 25658 2065 25692 3326
rect 26544 3307 26578 3326
rect 25658 2031 25673 2065
rect 26563 2012 26578 3307
rect 26597 3273 26632 3307
rect 26597 2012 26631 3273
rect 26597 1978 26612 2012
rect 27502 1959 27517 3307
rect 27536 1959 27570 3361
rect 27536 1925 27551 1959
<< error_s >>
rect 28421 3820 28456 3854
rect 28422 3801 28456 3820
rect 28441 1906 28456 3801
rect 28475 3767 28510 3801
rect 28475 1906 28509 3767
rect 37354 2446 37356 3848
rect 37457 1970 38126 10385
rect 38222 8508 38228 9860
rect 45380 2446 45382 3848
rect 45483 1970 46152 10385
rect 46248 8508 46254 9860
rect 54004 2006 54142 2024
rect 54038 1972 54176 1990
rect 28475 1872 28490 1906
rect 54046 1046 54066 1302
rect 54074 1074 54122 1274
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
use opamp  x1
timestamp 1695307921
transform 1 0 6372 0 1 1800
box 0 -1200 23059 8696
use switch  x2
timestamp 1695359377
transform 1 0 29484 0 1 1400
box -114 -950 8642 11418
use switch  x3
timestamp 1695359377
transform 1 0 37510 0 1 1400
box -114 -950 8642 11418
use switch  x4
timestamp 1695359377
transform 1 0 45536 0 1 1400
box -114 -950 8642 11418
use not  x5
timestamp 1695355038
transform 1 0 53562 0 1 1000
box 476 -578 1868 990
use not  x6
timestamp 1695355038
transform 1 0 54393 0 1 1000
box 476 -578 1868 990
use not  x7
timestamp 1695355038
transform 1 0 55224 0 1 1000
box 476 -578 1868 990
use sky130_fd_pr__cap_mim_m3_1_3HBNLG  XC1
timestamp 1695196838
transform 1 0 3186 0 1 3640
box -3186 -3040 3186 3040
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 sw1
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 opbias
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 shin
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 shout
port 3 nsew
<< end >>
