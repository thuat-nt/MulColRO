magic
tech sky130A
magscale 1 2
timestamp 1698053393
<< nwell >>
rect -487 -4219 487 4219
<< pmoslvt >>
rect -291 -4000 -221 4000
rect -163 -4000 -93 4000
rect -35 -4000 35 4000
rect 93 -4000 163 4000
rect 221 -4000 291 4000
<< pdiff >>
rect -349 3988 -291 4000
rect -349 -3988 -337 3988
rect -303 -3988 -291 3988
rect -349 -4000 -291 -3988
rect -221 3988 -163 4000
rect -221 -3988 -209 3988
rect -175 -3988 -163 3988
rect -221 -4000 -163 -3988
rect -93 3988 -35 4000
rect -93 -3988 -81 3988
rect -47 -3988 -35 3988
rect -93 -4000 -35 -3988
rect 35 3988 93 4000
rect 35 -3988 47 3988
rect 81 -3988 93 3988
rect 35 -4000 93 -3988
rect 163 3988 221 4000
rect 163 -3988 175 3988
rect 209 -3988 221 3988
rect 163 -4000 221 -3988
rect 291 3988 349 4000
rect 291 -3988 303 3988
rect 337 -3988 349 3988
rect 291 -4000 349 -3988
<< pdiffc >>
rect -337 -3988 -303 3988
rect -209 -3988 -175 3988
rect -81 -3988 -47 3988
rect 47 -3988 81 3988
rect 175 -3988 209 3988
rect 303 -3988 337 3988
<< nsubdiff >>
rect -451 4149 -355 4183
rect 355 4149 451 4183
rect -451 4087 -417 4149
rect 417 4087 451 4149
rect -451 -4149 -417 -4087
rect 417 -4149 451 -4087
rect -451 -4183 -355 -4149
rect 355 -4183 451 -4149
<< nsubdiffcont >>
rect -355 4149 355 4183
rect -451 -4087 -417 4087
rect 417 -4087 451 4087
rect -355 -4183 355 -4149
<< poly >>
rect -291 4081 -221 4097
rect -291 4047 -275 4081
rect -237 4047 -221 4081
rect -291 4000 -221 4047
rect -163 4081 -93 4097
rect -163 4047 -147 4081
rect -109 4047 -93 4081
rect -163 4000 -93 4047
rect -35 4081 35 4097
rect -35 4047 -19 4081
rect 19 4047 35 4081
rect -35 4000 35 4047
rect 93 4081 163 4097
rect 93 4047 109 4081
rect 147 4047 163 4081
rect 93 4000 163 4047
rect 221 4081 291 4097
rect 221 4047 237 4081
rect 275 4047 291 4081
rect 221 4000 291 4047
rect -291 -4047 -221 -4000
rect -291 -4081 -275 -4047
rect -237 -4081 -221 -4047
rect -291 -4097 -221 -4081
rect -163 -4047 -93 -4000
rect -163 -4081 -147 -4047
rect -109 -4081 -93 -4047
rect -163 -4097 -93 -4081
rect -35 -4048 35 -4000
rect -35 -4082 -16 -4048
rect 18 -4082 35 -4048
rect -35 -4097 35 -4082
rect 93 -4047 163 -4000
rect 93 -4081 109 -4047
rect 147 -4081 163 -4047
rect 93 -4097 163 -4081
rect 221 -4047 291 -4000
rect 221 -4081 237 -4047
rect 275 -4081 291 -4047
rect 221 -4097 291 -4081
<< polycont >>
rect -275 4047 -237 4081
rect -147 4047 -109 4081
rect -19 4047 19 4081
rect 109 4047 147 4081
rect 237 4047 275 4081
rect -275 -4081 -237 -4047
rect -147 -4081 -109 -4047
rect -16 -4082 18 -4048
rect 109 -4081 147 -4047
rect 237 -4081 275 -4047
<< locali >>
rect -451 4149 -355 4183
rect 355 4149 451 4183
rect -451 4087 -417 4149
rect 417 4087 451 4149
rect -36 4081 34 4082
rect -291 4047 -275 4081
rect -237 4047 -221 4081
rect -163 4047 -147 4081
rect -109 4047 -93 4081
rect -36 4047 -19 4081
rect 19 4047 35 4081
rect 93 4047 109 4081
rect 147 4047 163 4081
rect 221 4047 237 4081
rect 275 4047 291 4081
rect -36 4044 34 4047
rect -337 3988 -303 4004
rect -337 -4004 -303 -3988
rect -209 3988 -175 4004
rect -209 -4004 -175 -3988
rect -81 3988 -47 4004
rect -81 -4004 -47 -3988
rect 47 3988 81 4004
rect 47 -4004 81 -3988
rect 175 3988 209 4004
rect 175 -4004 209 -3988
rect 303 3988 337 4004
rect 303 -4004 337 -3988
rect -291 -4081 -275 -4047
rect -237 -4081 -221 -4047
rect -163 -4081 -147 -4047
rect -109 -4081 -93 -4047
rect -34 -4082 -16 -4048
rect 18 -4082 36 -4048
rect 93 -4081 109 -4047
rect 147 -4081 163 -4047
rect 221 -4081 237 -4047
rect 275 -4081 291 -4047
rect -34 -4084 36 -4082
rect -451 -4149 -417 -4087
rect 417 -4149 451 -4087
rect -451 -4183 -355 -4149
rect 355 -4183 451 -4149
<< viali >>
rect -275 4047 -237 4081
rect -147 4047 -109 4081
rect -19 4047 19 4081
rect 109 4047 147 4081
rect 237 4047 275 4081
rect -337 -3988 -303 3988
rect -209 -3988 -175 3988
rect -81 -3988 -47 3988
rect 47 -3988 81 3988
rect 175 -3988 209 3988
rect 303 -3988 337 3988
rect -275 -4081 -237 -4047
rect -147 -4081 -109 -4047
rect -16 -4082 18 -4048
rect 109 -4081 147 -4047
rect 237 -4081 275 -4047
<< metal1 >>
rect -290 4081 290 4096
rect -290 4047 -275 4081
rect -237 4047 -147 4081
rect -109 4047 -19 4081
rect 19 4047 109 4081
rect 147 4047 237 4081
rect 275 4047 290 4081
rect -290 4032 290 4047
rect -380 3988 -258 4002
rect -380 3780 -337 3988
rect -303 3780 -258 3988
rect -380 3464 -360 3780
rect -282 3464 -258 3780
rect -380 3302 -337 3464
rect -343 -3988 -337 3302
rect -303 3302 -258 3464
rect -215 3988 -169 4000
rect -303 -3988 -297 3302
rect -215 -3202 -209 3988
rect -260 -3388 -209 -3202
rect -175 -3202 -169 3988
rect -124 3988 0 4000
rect -124 3756 -81 3988
rect -47 3756 0 3988
rect -124 3442 -106 3756
rect -20 3442 0 3756
rect -124 3300 -81 3442
rect -175 -3388 -126 -3202
rect -260 -3884 -234 -3388
rect -148 -3884 -126 -3388
rect -260 -3968 -209 -3884
rect -343 -4000 -297 -3988
rect -215 -3988 -209 -3968
rect -175 -3968 -126 -3884
rect -175 -3988 -169 -3968
rect -215 -4000 -169 -3988
rect -87 -3988 -81 3300
rect -47 3300 0 3442
rect 41 3988 87 4000
rect -47 -3988 -41 3300
rect 41 -3198 47 3988
rect 2 -3374 47 -3198
rect 81 -3198 87 3988
rect 130 3988 254 4002
rect 130 3758 175 3988
rect 209 3758 254 3988
rect 130 3444 152 3758
rect 238 3444 254 3758
rect 130 3302 175 3444
rect 81 -3374 136 -3198
rect 2 -3870 26 -3374
rect 112 -3870 136 -3374
rect 2 -3964 47 -3870
rect -87 -4000 -41 -3988
rect 41 -3988 47 -3964
rect 81 -3964 136 -3870
rect 81 -3988 87 -3964
rect 41 -4000 87 -3988
rect 169 -3988 175 3302
rect 209 3302 254 3444
rect 297 3988 343 4000
rect 209 -3988 215 3302
rect 297 -3196 303 3988
rect 256 -3374 303 -3196
rect 337 -3196 343 3988
rect 337 -3374 390 -3196
rect 256 -3870 278 -3374
rect 364 -3870 390 -3374
rect 256 -3962 303 -3870
rect 169 -4000 215 -3988
rect 297 -3988 303 -3962
rect 337 -3962 390 -3870
rect 337 -3988 343 -3962
rect 297 -4000 343 -3988
rect -292 -4047 294 -4036
rect -292 -4081 -275 -4047
rect -237 -4081 -147 -4047
rect -109 -4048 109 -4047
rect -109 -4081 -16 -4048
rect -292 -4082 -16 -4081
rect 18 -4081 109 -4048
rect 147 -4081 237 -4047
rect 275 -4081 294 -4047
rect 18 -4082 294 -4081
rect -292 -4098 294 -4082
rect -40 -4100 42 -4098
<< via1 >>
rect -360 3464 -337 3780
rect -337 3464 -303 3780
rect -303 3464 -282 3780
rect -106 3442 -81 3756
rect -81 3442 -47 3756
rect -47 3442 -20 3756
rect -234 -3884 -209 -3388
rect -209 -3884 -175 -3388
rect -175 -3884 -148 -3388
rect 152 3444 175 3758
rect 175 3444 209 3758
rect 209 3444 238 3758
rect 26 -3870 47 -3374
rect 47 -3870 81 -3374
rect 81 -3870 112 -3374
rect 278 -3870 303 -3374
rect 303 -3870 337 -3374
rect 337 -3870 364 -3374
<< metal2 >>
rect -382 3780 -258 3826
rect -382 3464 -360 3780
rect -282 3464 -258 3780
rect -382 3412 -258 3464
rect -124 3756 0 3810
rect -124 3442 -106 3756
rect -20 3442 0 3756
rect -124 3396 0 3442
rect 132 3758 256 3814
rect 132 3444 152 3758
rect 238 3444 256 3758
rect 132 3400 256 3444
rect -250 -3388 -130 -3344
rect -250 -3884 -234 -3388
rect -148 -3884 -130 -3388
rect -250 -3910 -130 -3884
rect 12 -3374 132 -3340
rect 12 -3870 26 -3374
rect 112 -3870 132 -3374
rect 12 -3906 132 -3870
rect 262 -3374 382 -3328
rect 262 -3870 278 -3374
rect 364 -3870 382 -3374
rect 262 -3894 382 -3870
<< properties >>
string FIXED_BBOX -434 -4166 434 4166
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 40.0 l 0.35 m 1 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
