magic
tech sky130A
magscale 1 2
timestamp 1695908076
<< locali >>
rect 878 9600 11320 10390
rect 878 9528 2036 9600
rect 2212 9528 11320 9600
rect 878 9386 11320 9528
rect 3434 6974 11220 7188
rect 1020 6772 11220 6974
rect 1020 6760 3518 6772
rect 896 6164 1024 6192
rect 11226 6164 11276 6196
rect 896 6130 11276 6164
rect 896 6054 11238 6130
rect 896 5826 9242 6054
rect 9736 5826 11238 6054
rect 896 5142 11238 5826
rect 896 5130 1024 5142
<< viali >>
rect 2036 9528 2212 9600
rect 9242 5826 9736 6054
<< metal1 >>
rect 1994 9600 2242 9612
rect 1994 9524 2032 9600
rect 2218 9524 2242 9600
rect 1994 9518 2242 9524
rect 644 8318 844 8376
rect 644 8226 670 8318
rect 826 8226 844 8318
rect 644 8176 844 8226
rect 1368 8336 2862 9366
rect 3078 9130 3202 9194
rect 3078 8828 3134 9130
rect 3194 8828 3202 9130
rect 3078 8776 3202 8828
rect 7022 8508 7222 8584
rect 7022 8452 7070 8508
rect 7168 8452 7222 8508
rect 7022 8384 7222 8452
rect 1368 8222 1922 8336
rect 2336 8222 2862 8336
rect 1062 7670 1158 7736
rect 1062 7362 1078 7670
rect 1134 7362 1158 7670
rect 1062 7324 1158 7362
rect 1368 7170 2862 8222
rect 4662 8044 4748 8060
rect 4662 7984 4672 8044
rect 4736 7984 4748 8044
rect 4662 7968 4748 7984
rect 4668 7966 4732 7968
rect 5810 7732 8316 8190
rect 5810 7676 6764 7732
rect 7376 7676 8316 7732
rect 5810 7210 8316 7676
rect 9708 7424 9798 7436
rect 9708 7358 9730 7424
rect 9784 7358 9798 7424
rect 9708 7346 9798 7358
rect 1210 6716 1800 6728
rect 1210 6662 1274 6716
rect 1680 6662 1800 6716
rect 1210 6642 1800 6662
rect 1036 6524 11218 6576
rect 1036 6390 6960 6524
rect 7198 6390 11218 6524
rect 1036 6332 11218 6390
rect 9214 6262 9798 6290
rect 9214 6200 9346 6262
rect 9638 6200 9798 6262
rect 9214 6190 9798 6200
rect 9188 6054 9818 6086
rect 9188 5826 9242 6054
rect 9736 5826 9818 6054
rect 9188 5800 9818 5826
<< via1 >>
rect 2032 9528 2036 9600
rect 2036 9528 2212 9600
rect 2212 9528 2218 9600
rect 2032 9524 2218 9528
rect 670 8226 826 8318
rect 3134 8828 3194 9130
rect 7070 8452 7168 8508
rect 1922 8222 2336 8336
rect 1078 7362 1134 7670
rect 4672 7984 4736 8044
rect 6764 7676 7376 7732
rect 9730 7358 9784 7424
rect 1274 6662 1680 6716
rect 6960 6390 7198 6524
rect 9346 6200 9638 6262
rect 9242 5826 9736 6054
<< metal2 >>
rect 1432 9600 2816 9646
rect 1432 9524 2032 9600
rect 2218 9524 2816 9600
rect 1432 9224 2816 9524
rect 1056 9130 3204 9224
rect 1056 8828 3134 9130
rect 3194 8828 3204 9130
rect 1056 8734 3204 8828
rect 6690 8508 7584 8744
rect 6690 8452 7070 8508
rect 7168 8452 7584 8508
rect 816 8384 1216 8386
rect 816 8378 3232 8384
rect 400 8336 3232 8378
rect 400 8318 1922 8336
rect 400 8226 670 8318
rect 826 8226 1922 8318
rect 400 8222 1922 8226
rect 2336 8222 3232 8336
rect 400 8174 3232 8222
rect 400 8164 1216 8174
rect 3142 8170 3232 8174
rect 816 8148 1216 8164
rect 6690 8072 7584 8452
rect 4648 8044 9818 8072
rect 4648 7984 4672 8044
rect 4736 7984 9818 8044
rect 4648 7958 9818 7984
rect 1048 7670 3214 7792
rect 1048 7362 1078 7670
rect 1134 7362 3214 7670
rect 4644 7748 9814 7762
rect 4644 7732 6908 7748
rect 7276 7732 9814 7748
rect 4644 7676 6764 7732
rect 7376 7676 9814 7732
rect 4644 7662 6908 7676
rect 7276 7662 9814 7676
rect 4644 7648 9814 7662
rect 1048 7304 3214 7362
rect 4644 7424 9814 7450
rect 4644 7358 9730 7424
rect 9784 7358 9814 7424
rect 4644 7336 9814 7358
rect 1320 6738 1674 7304
rect 1180 6716 1830 6738
rect 1180 6662 1274 6716
rect 1680 6662 1830 6716
rect 1180 6588 1830 6662
rect 6736 6588 7432 6742
rect 9254 6740 9654 7336
rect 1180 6526 7432 6588
rect 1180 6524 6968 6526
rect 1180 6390 6960 6524
rect 7216 6404 7432 6526
rect 7198 6390 7432 6404
rect 1180 6312 7432 6390
rect 1180 6184 1830 6312
rect 6736 6182 7432 6312
rect 9150 6384 9846 6740
rect 9150 6262 9850 6384
rect 9150 6200 9346 6262
rect 9638 6200 9850 6262
rect 9150 6054 9850 6200
rect 9150 5826 9242 6054
rect 9736 5826 9850 6054
rect 9150 5800 9850 5826
<< via2 >>
rect 6908 7732 7276 7748
rect 6908 7676 7276 7732
rect 6908 7662 7276 7676
rect 6968 6524 7216 6526
rect 6968 6404 7198 6524
rect 7198 6404 7216 6524
<< metal3 >>
rect 6848 7748 7356 7762
rect 6848 7662 6908 7748
rect 7276 7662 7356 7748
rect 6848 6526 7356 7662
rect 6848 6404 6968 6526
rect 7216 6404 7356 6526
rect 6848 6362 7356 6404
use sky130_fd_pr__nfet_01v8_lvt_T4BG7Y  XM1
timestamp 1695195131
transform 0 1 6124 -1 0 6460
box -396 -5210 396 5210
use sky130_fd_pr__nfet_01v8_lvt_6TMDZ9  XM2
timestamp 1695195131
transform 1 0 7230 0 1 7704
box -2696 -610 2696 610
use sky130_fd_pr__pfet_01v8_lvt_B5Z988  XM10
timestamp 1695195131
transform 1 0 2134 0 1 8267
box -1196 -1219 1196 1219
<< labels >>
flabel metal1 7022 8384 7222 8584 0 FreeSans 256 0 0 0 Ib
port 1 nsew
flabel metal1 644 8176 844 8376 0 FreeSans 256 0 0 0 Vtune
port 0 nsew
rlabel locali 2212 9386 11320 10390 1 VDD
port 3 nsew
rlabel locali 990 5142 11238 6164 1 GROUND
port 2 nsew
<< end >>
