magic
tech sky130A
timestamp 1696676405
<< metal1 >>
rect 9308 15366 9872 15369
rect 8713 15315 9872 15366
rect 8713 15100 8794 15315
rect 9778 15100 9872 15315
rect 3208 13018 3308 13030
rect 3208 12938 3214 13018
rect 3297 12938 3308 13018
rect 3208 12930 3308 12938
rect 2201 8252 2335 8281
rect 2201 8193 2237 8252
rect 2298 8193 2335 8252
rect 2201 6239 2335 8193
rect 2962 6869 3071 12775
rect 3232 8489 3332 8497
rect 3232 8403 3238 8489
rect 3324 8403 3332 8489
rect 3232 8397 3332 8403
rect 2574 6359 2675 6360
rect 2574 6348 2768 6359
rect 2574 6276 2581 6348
rect 2658 6276 2768 6348
rect 2574 6271 2768 6276
rect 2667 6270 2768 6271
rect 2957 6239 3054 6391
rect 2201 6232 3054 6239
rect 2201 6134 3057 6232
rect 2957 6132 3057 6134
rect 3272 6005 3377 6397
rect 3707 6005 4268 11002
rect 8713 6110 9872 15100
rect 10261 10497 10361 10506
rect 10261 10416 10269 10497
rect 10353 10416 10361 10497
rect 10261 10406 10361 10416
rect 8713 6090 9855 6110
rect 3260 5878 4285 6005
rect 3260 5669 3331 5878
rect 4208 5669 4285 5878
rect 3260 5637 4285 5669
<< via1 >>
rect 8794 15100 9778 15315
rect 3214 12938 3297 13018
rect 2237 8193 2298 8252
rect 3238 8403 3324 8489
rect 2581 6276 2658 6348
rect 10269 10416 10353 10497
rect 3331 5669 4208 5878
<< metal2 >>
rect 2120 15315 10436 16746
rect 2120 15100 8794 15315
rect 9778 15100 10436 15315
rect 2120 15037 10436 15100
rect 2192 8252 2351 8275
rect 2192 8193 2237 8252
rect 2298 8193 2351 8252
rect 2192 8165 2351 8193
rect 2576 6348 2684 15037
rect 4748 13073 4778 13076
rect 3047 13072 4778 13073
rect 3047 13018 5263 13072
rect 3047 12938 3214 13018
rect 3297 12938 5270 13018
rect 3047 12839 5270 12938
rect 3057 12816 5270 12839
rect 2947 12742 3094 12769
rect 2947 12682 2988 12742
rect 3045 12682 3094 12742
rect 2947 12659 3094 12682
rect 4916 12586 5202 12816
rect 5773 12758 5891 12775
rect 5773 12679 5790 12758
rect 5880 12679 5891 12758
rect 5773 12667 5891 12679
rect 7877 10497 10395 14832
rect 7877 10416 10269 10497
rect 10353 10416 10395 10497
rect 3073 8489 4786 8556
rect 3065 8403 3238 8489
rect 3324 8403 5278 8489
rect 3065 8318 5278 8403
rect 4916 8055 5202 8318
rect 5789 8245 5889 8269
rect 5789 8179 5805 8245
rect 5876 8179 5889 8245
rect 5789 8144 5889 8179
rect 2576 6276 2581 6348
rect 2658 6276 2684 6348
rect 2576 6273 2684 6276
rect 7877 6134 10395 10416
rect 2100 5878 10423 5924
rect 2100 5669 3331 5878
rect 4208 5669 10423 5878
rect 2100 4211 10423 5669
<< via2 >>
rect 2237 8193 2298 8252
rect 2988 12682 3045 12742
rect 5790 12679 5880 12758
rect 5805 8179 5876 8245
<< metal3 >>
rect 2947 12758 5902 12781
rect 2947 12742 5790 12758
rect 2947 12682 2988 12742
rect 3045 12682 5790 12742
rect 2947 12679 5790 12682
rect 5880 12679 5902 12758
rect 2947 12656 5902 12679
rect 5775 8279 5905 8283
rect 2180 8252 2576 8279
rect 2180 8193 2237 8252
rect 2298 8193 2576 8252
rect 2180 8154 2576 8193
rect 2684 8245 5905 8279
rect 2684 8179 5805 8245
rect 5876 8179 5905 8245
rect 2684 8154 5905 8179
rect 5775 8141 5905 8154
use not  x1
timestamp 1696661316
transform 0 -1 3093 1 0 6035
box 236 -289 934 518
use switch  x5
timestamp 1696676133
transform 0 1 4161 -1 0 14889
box -20 -459 4321 5137
use switch  x6
timestamp 1696676133
transform 0 1 4170 -1 0 10392
box -20 -459 4321 5137
<< labels >>
flabel metal1 2957 6132 3057 6232 0 FreeSans 128 0 0 0 SEL0
port 0 nsew
flabel metal1 3232 8397 3332 8497 0 FreeSans 128 0 0 0 IN1
port 1 nsew
flabel metal1 10261 10406 10361 10506 0 FreeSans 128 0 0 0 OUT
port 2 nsew
rlabel metal2 2120 15037 10436 16746 1 VDD
port 5 nsew
rlabel metal2 2100 4211 10423 5924 1 GROUND
port 6 nsew
flabel metal1 3208 12930 3308 13030 0 FreeSans 128 0 0 0 IN0
port 3 nsew
<< end >>
