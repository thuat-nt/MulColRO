magic
tech sky130A
magscale 1 2
timestamp 1695440875
<< nwell >>
rect -825 -719 825 719
<< pmoslvt >>
rect -629 -500 -29 500
rect 29 -500 629 500
<< pdiff >>
rect -687 488 -629 500
rect -687 -488 -675 488
rect -641 -488 -629 488
rect -687 -500 -629 -488
rect -29 488 29 500
rect -29 -488 -17 488
rect 17 -488 29 488
rect -29 -500 29 -488
rect 629 488 687 500
rect 629 -488 641 488
rect 675 -488 687 488
rect 629 -500 687 -488
<< pdiffc >>
rect -675 -488 -641 488
rect -17 -488 17 488
rect 641 -488 675 488
<< nsubdiff >>
rect -789 649 -693 683
rect 693 649 789 683
rect -789 587 -755 649
rect 755 587 789 649
rect -789 -649 -755 -587
rect 755 -649 789 -587
rect -789 -683 -693 -649
rect 693 -683 789 -649
<< nsubdiffcont >>
rect -693 649 693 683
rect -789 -587 -755 587
rect 755 -587 789 587
rect -693 -683 693 -649
<< poly >>
rect -629 581 -29 597
rect -629 547 -613 581
rect -45 547 -29 581
rect -629 500 -29 547
rect 29 581 629 597
rect 29 547 45 581
rect 613 547 629 581
rect 29 500 629 547
rect -629 -547 -29 -500
rect -629 -581 -613 -547
rect -45 -581 -29 -547
rect -629 -597 -29 -581
rect 29 -547 629 -500
rect 29 -581 45 -547
rect 613 -581 629 -547
rect 29 -597 629 -581
<< polycont >>
rect -613 547 -45 581
rect 45 547 613 581
rect -613 -581 -45 -547
rect 45 -581 613 -547
<< locali >>
rect -789 649 -693 683
rect 693 649 789 683
rect -789 587 -755 649
rect 755 587 789 649
rect -629 547 -613 581
rect -45 547 -29 581
rect 29 547 45 581
rect 613 547 629 581
rect -675 488 -641 504
rect -675 -504 -641 -488
rect -17 488 17 504
rect -17 -504 17 -488
rect 641 488 675 504
rect 641 -504 675 -488
rect -629 -581 -613 -547
rect -45 -581 -29 -547
rect 29 -581 45 -547
rect 613 -581 629 -547
rect -789 -649 -755 -587
rect 755 -649 789 -587
rect -789 -683 -693 -649
rect 693 -683 789 -649
<< viali >>
rect -613 547 -45 581
rect 45 547 613 581
rect -675 -488 -641 488
rect -17 -488 17 488
rect 641 -488 675 488
rect -613 -581 -45 -547
rect 45 -581 613 -547
<< metal1 >>
rect -625 581 -33 587
rect -625 547 -613 581
rect -45 547 -33 581
rect -625 541 -33 547
rect 33 581 625 587
rect 33 547 45 581
rect 613 547 625 581
rect 33 541 625 547
rect -681 488 -635 500
rect -681 -488 -675 488
rect -641 -488 -635 488
rect -681 -500 -635 -488
rect -23 488 23 500
rect -23 -488 -17 488
rect 17 -488 23 488
rect -23 -500 23 -488
rect 635 488 681 500
rect 635 -488 641 488
rect 675 -488 681 488
rect 635 -500 681 -488
rect -625 -547 -33 -541
rect -625 -581 -613 -547
rect -45 -581 -33 -547
rect -625 -587 -33 -581
rect 33 -547 625 -541
rect 33 -581 45 -547
rect 613 -581 625 -547
rect 33 -587 625 -581
<< labels >>
rlabel poly -629 500 -29 547 1 G
rlabel nsubdiffcont -693 649 693 683 1 B
rlabel locali -675 488 -641 504 1 D
rlabel locali -17 488 17 504 1 S
<< properties >>
string FIXED_BBOX -772 -666 772 666
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 5.0 l 3.0 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
