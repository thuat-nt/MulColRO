magic
tech sky130A
timestamp 1698059410
<< metal1 >>
rect 57623 18942 58045 18988
rect 57623 18296 57672 18942
rect 57995 18296 58045 18942
rect 57623 3779 58045 18296
rect 58315 9617 59176 9659
rect 58315 9467 58621 9617
rect 58869 9467 59176 9617
rect 58315 9413 59176 9467
rect 57623 3772 58745 3779
rect 57623 3255 58755 3772
rect 58355 -3096 58755 3255
rect 62280 -3381 62784 -1071
rect 62280 -3670 62313 -3381
rect 62755 -3670 62784 -3381
rect 62280 -3706 62784 -3670
<< via1 >>
rect 57672 18296 57995 18942
rect 58621 9467 58869 9617
rect 62313 -3670 62755 -3381
<< metal2 >>
rect 19319 25742 65574 26370
rect 19319 23492 37366 25742
rect 42889 23492 65574 25742
rect 19319 20274 65574 23492
rect 19284 18942 65574 20274
rect 19284 18678 57672 18942
rect 17147 18076 17722 18214
rect 17147 16936 17253 18076
rect 17636 16936 17722 18076
rect 15946 11863 16820 11866
rect 4827 11859 16820 11863
rect 4827 11675 16832 11859
rect 4827 10740 5044 11675
rect 5899 10740 16832 11675
rect 4827 10485 16832 10740
rect 15946 600 16820 10485
rect 17147 7203 17722 16936
rect 19284 16395 38912 18678
rect 53011 18296 57672 18678
rect 57995 18678 65574 18942
rect 57995 18296 59002 18678
rect 53011 18178 59002 18296
rect 58535 9617 58943 9664
rect 58535 9467 58621 9617
rect 58869 9467 58943 9617
rect 58535 9418 58943 9467
rect 17147 7001 19308 7203
rect 17147 6245 18776 7001
rect 19159 6245 19308 7001
rect 17147 6106 19308 6245
rect 15946 527 18450 600
rect 15946 139 18112 527
rect 18376 139 18450 527
rect 15946 71 18450 139
rect 20551 -2749 37374 1499
rect 62048 -2513 62288 -2471
rect 62048 -2726 62072 -2513
rect 62244 -2726 62288 -2513
rect 20295 -3288 57589 -2749
rect 62048 -2759 62288 -2726
rect 20295 -3379 62795 -3288
rect 63115 -3379 65005 9302
rect 20295 -3381 65005 -3379
rect 20295 -3670 62313 -3381
rect 62755 -3670 65005 -3381
rect 20295 -6171 65005 -3670
rect 20295 -7046 38742 -6171
rect 20352 -8421 38742 -7046
rect 44265 -8421 65005 -6171
rect 20352 -9138 65005 -8421
rect 20352 -9280 64864 -9138
<< via2 >>
rect 37366 23492 42889 25742
rect 17253 16936 17636 18076
rect 5044 10740 5899 11675
rect 59240 16264 59470 16480
rect 59330 11787 59472 11961
rect 66031 10139 66434 17957
rect 58621 9467 58869 9617
rect 18776 6245 19159 7001
rect 18112 139 18376 527
rect 62072 -2726 62244 -2513
rect 38742 -8421 44265 -6171
<< metal3 >>
rect 36827 25742 43556 26184
rect 36827 23492 37366 25742
rect 42889 23492 43556 25742
rect 36827 23021 43556 23492
rect 36979 21707 38111 21859
rect 36979 20642 37198 21707
rect 37942 20642 38111 21707
rect 17189 18076 17732 18182
rect 17189 16936 17253 18076
rect 17636 16936 17732 18076
rect 17189 16798 17732 16936
rect 17164 15920 17687 16112
rect 17164 14885 17282 15920
rect 17602 14885 17687 15920
rect 4782 13804 16882 14023
rect 4782 12833 4980 13804
rect 5891 12833 16882 13804
rect 4782 12606 16882 12833
rect 4927 11675 5998 11785
rect 4927 10740 5044 11675
rect 5899 10740 5998 11675
rect 4927 10592 5998 10740
rect 15927 -183 16850 12606
rect 17164 12184 17687 14885
rect 36979 13214 38111 20642
rect 65896 17957 66548 18187
rect 59216 16480 59502 16493
rect 59216 16264 59240 16480
rect 59470 16264 59502 16480
rect 59216 16250 59502 16264
rect 17164 11790 19405 12184
rect 35003 11893 38111 13214
rect 59307 11961 59510 11978
rect 35003 11381 38069 11893
rect 59307 11787 59330 11961
rect 59472 11787 59510 11961
rect 59307 11766 59510 11787
rect 35003 10776 37259 11381
rect 37971 10776 38069 11381
rect 35003 10693 38069 10776
rect 65896 10139 66031 17957
rect 66434 10139 66548 17957
rect 65896 9986 66548 10139
rect 58535 9617 58943 9664
rect 58535 9467 58621 9617
rect 58869 9467 58943 9617
rect 58535 9418 58943 9467
rect 18691 7001 19330 7192
rect 18691 6245 18776 7001
rect 19159 6245 19330 7001
rect 18691 6095 19330 6245
rect 56856 3249 57526 3251
rect 37301 600 37794 3246
rect 56856 2795 59121 3249
rect 18050 527 37794 600
rect 18050 139 18112 527
rect 18376 139 37794 527
rect 18050 77 37794 139
rect 37301 59 37794 77
rect 15927 -199 47425 -183
rect 56856 -199 57526 2795
rect 15927 -805 57526 -199
rect 15927 -806 47425 -805
rect 56856 -813 57526 -805
rect 60524 -929 60722 -807
rect 62043 -2360 62326 -2283
rect 62043 -2513 62074 -2360
rect 62043 -2726 62072 -2513
rect 62043 -2851 62074 -2726
rect 62271 -2851 62326 -2360
rect 62043 -2927 62326 -2851
rect 37825 -6171 44986 -5785
rect 37825 -8421 38742 -6171
rect 44265 -8421 44986 -6171
rect 37825 -8936 44986 -8421
<< via3 >>
rect 37366 23492 42889 25742
rect 37198 20642 37942 21707
rect 17253 16936 17636 18076
rect 17282 14885 17602 15920
rect 4980 12833 5891 13804
rect 5044 10740 5899 11675
rect 18970 13719 19191 14755
rect 39425 16602 39886 17086
rect 59240 16264 59470 16480
rect 39439 15480 39900 15964
rect 39460 12098 39921 12582
rect 59330 11787 59472 11961
rect 37259 10776 37971 11381
rect 39453 11018 39914 11502
rect 39467 9938 39928 10422
rect 66031 10139 66434 17957
rect 58621 9467 58869 9617
rect 18887 3254 19451 3965
rect 39320 1119 39784 1590
rect 62074 -2513 62271 -2360
rect 62074 -2726 62244 -2513
rect 62244 -2726 62271 -2513
rect 62074 -2851 62271 -2726
rect 38742 -8421 44265 -6171
<< metal4 >>
rect 36827 25742 43556 26184
rect 36827 23492 37366 25742
rect 42889 23492 43556 25742
rect 36827 23021 43556 23492
rect 15813 22390 16984 22555
rect 15813 21186 15970 22390
rect 16800 21186 16984 22390
rect 4896 13804 5967 13914
rect 4896 12833 4980 13804
rect 5891 12833 5967 13804
rect 4896 12721 5967 12833
rect 4927 11675 5998 11785
rect 4927 10740 5044 11675
rect 5899 10740 5998 11675
rect 4927 10592 5998 10740
rect 4737 9427 15548 9688
rect 4737 8565 4948 9427
rect 5784 8565 15548 9427
rect 4737 8273 15548 8565
rect 14723 1653 15548 8273
rect 15813 4446 16984 21186
rect 37063 21707 38111 21859
rect 37063 20642 37198 21707
rect 37942 20642 38111 21707
rect 37063 20440 38111 20642
rect 17902 20159 19186 20212
rect 17902 19055 18093 20159
rect 18931 19055 19186 20159
rect 17189 18076 17732 18182
rect 17189 16936 17253 18076
rect 17636 16936 17732 18076
rect 17189 16798 17732 16936
rect 17175 15920 17708 16101
rect 17175 14885 17282 15920
rect 17602 14885 17708 15920
rect 17175 14778 17708 14885
rect 17902 14992 19186 19055
rect 63664 17957 66501 18281
rect 39319 17086 40024 17220
rect 39319 16602 39425 17086
rect 39886 16602 40024 17086
rect 39319 16471 40024 16602
rect 59216 16480 59502 16493
rect 59216 16264 59240 16480
rect 59470 16264 59502 16480
rect 59216 16250 59502 16264
rect 39330 15964 40035 16085
rect 39330 15480 39439 15964
rect 39900 15480 40035 15964
rect 39330 15336 40035 15480
rect 17902 14755 19249 14992
rect 17902 13719 18970 14755
rect 19191 13719 19249 14755
rect 17902 13465 19249 13719
rect 39341 12582 40046 12725
rect 39341 12098 39460 12582
rect 39921 12098 40046 12582
rect 39341 11976 40046 12098
rect 56694 11961 59814 13302
rect 56694 11787 59330 11961
rect 59472 11787 59814 11961
rect 56694 11728 59814 11787
rect 39345 11502 40050 11626
rect 37145 11381 38069 11471
rect 37145 10776 37259 11381
rect 37971 10776 38069 11381
rect 39345 11018 39453 11502
rect 39914 11018 40050 11502
rect 39345 10877 40050 11018
rect 37145 9737 38069 10776
rect 39348 10422 40053 10567
rect 39348 9938 39467 10422
rect 39928 9938 40053 10422
rect 39348 9818 40053 9938
rect 63664 10139 66031 17957
rect 66434 10139 66501 17957
rect 58535 9617 58943 9664
rect 58535 9467 58621 9617
rect 58869 9467 58943 9617
rect 58535 9418 58943 9467
rect 63664 5887 66501 10139
rect 15813 3965 19702 4446
rect 15813 3254 18887 3965
rect 19451 3254 19702 3965
rect 59975 3517 66501 5887
rect 59975 3365 66498 3517
rect 15813 2794 19702 3254
rect 14723 1590 39835 1653
rect 14723 1119 39320 1590
rect 39784 1119 39835 1590
rect 14723 1074 39835 1119
rect 62058 -1806 62498 -1728
rect 62058 -2360 62101 -1806
rect 62058 -2851 62074 -2360
rect 62058 -3023 62101 -2851
rect 62423 -3023 62498 -1806
rect 62058 -3086 62498 -3023
rect 37825 -6171 44986 -5785
rect 37825 -8421 38742 -6171
rect 44265 -8421 44986 -6171
rect 37825 -8936 44986 -8421
<< via4 >>
rect 37366 23492 42889 25742
rect 15970 21186 16800 22390
rect 4980 12833 5891 13804
rect 5044 10740 5899 11675
rect 4948 8565 5784 9427
rect 37198 20642 37942 21707
rect 18093 19055 18931 20159
rect 17253 16936 17636 18076
rect 17282 14885 17602 15920
rect 39425 16602 39886 17086
rect 59240 16264 59470 16480
rect 39439 15480 39900 15964
rect 39460 12098 39921 12582
rect 39453 11018 39914 11502
rect 39467 9938 39928 10422
rect 58621 9467 58869 9617
rect 62101 -2360 62423 -1806
rect 62101 -2851 62271 -2360
rect 62271 -2851 62423 -2360
rect 62101 -3023 62423 -2851
rect 38742 -8421 44265 -6171
<< metal5 >>
rect 17869 25742 65634 26337
rect 17869 23492 37366 25742
rect 42889 23492 65634 25742
rect 17869 22808 65634 23492
rect 4768 22492 6091 22497
rect 4768 22488 6579 22492
rect 15740 22488 16963 22492
rect 4768 22390 17006 22488
rect 4768 21186 15970 22390
rect 16800 21186 17006 22390
rect 4768 21111 17006 21186
rect 4770 21091 17006 21111
rect 37030 21707 59798 21859
rect 37030 20642 37198 21707
rect 37942 20642 59798 21707
rect 37030 20457 59798 20642
rect 4784 20279 6579 20286
rect 15740 20279 19154 20286
rect 4784 20159 19154 20279
rect 4784 19055 18093 20159
rect 18931 19055 19154 20159
rect 4784 18907 19154 19055
rect 4800 18894 6123 18907
rect 4782 18182 6105 18190
rect 4782 18169 6579 18182
rect 15740 18169 17711 18182
rect 4782 18076 17711 18169
rect 4782 16936 17253 18076
rect 17636 16936 17711 18076
rect 4782 16804 17711 16936
rect 39259 17209 43875 17264
rect 39259 17086 43888 17209
rect 39259 16602 39425 17086
rect 39886 16602 43888 17086
rect 39259 16416 43888 16602
rect 4782 16112 6105 16114
rect 4782 16108 6579 16112
rect 15740 16108 17698 16112
rect 4782 15920 17698 16108
rect 4782 14885 17282 15920
rect 17602 14885 17698 15920
rect 39270 16088 42619 16128
rect 39270 15964 42631 16088
rect 39270 15480 39439 15964
rect 39900 15480 42631 15964
rect 39270 15306 42631 15480
rect 4782 14728 17698 14885
rect 4782 13804 6105 13992
rect 4782 12833 4980 13804
rect 5891 12833 6105 13804
rect 4782 12606 6105 12833
rect 6723 12821 8080 12899
rect 6723 12582 40092 12821
rect 6723 12098 39460 12582
rect 39921 12098 40092 12582
rect 6723 11907 40092 12098
rect 4827 11675 6150 11871
rect 4827 10740 5044 11675
rect 5899 10740 6150 11675
rect 4827 10485 6150 10740
rect 4737 9427 6060 9659
rect 4737 8565 4948 9427
rect 5784 8565 6060 9427
rect 4737 8273 6060 8565
rect 6723 7469 8080 11907
rect 40450 11668 41373 11669
rect 39292 11502 41394 11668
rect 39292 11018 39453 11502
rect 39914 11018 41394 11502
rect 39292 10835 41394 11018
rect 8908 10589 9899 10633
rect 8892 10422 40107 10589
rect 8892 9938 39467 10422
rect 39928 9938 40107 10422
rect 8892 9766 40107 9938
rect 4737 6062 8081 7469
rect 8908 5250 9899 9766
rect 4691 3850 9925 5250
rect 4691 3005 6014 3025
rect 40450 3005 41373 10835
rect 4691 1910 41373 3005
rect 4691 1642 41370 1910
rect 4691 1639 41316 1642
rect 41556 816 42631 15306
rect 4646 -562 42631 816
rect 4646 -573 42407 -562
rect 43008 -1336 43888 16416
rect 57957 16480 59798 20457
rect 57957 16264 59240 16480
rect 59470 16264 59798 16480
rect 57957 16200 59798 16264
rect 58318 9617 59170 9661
rect 58318 9467 58621 9617
rect 58869 9467 59170 9617
rect 4556 -2739 43889 -1336
rect 58318 -3444 59170 9467
rect 62050 -1721 62931 -1714
rect 66613 -1721 67981 -1711
rect 62050 -1806 67981 -1721
rect 62050 -3023 62101 -1806
rect 62423 -3023 67981 -1806
rect 62050 -3097 67981 -3023
rect 62050 -3106 67975 -3097
rect 62473 -3111 67975 -3106
rect 4511 -4861 60239 -3444
rect 58318 -4865 59170 -4861
rect 17282 -6171 65047 -5619
rect 17282 -8421 38742 -6171
rect 44265 -8421 65047 -6171
rect 17282 -9148 65047 -8421
use diffamp  x1
timestamp 1696157832
transform 1 0 5022 0 1 15569
box 13700 -15857 30592 2342
use integrator  x2
timestamp 1698059410
transform 1 0 28984 0 1 2100
box 7314 -5062 28629 18146
use mux2_1  x3
timestamp 1698059410
transform 1 0 56116 0 1 3427
box 2100 4211 10436 16746
use buffer  x7
timestamp 1698059410
transform 0 -1 63946 -1 0 6377
box 2815 1163 9644 5591
<< labels >>
rlabel metal5 17282 -9148 65047 -5619 1 VSS
port 2 nsew
rlabel metal5 17869 22808 65634 26337 1 VDD
port 1 nsew
rlabel metal5 4768 21111 6091 22497 1 AIn0
port 3 nsew
rlabel metal5 4800 18894 6123 20280 1 AIn1
port 4 nsew
rlabel metal5 4782 16804 6105 18190 1 AIn2
port 5 nsew
rlabel metal5 4782 14728 6105 16114 1 AIn3
port 6 nsew
rlabel metal5 4782 12606 6105 13992 1 AIn4
port 7 nsew
rlabel metal5 4827 10485 6150 11871 1 AIn5
port 8 nsew
rlabel metal5 4737 8273 6060 9659 1 REG0
port 9 nsew
rlabel metal5 4737 6062 6060 7448 1 REG1
port 10 nsew
rlabel metal5 4691 3850 6014 5236 1 REG2
port 11 nsew
rlabel metal5 4691 1639 6014 3025 1 REG3
port 12 nsew
rlabel metal5 4646 -573 5969 813 1 REG4
port 13 nsew
rlabel metal5 4556 -2739 5879 -1353 1 REG5
port 14 nsew
rlabel metal5 4511 -4861 5834 -3475 1 REG6
port 15 nsew
rlabel metal5 66658 -3097 67981 -1711 1 AOut
port 16 nsew
<< end >>
