magic
tech sky130A
timestamp 1695566345
<< metal5 >>
rect 159883 79815 160788 79848
rect 158076 79781 160788 79815
rect 158076 77707 230680 79781
rect 158076 77630 160788 77707
rect 158107 32740 159113 77630
rect 159883 68485 160788 77630
rect 158107 31332 161324 32740
rect 227664 32673 228535 77707
rect 229791 68682 230680 77707
rect 227664 31332 231149 32673
use ColROs  x1
timestamp 1695566025
transform 1 0 155113 0 1 47394
box 4511 -9280 67981 26370
use ColROs  x2
timestamp 1695566025
transform 1 0 155163 0 1 10210
box 4511 -9280 67981 26370
use ColROs  x3
timestamp 1695566025
transform 1 0 224981 0 1 10215
box 4511 -9280 67981 26370
use ColROs  x5
timestamp 1695566025
transform 1 0 225021 0 1 47591
box 4511 -9280 67981 26370
<< labels >>
rlabel metal5 158076 77630 160430 79815 1 REF
port 1 nsew
<< end >>
