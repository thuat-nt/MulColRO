magic
tech sky130A
magscale 1 2
timestamp 1695377223
<< error_p >>
rect 253023 62300 253058 62334
rect 253024 62281 253058 62300
rect 236957 62142 236992 62176
rect 236958 62123 236992 62142
rect 235380 60863 235395 61729
rect 235414 60863 235448 61783
rect 235414 60829 235429 60863
rect 236977 60810 236992 62123
rect 237011 62089 237046 62123
rect 237011 60810 237045 62089
rect 244380 61983 244415 62017
rect 246689 62000 246723 62018
rect 244381 61964 244415 61983
rect 237011 60776 237026 60810
rect 244400 60651 244415 61964
rect 244434 61930 244469 61964
rect 244434 60651 244468 61930
rect 244434 60617 244449 60651
rect 246653 60598 246723 62000
rect 250207 61840 250241 61894
rect 246653 60562 246706 60598
rect 250226 60545 250241 61840
rect 250260 61806 250295 61840
rect 251145 61806 251180 61840
rect 250260 60545 250294 61806
rect 251146 61787 251180 61806
rect 250260 60511 250275 60545
rect 251165 60492 251180 61787
rect 251199 61753 251234 61787
rect 251199 60492 251233 61753
rect 251199 60458 251214 60492
rect 252104 60439 252119 61787
rect 252138 60439 252172 61841
rect 252138 60405 252153 60439
rect 253043 60386 253058 62281
rect 253077 62247 253112 62281
rect 253077 60386 253111 62247
rect 261956 60926 261958 62328
rect 262059 60450 262728 68865
rect 262824 66988 262830 68340
rect 269982 60926 269984 62328
rect 270085 60450 270754 68865
rect 270850 66988 270856 68340
rect 278606 60486 278744 60504
rect 278640 60452 278778 60470
rect 253077 60352 253092 60386
rect 278648 59526 278668 59782
rect 278676 59554 278724 59754
rect 66576 51260 72496 55460
rect 76422 55009 76456 59113
rect 77097 55082 77119 55299
rect 77541 55082 77559 55299
rect 77119 55009 77541 55045
rect 74558 54998 77541 55009
rect 77939 54998 78146 55045
rect 74558 54975 78146 54998
rect 74399 51350 74401 52752
rect 72535 51300 72536 51301
rect 72784 51300 72848 51316
rect 72536 51299 72537 51300
rect 72848 51260 72864 51300
rect 66576 50877 74150 51260
rect 74558 50877 74592 54975
rect 74992 54923 75039 54954
rect 74980 54907 75039 54923
rect 75302 54907 75349 54954
rect 75650 54923 75697 54954
rect 75638 54907 75697 54923
rect 75960 54907 76007 54954
rect 76308 54923 76354 54954
rect 76296 54907 76354 54923
rect 74734 54873 75349 54907
rect 75392 54873 76007 54907
rect 76050 54873 76354 54907
rect 74980 54826 75038 54873
rect 75638 54826 75696 54873
rect 76296 54826 76354 54873
rect 74661 54814 74706 54825
rect 74672 51026 74706 54814
rect 74992 51038 75026 54826
rect 75319 54814 75364 54825
rect 75330 51026 75364 54814
rect 75650 51038 75684 54826
rect 75977 54814 76022 54825
rect 75988 51026 76022 54814
rect 76308 51038 76342 54826
rect 74660 50979 74719 51026
rect 74964 50979 75011 51026
rect 75318 50979 75377 51026
rect 75622 50979 75669 51026
rect 75976 50979 76035 51026
rect 76280 50979 76327 51026
rect 74660 50945 75011 50979
rect 75054 50945 75669 50979
rect 75712 50945 76327 50979
rect 74660 50929 74718 50945
rect 75318 50929 75376 50945
rect 75976 50929 76034 50945
rect 74660 50914 74675 50929
rect 74672 50877 74706 50911
rect 75330 50877 75364 50911
rect 75988 50877 76022 50911
rect 76422 50877 76456 54975
rect 76515 54946 76613 54975
rect 76487 54918 76557 54926
rect 76597 53174 76613 54526
rect 77119 54448 77541 54975
rect 77879 54867 77919 54882
rect 77879 54839 77891 54854
rect 66576 50843 76456 50877
rect 77939 50968 78146 54975
rect 78755 51520 78781 51708
rect 78789 51520 78815 51674
rect 79405 51576 79439 59028
rect 80894 55050 81563 59245
rect 86097 59180 87701 59214
rect 81659 57368 81665 58720
rect 80894 55014 83217 55050
rect 79629 54980 83217 55014
rect 78751 51110 79213 51520
rect 78713 51012 78727 51110
rect 78741 51040 79213 51110
rect 79405 51494 79509 51576
rect 79405 51052 79439 51494
rect 78151 50968 78397 50974
rect 77939 50962 78629 50968
rect 77939 50900 78146 50962
rect 78221 50956 78629 50962
rect 78169 50940 78369 50946
rect 78169 50934 78629 50940
rect 78193 50928 78629 50934
rect 78751 50900 79213 51040
rect 79297 50962 79389 50986
rect 79455 50962 79553 50986
rect 79297 50960 79321 50962
rect 79325 50934 79417 50958
rect 79427 50934 79525 50958
rect 79531 50956 79553 50962
rect 79325 50932 79349 50934
rect 79475 50900 79525 50934
rect 79629 50900 79663 54980
rect 80063 54928 80101 54950
rect 80051 54912 80109 54928
rect 80373 54912 80411 54950
rect 80721 54928 80759 54950
rect 80709 54912 80767 54928
rect 80894 54912 83217 54980
rect 79805 54878 80411 54912
rect 80463 54878 83217 54912
rect 80051 54840 80109 54878
rect 80709 54840 80767 54878
rect 79732 54828 79777 54839
rect 79743 51040 79777 54828
rect 80063 51052 80097 54840
rect 80390 54828 80435 54839
rect 80401 51040 80435 54828
rect 80721 51052 80755 54840
rect 79731 51002 79789 51040
rect 80035 51002 80073 51040
rect 80389 51002 80447 51040
rect 80693 51002 80731 51040
rect 80894 51002 83217 54878
rect 88817 51306 88819 52708
rect 79731 50968 80073 51002
rect 80125 50968 80731 51002
rect 80783 50968 83217 51002
rect 79731 50952 79789 50968
rect 80389 50952 80447 50968
rect 79731 50937 79746 50952
rect 79743 50900 79777 50934
rect 80401 50900 80435 50934
rect 80894 50900 83217 50968
rect 77939 50866 83217 50900
rect 86097 50866 87487 50900
rect 66576 49540 74150 50843
rect 68189 49500 68190 49501
rect 68190 49499 68191 49500
rect 68230 48860 74150 49540
rect 74558 48860 74592 50843
rect 77939 50830 78146 50866
rect 79629 48860 79663 50866
rect 80894 50807 83217 50866
rect 88920 50830 89589 55045
rect 89685 53168 89691 54520
rect 119439 52680 119474 52714
rect 119440 52661 119474 52680
rect 103373 52522 103408 52556
rect 103374 52503 103408 52522
rect 101796 51243 101811 52109
rect 101830 51243 101864 52163
rect 101830 51209 101845 51243
rect 103393 51190 103408 52503
rect 103427 52469 103462 52503
rect 103427 51190 103461 52469
rect 110796 52363 110831 52397
rect 113105 52380 113139 52398
rect 110797 52344 110831 52363
rect 94027 49834 94061 50174
rect 97545 49094 97579 51186
rect 103427 51156 103442 51190
rect 110816 51031 110831 52344
rect 110850 52310 110885 52344
rect 110850 51031 110884 52310
rect 110850 50997 110865 51031
rect 113069 50978 113139 52380
rect 116623 52220 116657 52274
rect 113069 50942 113122 50978
rect 116642 50925 116657 52220
rect 116676 52186 116711 52220
rect 117561 52186 117596 52220
rect 116676 50925 116710 52186
rect 117562 52167 117596 52186
rect 116676 50891 116691 50925
rect 117581 50872 117596 52167
rect 117615 52133 117650 52167
rect 117615 50872 117649 52133
rect 117615 50838 117630 50872
rect 118520 50819 118535 52167
rect 118554 50819 118588 52221
rect 118554 50785 118569 50819
rect 119459 50766 119474 52661
rect 119493 52627 119528 52661
rect 119493 50766 119527 52627
rect 128372 51306 128374 52708
rect 128475 50830 129144 59245
rect 129240 57368 129246 58720
rect 136996 50866 137134 50884
rect 137030 50832 137168 50850
rect 119493 50732 119508 50766
rect 283023 15912 283058 15946
rect 283024 15893 283058 15912
rect 266957 15754 266992 15788
rect 266958 15735 266992 15754
rect 265380 14475 265395 15341
rect 265414 14475 265448 15395
rect 265414 14441 265429 14475
rect 266977 14422 266992 15735
rect 267011 15701 267046 15735
rect 267011 14422 267045 15701
rect 274380 15595 274415 15629
rect 276689 15612 276723 15630
rect 274381 15576 274415 15595
rect 267011 14388 267026 14422
rect 274400 14263 274415 15576
rect 274434 15542 274469 15576
rect 274434 14263 274468 15542
rect 274434 14229 274449 14263
rect 276653 14210 276723 15612
rect 280207 15452 280241 15506
rect 276653 14174 276706 14210
rect 280226 14157 280241 15452
rect 280260 15418 280295 15452
rect 281145 15418 281180 15452
rect 280260 14157 280294 15418
rect 281146 15399 281180 15418
rect 280260 14123 280275 14157
rect 281165 14104 281180 15399
rect 281199 15365 281234 15399
rect 281199 14104 281233 15365
rect 281199 14070 281214 14104
rect 282104 14051 282119 15399
rect 282138 14051 282172 15453
rect 282138 14017 282153 14051
rect 283043 13998 283058 15893
rect 283077 15859 283112 15893
rect 283077 13998 283111 15859
rect 283077 13964 283092 13998
rect 170785 5176 170820 5210
rect 170786 5157 170820 5176
rect 154719 5018 154754 5052
rect 154720 4999 154754 5018
rect 153142 3739 153157 4605
rect 153176 3739 153210 4659
rect 153176 3705 153191 3739
rect 154739 3686 154754 4999
rect 154773 4965 154808 4999
rect 154773 3686 154807 4965
rect 162142 4859 162177 4893
rect 164451 4876 164485 4894
rect 162143 4840 162177 4859
rect 154773 3652 154788 3686
rect 162162 3527 162177 4840
rect 162196 4806 162231 4840
rect 162196 3527 162230 4806
rect 162196 3493 162211 3527
rect 164415 3474 164485 4876
rect 167969 4716 168003 4770
rect 164415 3438 164468 3474
rect 167988 3421 168003 4716
rect 168022 4682 168057 4716
rect 168907 4682 168942 4716
rect 168022 3421 168056 4682
rect 168908 4663 168942 4682
rect 168022 3387 168037 3421
rect 168927 3368 168942 4663
rect 168961 4629 168996 4663
rect 168961 3368 168995 4629
rect 168961 3334 168976 3368
rect 169866 3315 169881 4663
rect 169900 3315 169934 4717
rect 169900 3281 169915 3315
rect 170805 3262 170820 5157
rect 170839 5123 170874 5157
rect 170839 3262 170873 5123
rect 179718 3802 179720 5204
rect 179821 3326 180490 11741
rect 180586 9864 180592 11216
rect 187744 3802 187746 5204
rect 187847 3326 188516 11741
rect 188612 9864 188618 11216
rect 195770 3802 195772 5204
rect 195873 3326 196542 11741
rect 196638 9864 196644 11216
rect 170839 3228 170854 3262
use diffamp  x1
timestamp 1695351391
transform 1 0 53 0 1 2200
box 28606 -27970 57968 1616
use integrator  x2
timestamp 1695316725
transform 1 0 60124 0 1 48860
box 0 -3600 78298 10660
use cds  x4
timestamp 1695365668
transform 1 0 135992 0 1 1356
box 0 -1600 68576 12818
use s&h  x5
timestamp 1695365668
transform 1 0 224602 0 1 58480
box 0 -1200 57092 12818
use mux4_1  x6
timestamp 1695377223
transform 1 0 246874 0 1 -25244
box 23126 -7250 55042 27920
use buffer  x7
timestamp 1695307921
transform 1 0 260974 0 1 12092
box 0 -800 23059 10496
<< end >>
