magic
tech sky130A
magscale 1 2
timestamp 1696652587
<< error_p >>
rect -31 172 31 178
rect -31 138 -19 172
rect -31 132 31 138
rect -31 -138 31 -132
rect -31 -172 -19 -138
rect -31 -178 31 -172
<< pwell >>
rect -231 -310 231 310
<< nmoslvt >>
rect -35 -100 35 100
<< ndiff >>
rect -93 88 -35 100
rect -93 -88 -81 88
rect -47 -88 -35 88
rect -93 -100 -35 -88
rect 35 88 93 100
rect 35 -88 47 88
rect 81 -88 93 88
rect 35 -100 93 -88
<< ndiffc >>
rect -81 -88 -47 88
rect 47 -88 81 88
<< psubdiff >>
rect -195 240 -99 274
rect 99 240 195 274
rect -195 178 -161 240
rect 161 178 195 240
rect -195 -240 -161 -178
rect 161 -240 195 -178
rect -195 -274 -99 -240
rect 99 -274 195 -240
<< psubdiffcont >>
rect -99 240 99 274
rect -195 -178 -161 178
rect 161 -178 195 178
rect -99 -274 99 -240
<< poly >>
rect -35 172 35 188
rect -35 138 -19 172
rect 19 138 35 172
rect -35 100 35 138
rect -35 -138 35 -100
rect -35 -172 -19 -138
rect 19 -172 35 -138
rect -35 -188 35 -172
<< polycont >>
rect -19 138 19 172
rect -19 -172 19 -138
<< locali >>
rect -195 240 -99 274
rect 99 240 195 274
rect -195 178 -161 240
rect 161 178 195 240
rect -35 138 -19 172
rect 19 138 35 172
rect -81 88 -47 104
rect -81 -104 -47 -88
rect 47 88 81 104
rect 47 -104 81 -88
rect -35 -172 -19 -138
rect 19 -172 35 -138
rect -195 -240 -161 -178
rect 161 -240 195 -178
rect -195 -274 -99 -240
rect 99 -274 195 -240
<< viali >>
rect -19 138 19 172
rect -81 -88 -47 88
rect 47 -88 81 88
rect -19 -172 19 -138
<< metal1 >>
rect -31 172 31 178
rect -31 138 -19 172
rect 19 138 31 172
rect -31 132 31 138
rect -87 88 -41 100
rect -87 -88 -81 88
rect -47 -88 -41 88
rect -87 -100 -41 -88
rect 41 88 87 100
rect 41 -88 47 88
rect 81 -88 87 88
rect 41 -100 87 -88
rect -31 -138 31 -132
rect -31 -172 -19 -138
rect 19 -172 31 -138
rect -31 -178 31 -172
<< properties >>
string FIXED_BBOX -178 -257 178 257
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 1.0 l 0.35 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
