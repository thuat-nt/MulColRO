magic
tech sky130A
magscale 1 2
timestamp 1695908076
<< nwell >>
rect -1154 -719 1154 719
<< pmoslvt >>
rect -958 -500 -358 500
rect -300 -500 300 500
rect 358 -500 958 500
<< pdiff >>
rect -1016 488 -958 500
rect -1016 -488 -1004 488
rect -970 -488 -958 488
rect -1016 -500 -958 -488
rect -358 488 -300 500
rect -358 -488 -346 488
rect -312 -488 -300 488
rect -358 -500 -300 -488
rect 300 488 358 500
rect 300 -488 312 488
rect 346 -488 358 488
rect 300 -500 358 -488
rect 958 488 1016 500
rect 958 -488 970 488
rect 1004 -488 1016 488
rect 958 -500 1016 -488
<< pdiffc >>
rect -1004 -488 -970 488
rect -346 -488 -312 488
rect 312 -488 346 488
rect 970 -488 1004 488
<< nsubdiff >>
rect -1118 649 -1022 683
rect 1022 649 1118 683
rect -1118 587 -1084 649
rect 1084 587 1118 649
rect -1118 -649 -1084 -587
rect 1084 -649 1118 -587
rect -1118 -683 -1022 -649
rect 1022 -683 1118 -649
<< nsubdiffcont >>
rect -1022 649 1022 683
rect -1118 -587 -1084 587
rect 1084 -587 1118 587
rect -1022 -683 1022 -649
<< poly >>
rect -958 581 -358 597
rect -958 547 -942 581
rect -374 547 -358 581
rect -958 500 -358 547
rect -300 581 300 597
rect -300 547 -284 581
rect 284 547 300 581
rect -300 500 300 547
rect 358 581 958 597
rect 358 547 374 581
rect 942 547 958 581
rect 358 500 958 547
rect -958 -547 -358 -500
rect -958 -581 -942 -547
rect -374 -581 -358 -547
rect -958 -597 -358 -581
rect -300 -547 300 -500
rect -300 -581 -284 -547
rect 284 -581 300 -547
rect -300 -597 300 -581
rect 358 -547 958 -500
rect 358 -581 374 -547
rect 942 -581 958 -547
rect 358 -597 958 -581
<< polycont >>
rect -942 547 -374 581
rect -284 547 284 581
rect 374 547 942 581
rect -942 -581 -374 -547
rect -284 -581 284 -547
rect 374 -581 942 -547
<< locali >>
rect -1118 649 -1022 683
rect 1022 649 1118 683
rect -1118 587 -1084 649
rect 1084 587 1118 649
rect -958 547 -942 581
rect -374 547 -358 581
rect -300 547 -284 581
rect 284 547 300 581
rect 358 547 374 581
rect 942 547 958 581
rect -1004 488 -970 504
rect -1004 -504 -970 -488
rect -346 488 -312 504
rect -346 -504 -312 -488
rect 312 488 346 504
rect 312 -504 346 -488
rect 970 488 1004 504
rect 970 -504 1004 -488
rect -958 -581 -942 -547
rect -374 -581 -358 -547
rect -300 -581 -284 -547
rect 284 -581 300 -547
rect 358 -581 374 -547
rect 942 -581 958 -547
rect -1118 -649 -1084 -587
rect 1084 -649 1118 -587
rect -1118 -683 -1022 -649
rect 1022 -683 1118 -649
<< viali >>
rect -942 547 -374 581
rect -284 547 284 581
rect 374 547 942 581
rect -1004 -488 -970 488
rect -346 -488 -312 488
rect 312 -488 346 488
rect 970 -488 1004 488
rect -942 -581 -374 -547
rect -284 -581 284 -547
rect 374 -581 942 -547
<< metal1 >>
rect -954 581 -362 587
rect -954 547 -942 581
rect -374 547 -362 581
rect -954 541 -362 547
rect -296 581 296 587
rect -296 547 -284 581
rect 284 547 296 581
rect -296 541 296 547
rect 362 581 954 587
rect 362 547 374 581
rect 942 547 954 581
rect 362 541 954 547
rect -1010 488 -964 500
rect -1010 -488 -1004 488
rect -970 -488 -964 488
rect -1010 -500 -964 -488
rect -352 488 -306 500
rect -352 -488 -346 488
rect -312 -488 -306 488
rect -352 -500 -306 -488
rect 306 488 352 500
rect 306 -488 312 488
rect 346 -488 352 488
rect 306 -500 352 -488
rect 964 488 1010 500
rect 964 -488 970 488
rect 1004 -488 1010 488
rect 964 -500 1010 -488
rect -954 -547 -362 -541
rect -954 -581 -942 -547
rect -374 -581 -362 -547
rect -954 -587 -362 -581
rect -296 -547 296 -541
rect -296 -581 -284 -547
rect 284 -581 296 -547
rect -296 -587 296 -581
rect 362 -547 954 -541
rect 362 -581 374 -547
rect 942 -581 954 -547
rect 362 -587 954 -581
<< labels >>
rlabel poly -958 500 -358 547 1 G
rlabel locali -346 488 -312 504 1 S
rlabel locali -1004 488 -970 504 1 D
rlabel nsubdiffcont -1118 -587 -1084 587 1 B
<< properties >>
string FIXED_BBOX -1101 -666 1101 666
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 5.0 l 3.0 m 1 nf 3 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
