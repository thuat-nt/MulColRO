magic
tech sky130A
timestamp 1698140848
<< metal4 >>
rect 37444 386004 38883 405005
rect 37444 384883 37557 386004
rect 38764 384883 38883 386004
rect 37444 384753 38883 384883
rect 63390 398361 66908 400977
rect 63390 396027 63606 398361
rect 66692 396027 66908 398361
rect 63390 383496 66908 396027
rect 76674 386046 78113 405046
rect 76674 384925 76768 386046
rect 77975 384925 78113 386046
rect 76674 384794 78113 384925
rect 102608 398450 106126 400972
rect 102608 396116 102862 398450
rect 105948 396116 106126 398450
rect 63390 381162 63606 383496
rect 66692 381162 66908 383496
rect 63390 380912 66908 381162
rect 102608 383518 106126 396116
rect 114584 386313 116023 405345
rect 114584 385192 114661 386313
rect 115868 385192 116023 386313
rect 114584 385093 116023 385192
rect 140445 398523 143963 401515
rect 140445 396189 140726 398523
rect 143812 396189 143963 398523
rect 102608 381184 102831 383518
rect 105917 381184 106126 383518
rect 140445 383896 143963 396189
rect 153451 386611 154890 405525
rect 153451 385490 153587 386611
rect 154794 385490 154890 386611
rect 153451 385273 154890 385490
rect 179417 398458 182935 401488
rect 179417 396124 179657 398458
rect 182743 396124 182935 398458
rect 140445 381562 140677 383896
rect 143763 381562 143963 383896
rect 140445 381450 143963 381562
rect 179417 384020 182935 396124
rect 179417 381686 179656 384020
rect 182742 381686 182935 384020
rect 179417 381423 182935 381686
rect 102608 380907 106126 381184
rect 37855 323770 39216 323940
rect 37855 322844 38034 323770
rect 39076 322844 39216 323770
rect 37855 320080 39216 322844
rect 37855 319542 38087 320080
rect 38983 319542 39216 320080
rect 37855 319220 39216 319542
rect 40095 323794 41301 323986
rect 40095 322942 40270 323794
rect 41159 322942 41301 323794
rect 40095 318344 41301 322942
rect 40095 317866 40251 318344
rect 41080 317866 41301 318344
rect 40095 317470 41301 317866
rect 42148 323798 43578 324142
rect 42148 323032 42381 323798
rect 43363 323032 43578 323798
rect 42148 316711 43578 323032
rect 42148 316172 42379 316711
rect 43298 316172 43578 316711
rect 42148 315777 43578 316172
rect 44462 323927 45830 324160
rect 44462 323026 44568 323927
rect 45643 323026 45830 323927
rect 44462 314950 45830 323026
rect 44462 314364 44738 314950
rect 45654 314364 45830 314950
rect 44462 313966 45830 314364
rect 46591 323944 48075 324162
rect 46591 322991 46799 323944
rect 47805 322991 48075 323944
rect 46591 313156 48075 322991
rect 46591 312524 46789 313156
rect 47763 312524 48075 313156
rect 46591 312248 48075 312524
rect 48886 311415 50208 324679
rect 48886 310813 48994 311415
rect 50039 310813 50208 311415
rect 48886 310492 50208 310813
rect 51087 309652 52388 324875
rect 51087 308894 51195 309652
rect 52269 308894 52388 309652
rect 51087 308728 52388 308894
rect 53177 307847 54515 324723
rect 53177 307146 53340 307847
rect 54333 307146 54515 307847
rect 53177 307013 54515 307146
rect 55265 324012 56638 324755
rect 55265 323020 55434 324012
rect 56426 323020 56638 324012
rect 55265 305994 56638 323020
rect 55265 305325 55424 305994
rect 56440 305325 56638 305994
rect 55265 305114 56638 305325
rect 57385 323867 58756 324198
rect 57385 323099 57526 323867
rect 58627 323099 58756 323867
rect 57385 304023 58756 323099
rect 59455 324021 60892 324246
rect 59455 323044 59607 324021
rect 60729 323044 60892 324021
rect 59455 321960 60892 323044
rect 57385 303228 57572 304023
rect 58660 303228 58756 304023
rect 57385 303111 58756 303228
rect 59447 312937 60892 321960
rect 61675 324030 63070 324194
rect 61675 323053 61824 324030
rect 62946 323053 63070 324030
rect 59447 300083 60876 312937
rect 61675 302251 63070 323053
rect 77047 323761 78408 323963
rect 77047 322835 77229 323761
rect 78271 322835 78408 323761
rect 77047 320160 78408 322835
rect 77047 319622 77245 320160
rect 78141 319622 78408 320160
rect 77047 319243 78408 319622
rect 79332 323849 80538 324082
rect 79332 322997 79487 323849
rect 80376 322997 80538 323849
rect 79332 318408 80538 322997
rect 79332 317930 79544 318408
rect 80373 317930 80538 318408
rect 79332 317566 80538 317930
rect 81401 323837 82831 324141
rect 81401 323071 81612 323837
rect 82594 323071 82831 323837
rect 81401 316751 82831 323071
rect 81401 316212 81679 316751
rect 82598 316212 82831 316751
rect 81401 315776 82831 316212
rect 83665 323927 85033 324140
rect 83665 323026 83783 323927
rect 84858 323026 85033 323927
rect 83665 314903 85033 323026
rect 83665 314317 83899 314903
rect 84815 314317 85033 314903
rect 83665 313946 85033 314317
rect 85787 324043 87271 324123
rect 85787 323090 86010 324043
rect 87016 323090 87271 324043
rect 85787 313196 87271 323090
rect 85787 312564 86011 313196
rect 86985 312564 87271 313196
rect 85787 312209 87271 312564
rect 88144 311411 89466 324660
rect 88144 310809 88283 311411
rect 89328 310809 89466 311411
rect 88144 310473 89466 310809
rect 90298 309671 91599 324756
rect 90298 308913 90438 309671
rect 91512 308913 91599 309671
rect 90298 308729 91599 308913
rect 92426 307919 93764 324687
rect 92426 307218 92608 307919
rect 93601 307218 93764 307919
rect 92426 306977 93764 307218
rect 94528 324099 95901 324777
rect 94528 323107 94710 324099
rect 95702 323107 95901 324099
rect 94528 306028 95901 323107
rect 94528 305359 94675 306028
rect 95691 305359 95901 306028
rect 94528 305136 95901 305359
rect 96602 323941 97979 324254
rect 96602 323173 96755 323941
rect 97856 323173 97979 323941
rect 96602 304009 97979 323173
rect 98643 324068 100080 324329
rect 98643 323129 98945 324068
rect 99912 323129 100080 324068
rect 98643 313020 100080 323129
rect 100891 324098 102287 324239
rect 100891 323046 100983 324098
rect 102204 323046 102287 324098
rect 96602 303241 96749 304009
rect 97850 303241 97979 304009
rect 96602 303111 97979 303241
rect 61675 301369 61817 302251
rect 62972 301369 63070 302251
rect 61675 301313 63070 301369
rect 98645 300221 100074 313020
rect 100891 302220 102287 323046
rect 114872 324037 116233 324138
rect 114872 323111 114991 324037
rect 116033 323111 116233 324037
rect 114872 320169 116233 323111
rect 114872 319631 115077 320169
rect 115973 319631 116233 320169
rect 114872 319418 116233 319631
rect 117145 324096 118351 324245
rect 117145 323244 117330 324096
rect 118219 323244 118351 324096
rect 117145 318436 118351 323244
rect 117145 317958 117327 318436
rect 118156 317958 118351 318436
rect 117145 317729 118351 317958
rect 119243 324073 120673 324354
rect 119243 323307 119508 324073
rect 120490 323307 120673 324073
rect 119243 316751 120673 323307
rect 119243 316212 119520 316751
rect 120439 316212 120673 316751
rect 119243 315989 120673 316212
rect 121499 324176 122867 324405
rect 121499 323275 121624 324176
rect 122699 323275 122867 324176
rect 121499 314962 122867 323275
rect 121499 314376 121739 314962
rect 122655 314376 122867 314962
rect 121499 314211 122867 314376
rect 123629 324275 125113 324335
rect 123629 323322 123897 324275
rect 124903 323322 125113 324275
rect 123629 313172 125113 323322
rect 123629 312540 123895 313172
rect 124869 312540 125113 313172
rect 123629 312421 125113 312540
rect 125962 311426 127284 324679
rect 125962 310824 126123 311426
rect 127168 310824 127284 311426
rect 125962 310492 127284 310824
rect 128125 309662 129426 324756
rect 128125 308904 128218 309662
rect 129292 308904 129426 309662
rect 128125 308718 129426 308904
rect 130274 307905 131612 324710
rect 130274 307204 130464 307905
rect 131457 307204 131612 307905
rect 130274 307000 131612 307204
rect 132282 324332 133655 324879
rect 175465 324739 176902 324879
rect 132282 323340 132542 324332
rect 133534 323340 133655 324332
rect 132282 306057 133655 323340
rect 132282 305388 132446 306057
rect 133462 305388 133655 306057
rect 132282 305238 133655 305388
rect 134447 324343 135823 324525
rect 134447 323366 134594 324343
rect 135706 323366 135823 324343
rect 134447 304059 135823 323366
rect 136536 324409 137973 324553
rect 136536 323315 136634 324409
rect 137879 323315 137973 324409
rect 136536 321844 137973 323315
rect 138731 324378 140131 324523
rect 138731 323284 138808 324378
rect 140053 323284 140131 324378
rect 136536 313244 137985 321844
rect 134447 303175 134595 304059
rect 135694 303175 135823 304059
rect 134447 303112 135823 303175
rect 100891 301404 101004 302220
rect 102174 301404 102287 302220
rect 100891 301312 102287 301404
rect 136556 299967 137985 313244
rect 138731 302211 140131 323284
rect 175465 323608 175591 324739
rect 176823 323608 176902 324739
rect 175465 322129 176902 323608
rect 138731 301409 138837 302211
rect 140038 301409 140131 302211
rect 138731 301312 140131 301409
rect 175453 313570 176902 322129
rect 175453 300252 176882 313570
<< via4 >>
rect 37557 384883 38764 386004
rect 63606 396027 66692 398361
rect 76768 384925 77975 386046
rect 102862 396116 105948 398450
rect 63606 381162 66692 383496
rect 114661 385192 115868 386313
rect 140726 396189 143812 398523
rect 102831 381184 105917 383518
rect 153587 385490 154794 386611
rect 179657 396124 182743 398458
rect 140677 381562 143763 383896
rect 179656 381686 182742 384020
rect 38034 322844 39076 323770
rect 38087 319542 38983 320080
rect 40270 322942 41159 323794
rect 40251 317866 41080 318344
rect 42381 323032 43363 323798
rect 42379 316172 43298 316711
rect 44568 323026 45643 323927
rect 44738 314364 45654 314950
rect 46799 322991 47805 323944
rect 46789 312524 47763 313156
rect 48994 310813 50039 311415
rect 51195 308894 52269 309652
rect 53340 307146 54333 307847
rect 55434 323020 56426 324012
rect 55424 305325 56440 305994
rect 57526 323099 58627 323867
rect 59607 323044 60729 324021
rect 57572 303228 58660 304023
rect 61824 323053 62946 324030
rect 77229 322835 78271 323761
rect 77245 319622 78141 320160
rect 79487 322997 80376 323849
rect 79544 317930 80373 318408
rect 81612 323071 82594 323837
rect 81679 316212 82598 316751
rect 83783 323026 84858 323927
rect 83899 314317 84815 314903
rect 86010 323090 87016 324043
rect 86011 312564 86985 313196
rect 88283 310809 89328 311411
rect 90438 308913 91512 309671
rect 92608 307218 93601 307919
rect 94710 323107 95702 324099
rect 94675 305359 95691 306028
rect 96755 323173 97856 323941
rect 98945 323129 99912 324068
rect 100983 323046 102204 324098
rect 96749 303241 97850 304009
rect 61817 301369 62972 302251
rect 114991 323111 116033 324037
rect 115077 319631 115973 320169
rect 117330 323244 118219 324096
rect 117327 317958 118156 318436
rect 119508 323307 120490 324073
rect 119520 316212 120439 316751
rect 121624 323275 122699 324176
rect 121739 314376 122655 314962
rect 123897 323322 124903 324275
rect 123895 312540 124869 313172
rect 126123 310824 127168 311426
rect 128218 308904 129292 309662
rect 130464 307204 131457 307905
rect 132542 323340 133534 324332
rect 132446 305388 133462 306057
rect 134594 323366 135706 324343
rect 136634 323315 137879 324409
rect 138808 323284 140053 324378
rect 134595 303175 135694 304059
rect 101004 301404 102174 302220
rect 175591 323608 176823 324739
rect 138837 301409 140038 302211
<< metal5 >>
rect 31093 398523 183995 402258
rect 31093 398450 140726 398523
rect 31093 398361 102862 398450
rect 31093 396027 63606 398361
rect 66692 396116 102862 398361
rect 105948 396189 140726 398450
rect 143812 398458 183995 398523
rect 143812 396189 179657 398458
rect 105948 396124 179657 396189
rect 182743 396124 183995 398458
rect 105948 396116 183995 396124
rect 66692 396027 183995 396116
rect 31093 395870 183995 396027
rect 31084 387420 183986 393808
rect 31433 380262 34973 387420
rect 70631 380262 74171 387420
rect 108484 379829 112024 387420
rect 147436 380349 150976 387420
rect 35626 322075 37066 323908
rect 74893 322075 76333 324043
rect 112705 322075 114145 324077
rect 151735 322075 153175 324483
rect 35607 321674 153175 322075
rect 35607 321065 153155 321674
rect 153857 320397 155218 324244
rect 153857 320230 155206 320397
rect 37855 320218 155206 320230
rect 35589 320169 155206 320218
rect 35589 320160 115077 320169
rect 35589 320080 77245 320160
rect 35589 319542 38087 320080
rect 38983 319622 77245 320080
rect 78141 319631 115077 320160
rect 115973 319631 155206 320169
rect 78141 319622 155206 319631
rect 38983 319542 155206 319622
rect 35589 319220 155206 319542
rect 35589 319208 73851 319220
rect 156152 318712 157358 324263
rect 156152 318480 157352 318712
rect 35620 318436 157352 318480
rect 35620 318408 117327 318436
rect 35620 318344 79544 318408
rect 35620 317866 40251 318344
rect 41080 317930 79544 318344
rect 80373 317958 117327 318408
rect 118156 317958 157352 318436
rect 80373 317930 157352 317958
rect 41080 317866 157352 317930
rect 35620 317470 157352 317866
rect 35714 316787 74095 316803
rect 158285 316787 159715 324335
rect 35714 316751 159715 316787
rect 35714 316711 81679 316751
rect 35714 316172 42379 316711
rect 43298 316212 81679 316711
rect 82598 316212 119520 316751
rect 120439 316212 159715 316751
rect 43298 316172 159715 316212
rect 35714 315970 159715 316172
rect 35714 315793 159696 315970
rect 42148 315777 159696 315793
rect 160441 315033 161836 324723
rect 44539 314989 161876 315033
rect 35747 314962 161876 314989
rect 35747 314950 121739 314962
rect 35747 314364 44738 314950
rect 45654 314903 121739 314950
rect 45654 314364 83899 314903
rect 35747 314317 83899 314364
rect 84815 314376 121739 314903
rect 122655 314376 161876 314962
rect 84815 314317 161876 314376
rect 35747 314023 161876 314317
rect 35747 313979 73992 314023
rect 162633 313210 164117 324335
rect 46531 313196 164117 313210
rect 46531 313176 86011 313196
rect 35747 313156 86011 313176
rect 35747 312524 46789 313156
rect 47763 312564 86011 313156
rect 86985 313172 164117 313196
rect 86985 312564 123895 313172
rect 47763 312540 123895 312564
rect 124869 312540 164117 313172
rect 47763 312524 164117 312540
rect 35747 312421 164117 312524
rect 35747 312200 164079 312421
rect 35747 312166 73995 312200
rect 35714 311505 73958 311521
rect 164908 311505 166230 324718
rect 35714 311426 166247 311505
rect 35714 311415 126123 311426
rect 35714 310813 48994 311415
rect 50039 311411 126123 311415
rect 50039 310813 88283 311411
rect 35714 310809 88283 310813
rect 89328 310824 126123 311411
rect 127168 310824 166247 311426
rect 89328 310809 166247 310824
rect 35714 310511 166247 310809
rect 48865 310495 166247 310511
rect 167116 309750 168417 324882
rect 51043 309722 168454 309750
rect 35713 309671 168454 309722
rect 35713 309652 90438 309671
rect 35713 308894 51195 309652
rect 52269 308913 90438 309652
rect 91512 309662 168454 309671
rect 91512 308913 128218 309662
rect 52269 308904 128218 308913
rect 129292 308904 168454 309662
rect 52269 308894 168454 308904
rect 35713 308740 168454 308894
rect 35713 308712 73882 308740
rect 167116 308735 168417 308740
rect 169219 308318 170557 324686
rect 169219 308007 170536 308318
rect 53165 307979 170536 308007
rect 35699 307919 170536 307979
rect 35699 307847 92608 307919
rect 35699 307146 53340 307847
rect 54333 307218 92608 307847
rect 93601 307905 170536 307919
rect 93601 307218 130464 307905
rect 54333 307204 130464 307218
rect 131457 307204 170536 307905
rect 54333 307146 170536 307204
rect 35699 306997 170536 307146
rect 35699 306969 73974 306997
rect 169219 306976 170536 306997
rect 35733 306155 73968 306159
rect 171310 306155 172683 324832
rect 35733 306057 172699 306155
rect 35733 306028 132446 306057
rect 35733 305994 94675 306028
rect 35733 305325 55424 305994
rect 56440 305359 94675 305994
rect 95691 305388 132446 306028
rect 133462 305388 172699 306057
rect 95691 305359 172699 305388
rect 56440 305325 172699 305359
rect 35733 305149 172699 305325
rect 55284 305145 172699 305149
rect 173391 304122 174784 324796
rect 57386 304107 174784 304122
rect 35733 304059 174784 304107
rect 35733 304023 134595 304059
rect 35733 303228 57572 304023
rect 58660 304009 134595 304023
rect 58660 303241 96749 304009
rect 97850 303241 134595 304009
rect 58660 303228 134595 303241
rect 35733 303175 134595 303228
rect 135694 303175 174784 304059
rect 35733 303112 174784 303175
rect 35733 303097 73822 303112
rect 173391 303105 174784 303112
rect 35799 302323 73831 302385
rect 177693 302323 179092 324803
rect 35799 302251 179094 302323
rect 35799 301375 61817 302251
rect 61654 301369 61817 301375
rect 62972 302220 179094 302251
rect 62972 301404 101004 302220
rect 102174 302211 179094 302220
rect 102174 301409 138837 302211
rect 140038 301409 179094 302211
rect 102174 301404 179094 301409
rect 62972 301369 179094 301404
rect 61654 301313 179094 301369
use ColROs  MulColROs[0]
timestamp 1698140848
transform 0 1 156602 1 0 318713
box 4511 -9280 67981 26370
use ColROs  MulColROs[1]
timestamp 1698140848
transform 0 1 117643 1 0 318433
box 4511 -9280 67981 26370
use ColROs  MulColROs[2]
timestamp 1698140848
transform 0 1 79800 1 0 318148
box 4511 -9280 67981 26370
use ColROs  MulColROs[3]
timestamp 1698140848
transform 0 1 40581 1 0 318102
box 4511 -9280 67981 26370
<< labels >>
rlabel metal5 31084 387420 183986 393808 1 VSS
port 1 nsew
rlabel metal5 31093 395870 183995 402258 1 VDD
port 2 nsew
rlabel metal4 37444 384753 38883 405005 1 AOut3
port 3 nsew
rlabel metal4 76674 384794 78113 405046 1 AOut2
port 4 nsew
rlabel metal4 114584 385093 116023 405345 1 AOut1
port 5 nsew
rlabel metal4 153451 385273 154890 405525 1 AOut0
port 6 nsew
rlabel metal5 35607 321065 153155 322075 1 REG6
port 7 nsew
rlabel metal5 35589 319208 73851 320218 1 REG5
port 8 nsew
rlabel metal5 35620 317470 74084 318480 1 REG4
port 9 nsew
rlabel metal5 35714 315793 74095 316803 1 REG3
port 10 nsew
rlabel metal5 35747 313979 73992 314989 1 REG2
port 11 nsew
rlabel metal5 35747 312166 73995 313176 1 REG1
port 12 nsew
rlabel metal5 35714 310511 73958 311521 1 REG0
port 13 nsew
rlabel metal5 35713 308712 73882 309722 1 AIn5
port 14 nsew
rlabel metal5 35699 306969 73974 307979 1 AIn4
port 15 nsew
rlabel metal5 35733 305149 73968 306159 1 AIn3
port 16 nsew
rlabel metal5 35733 303097 73822 304107 1 AIn2
port 17 nsew
rlabel metal5 35799 301375 73831 302385 1 AIn0
port 18 nsew
rlabel metal4 59447 300083 60876 321960 1 AIn_3
port 19 nsew
rlabel metal4 98645 300221 100074 322098 1 AIn_2
port 20 nsew
rlabel metal4 136556 299967 137985 321844 1 AIn_1
port 21 nsew
rlabel metal4 175453 300252 176882 322129 1 AIn_0
port 22 nsew
<< end >>
