magic
tech sky130A
magscale 1 2
timestamp 1695461801
<< error_s >>
rect 6494 7798 6528 8530
rect 7266 7892 7300 7926
rect 7924 7892 7958 7926
rect 9096 7894 9106 7948
rect 9212 7894 9220 7928
rect 9844 7894 9878 7928
rect 10502 7894 10536 7928
rect 11160 7894 11194 7928
rect 11274 7894 11308 8536
rect 7046 7858 8624 7892
rect 6494 7356 6538 7798
rect 6504 7076 6538 7356
rect 7046 7294 7080 7858
rect 7182 7722 7206 7824
rect 7266 7806 7313 7837
rect 7210 7790 7234 7796
rect 7254 7790 7313 7806
rect 7790 7790 7837 7837
rect 7210 7756 7837 7790
rect 7210 7750 7234 7756
rect 7254 7709 7312 7756
rect 7840 7722 7858 7824
rect 7924 7806 7971 7837
rect 7868 7790 7886 7796
rect 7912 7790 7971 7806
rect 8448 7790 8495 7837
rect 8590 7830 8624 7858
rect 8556 7796 8624 7830
rect 9150 7838 9160 7894
rect 9174 7860 12606 7894
rect 9174 7838 9184 7860
rect 7868 7756 8495 7790
rect 7868 7754 7886 7756
rect 7912 7754 7970 7756
rect 7868 7750 7970 7754
rect 7912 7726 7970 7750
rect 7888 7722 7970 7726
rect 7149 7697 7194 7708
rect 7160 7443 7194 7697
rect 7266 7455 7300 7709
rect 7807 7697 7852 7708
rect 7818 7443 7852 7697
rect 7860 7528 7882 7704
rect 7888 7500 7910 7722
rect 7912 7709 7970 7722
rect 7924 7455 7958 7709
rect 8465 7697 8510 7708
rect 8476 7443 8510 7697
rect 8590 7489 8650 7796
rect 8582 7455 8650 7489
rect 7148 7396 7207 7443
rect 7238 7402 7285 7443
rect 7230 7396 7285 7402
rect 7806 7396 7865 7443
rect 7896 7402 7943 7443
rect 7884 7396 7943 7402
rect 8464 7396 8522 7443
rect 7148 7362 7285 7396
rect 7328 7362 7943 7396
rect 7986 7362 8522 7396
rect 8556 7362 8570 7396
rect 7148 7346 7206 7362
rect 7230 7356 7250 7362
rect 7148 7331 7163 7346
rect 7258 7328 7278 7362
rect 7806 7346 7864 7362
rect 7884 7356 7908 7362
rect 7912 7328 7936 7362
rect 8464 7346 8522 7362
rect 8507 7331 8522 7346
rect 8590 7294 8624 7455
rect 9150 7300 9184 7838
rect 9186 7445 9218 7838
rect 9844 7808 9891 7839
rect 9832 7792 9891 7808
rect 9894 7792 9941 7839
rect 10502 7808 10549 7839
rect 10490 7792 10549 7808
rect 10552 7792 10599 7839
rect 11160 7808 11206 7839
rect 11148 7792 11206 7808
rect 11274 7792 11308 7860
rect 9326 7758 9941 7792
rect 9984 7758 10599 7792
rect 10642 7758 11206 7792
rect 11210 7758 11228 7792
rect 9230 7710 9254 7739
rect 9832 7711 9890 7758
rect 10490 7752 10564 7758
rect 10490 7732 10548 7752
rect 10490 7724 10574 7732
rect 10490 7711 10548 7724
rect 11148 7722 11206 7758
rect 11274 7733 11280 7765
rect 11284 7733 11308 7792
rect 11148 7711 11228 7722
rect 9258 7710 9282 7711
rect 9230 7699 9298 7710
rect 9230 7456 9254 7699
rect 9258 7449 9298 7699
rect 9844 7492 9884 7711
rect 9911 7706 9956 7710
rect 9894 7699 9956 7706
rect 9894 7520 9912 7699
rect 9844 7461 9878 7492
rect 9922 7449 9956 7699
rect 10502 7461 10536 7711
rect 10569 7699 10614 7710
rect 10580 7449 10614 7699
rect 11160 7472 11200 7711
rect 11204 7500 11228 7711
rect 11160 7461 11194 7472
rect 9252 7402 9311 7449
rect 9816 7402 9863 7449
rect 9910 7402 9969 7449
rect 10474 7402 10521 7449
rect 10568 7402 10627 7449
rect 11132 7402 11179 7449
rect 9252 7368 9863 7402
rect 9906 7368 10521 7402
rect 10564 7368 11179 7402
rect 9252 7352 9310 7368
rect 9910 7352 9968 7368
rect 10568 7352 10626 7368
rect 9252 7337 9267 7352
rect 11238 7300 11246 7334
rect 11274 7300 11308 7733
rect 6590 7260 8634 7294
rect 9150 7266 11308 7300
rect 7046 7156 7080 7260
rect 6940 7136 7602 7156
rect 6982 7116 7548 7136
rect 7046 7112 7080 7116
rect 7010 7088 7548 7112
rect 7046 7076 7080 7088
rect 8590 7076 8624 7260
rect 9150 7084 9184 7266
rect 6482 6492 6574 7076
rect 7010 6680 7474 7076
rect 7010 6490 7488 6680
rect 7492 6628 7548 6646
rect 7602 6628 7654 6646
rect 7450 6048 7488 6490
rect 7510 6108 7548 6620
rect 7602 6600 7626 6618
rect 7672 6490 8660 7076
rect 9114 5064 9974 7084
rect 10150 5072 11142 7092
rect 11310 6862 12738 7096
rect 11310 6534 12760 6862
rect 9290 4894 9304 5064
rect 9318 4922 9332 5064
rect 8648 3556 8674 4480
rect 8682 3556 8708 4446
rect 10580 3723 10614 5072
rect 11284 3630 11300 3664
rect 11310 3492 12738 6534
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
use opamp  opamp_0
timestamp 1695461801
transform 1 0 -6068 0 1 -644
box 0 -1200 19288 9014
use opamp  x1
timestamp 1695461801
transform 1 0 0 0 1 1800
box 0 -1200 19288 9014
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 opbias
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 in
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 out
port 2 nsew
<< end >>
