magic
tech sky130A
timestamp 1695441144
<< pwell >>
rect -248 -355 248 355
<< nmoslvt >>
rect -150 -250 150 250
<< ndiff >>
rect -179 244 -150 250
rect -179 -244 -173 244
rect -156 -244 -150 244
rect -179 -250 -150 -244
rect 150 244 179 250
rect 150 -244 156 244
rect 173 -244 179 244
rect 150 -250 179 -244
<< ndiffc >>
rect -173 -244 -156 244
rect 156 -244 173 244
<< psubdiff >>
rect -230 320 -182 337
rect 182 320 230 337
rect -230 289 -213 320
rect 213 289 230 320
rect -230 -320 -213 -289
rect 213 -320 230 -289
rect -230 -337 -182 -320
rect 182 -337 230 -320
<< psubdiffcont >>
rect -182 320 182 337
rect -230 -289 -213 289
rect 213 -289 230 289
rect -182 -337 182 -320
<< poly >>
rect -150 286 150 294
rect -150 269 -142 286
rect 142 269 150 286
rect -150 250 150 269
rect -150 -269 150 -250
rect -150 -286 -142 -269
rect 142 -286 150 -269
rect -150 -294 150 -286
<< polycont >>
rect -142 269 142 286
rect -142 -286 142 -269
<< locali >>
rect -230 320 -182 337
rect 182 320 230 337
rect -230 289 -213 320
rect 213 289 230 320
rect -150 269 -142 286
rect 142 269 150 286
rect -173 244 -156 252
rect -173 -252 -156 -244
rect 156 244 173 252
rect 156 -252 173 -244
rect -150 -286 -142 -269
rect 142 -286 150 -269
rect -230 -320 -213 -289
rect 213 -320 230 -289
rect -230 -337 -182 -320
rect 182 -337 230 -320
<< viali >>
rect -142 269 142 286
rect -173 -244 -156 244
rect 156 -244 173 244
rect -142 -286 142 -269
<< metal1 >>
rect -148 286 148 289
rect -148 269 -142 286
rect 142 269 148 286
rect -148 266 148 269
rect -176 244 -153 250
rect -176 -244 -173 244
rect -156 -244 -153 244
rect -176 -250 -153 -244
rect 153 244 176 250
rect 153 -244 156 244
rect 173 -244 176 244
rect 153 -250 176 -244
rect -148 -269 148 -266
rect -148 -286 -142 -269
rect 142 -286 148 -269
rect -148 -289 148 -286
<< labels >>
rlabel psubdiffcont -182 -337 182 -320 1 B
rlabel poly -150 250 150 269 1 G
rlabel locali 156 244 173 252 1 S
rlabel locali -173 244 -156 252 1 D
<< properties >>
string FIXED_BBOX -221 -328 221 328
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 5.0 l 3.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
