magic
tech sky130A
magscale 1 2
timestamp 1696665577
<< locali >>
rect 3474 8344 3884 8346
rect 3474 7934 4444 8344
rect 3474 7762 4214 7934
rect 4388 7762 4444 7934
rect 3474 7238 4444 7762
rect 3474 7216 3884 7238
rect 4214 1828 5094 2332
rect 4214 1654 4258 1828
rect 4422 1654 5094 1828
rect 4214 1220 5094 1654
<< viali >>
rect 4214 7762 4388 7934
rect 4258 1654 4422 1828
<< metal1 >>
rect -40 9086 8604 10274
rect 40 8060 148 8452
rect 40 7406 54 8060
rect 128 7406 148 8060
rect 40 7050 148 7406
rect 190 5046 638 8882
rect 190 4598 292 5046
rect 504 4598 638 5046
rect 190 688 638 4598
rect 848 5054 1296 8898
rect 1348 8060 1456 8464
rect 1348 7406 1368 8060
rect 1442 7406 1456 8060
rect 1348 7062 1456 7406
rect 848 4606 968 5054
rect 1180 4606 1296 5054
rect 688 2072 816 2446
rect 688 1616 714 2072
rect 784 1616 816 2072
rect 688 1094 816 1616
rect 848 704 1296 4606
rect 1510 5046 1958 8882
rect 1510 4598 1614 5046
rect 1826 4598 1958 5046
rect 1510 688 1958 4598
rect 2180 5054 2628 8882
rect 2668 8080 2776 8486
rect 2668 7426 2684 8080
rect 2758 7426 2776 8080
rect 2668 7084 2776 7426
rect 2180 4606 2310 5054
rect 2522 4606 2628 5054
rect 1998 2088 2126 2440
rect 1998 1632 2026 2088
rect 2096 1632 2126 2088
rect 1998 1088 2126 1632
rect 2180 688 2628 4606
rect 2832 5054 3280 8882
rect 4202 7934 4402 7948
rect 4202 7762 4214 7934
rect 4388 7762 4402 7934
rect 4202 7748 4402 7762
rect 4802 5398 4940 9086
rect 2832 4606 2956 5054
rect 3168 4606 3280 5054
rect 5300 4928 5748 8890
rect 5782 7838 5918 8204
rect 5782 7380 5800 7838
rect 5892 7380 5918 7838
rect 5782 7100 5918 7380
rect 2832 688 3280 4606
rect 5300 4480 5412 4928
rect 5624 4480 5748 4928
rect 4228 3404 4428 3444
rect 4228 3282 4284 3404
rect 4402 3282 4428 3404
rect 4228 3244 4428 3282
rect 3320 2110 3448 2470
rect 3320 1654 3348 2110
rect 3418 1654 3448 2110
rect 3320 1118 3448 1654
rect 4238 1828 4438 1844
rect 4238 1654 4258 1828
rect 4422 1654 4438 1828
rect 4238 1644 4438 1654
rect 4804 430 4942 4464
rect 5132 2164 5240 2478
rect 5132 1510 5152 2164
rect 5226 1510 5240 2164
rect 5132 1076 5240 1510
rect 5300 696 5748 4480
rect 5952 4924 6400 8894
rect 5952 4476 6078 4924
rect 6290 4476 6400 4924
rect 5952 994 6400 4476
rect 6610 4928 7058 8890
rect 7102 7810 7238 8186
rect 7102 7352 7118 7810
rect 7210 7352 7238 7810
rect 7102 7082 7238 7352
rect 6610 4480 6726 4928
rect 6938 4480 7058 4928
rect 6442 2136 6550 2484
rect 6442 1482 6466 2136
rect 6540 1482 6550 2136
rect 6442 1082 6550 1482
rect 5952 708 6402 994
rect 6610 696 7058 4480
rect 7274 4922 7722 8878
rect 7274 4474 7394 4922
rect 7606 4474 7722 4922
rect 7274 684 7722 4474
rect 7926 4910 8374 8884
rect 8410 7798 8546 8188
rect 8410 7340 8434 7798
rect 8526 7340 8546 7798
rect 8410 7084 8546 7340
rect 7926 4462 8038 4910
rect 8250 4462 8374 4910
rect 7764 2128 7872 2448
rect 7764 1474 7782 2128
rect 7856 1474 7872 2128
rect 7764 1046 7872 1474
rect 7926 690 8374 4462
rect -30 -918 8632 430
<< via1 >>
rect 54 7406 128 8060
rect 292 4598 504 5046
rect 1368 7406 1442 8060
rect 968 4606 1180 5054
rect 714 1616 784 2072
rect 1614 4598 1826 5046
rect 2684 7426 2758 8080
rect 2310 4606 2522 5054
rect 2026 1632 2096 2088
rect 4238 7784 4374 7920
rect 2956 4606 3168 5054
rect 5800 7380 5892 7838
rect 3604 4702 3784 4870
rect 3612 4698 3676 4702
rect 5412 4480 5624 4928
rect 4284 3282 4402 3404
rect 3348 1654 3418 2110
rect 4264 1664 4418 1818
rect 5152 1510 5226 2164
rect 6078 4476 6290 4924
rect 7118 7352 7210 7810
rect 6726 4480 6938 4928
rect 6466 1482 6540 2136
rect 7394 4474 7606 4922
rect 8434 7340 8526 7798
rect 8038 4462 8250 4910
rect 7782 1474 7856 2128
<< metal2 >>
rect 10 8344 3446 8744
rect 5116 8352 8552 8740
rect 3844 8344 8552 8352
rect 10 8080 8552 8344
rect 10 8060 2684 8080
rect 10 7406 54 8060
rect 128 7406 1368 8060
rect 1442 7426 2684 8060
rect 2758 7920 8552 8080
rect 2758 7784 4238 7920
rect 4374 7838 8552 7920
rect 4374 7784 5800 7838
rect 2758 7426 5800 7784
rect 1442 7406 5800 7426
rect 10 7380 5800 7406
rect 5892 7810 8552 7838
rect 5892 7380 7118 7810
rect 10 7352 7118 7380
rect 7210 7798 8552 7810
rect 7210 7352 8434 7798
rect 10 7340 8434 7352
rect 8526 7340 8552 7798
rect 10 7226 8552 7340
rect 10 7218 4188 7226
rect 10 6798 3446 7218
rect 3688 7216 3752 7218
rect 5116 6794 8552 7226
rect 28 5054 3446 5290
rect 28 5046 968 5054
rect 28 4598 292 5046
rect 504 4606 968 5046
rect 1180 5046 2310 5054
rect 1180 4606 1614 5046
rect 504 4598 1614 4606
rect 1826 4606 2310 5046
rect 2522 4606 2956 5054
rect 3168 4900 3446 5054
rect 5126 4928 8544 5168
rect 5126 4914 5412 4928
rect 3168 4870 3818 4900
rect 3168 4702 3604 4870
rect 3784 4702 3818 4870
rect 3168 4698 3612 4702
rect 3676 4698 3818 4702
rect 3168 4650 3818 4698
rect 4744 4684 5412 4914
rect 3168 4606 3446 4650
rect 1826 4598 3446 4606
rect 28 4376 3446 4598
rect 5126 4480 5412 4684
rect 5624 4924 6726 4928
rect 5624 4480 6078 4924
rect 5126 4476 6078 4480
rect 6290 4480 6726 4924
rect 6938 4922 8544 4928
rect 6938 4480 7394 4922
rect 6290 4476 7394 4480
rect 5126 4474 7394 4476
rect 7606 4910 8544 4922
rect 7606 4474 8038 4910
rect 5126 4462 8038 4474
rect 8250 4462 8544 4910
rect 5126 4254 8544 4462
rect 5126 3474 5310 4254
rect 4218 3404 5310 3474
rect 4218 3282 4284 3404
rect 4402 3282 5310 3404
rect 4218 3220 5310 3282
rect 4218 3216 5270 3220
rect 18 2328 3454 2782
rect 5112 2336 8548 2746
rect 3844 2328 8548 2336
rect 18 2164 8548 2328
rect 18 2110 5152 2164
rect 18 2088 3348 2110
rect 18 2072 2026 2088
rect 18 1616 714 2072
rect 784 1632 2026 2072
rect 2096 1654 3348 2088
rect 3418 1818 5152 2110
rect 3418 1664 4264 1818
rect 4418 1664 5152 1818
rect 3418 1654 5152 1664
rect 2096 1632 5152 1654
rect 784 1616 5152 1632
rect 18 1510 5152 1616
rect 5226 2136 8548 2164
rect 5226 1510 6466 2136
rect 18 1482 6466 1510
rect 6540 2128 8548 2136
rect 6540 1482 7782 2128
rect 18 1474 7782 1482
rect 7856 1474 8548 2128
rect 18 1210 8548 1474
rect 18 1202 4066 1210
rect 18 836 3454 1202
rect 3688 1200 3752 1202
rect 5112 808 8548 1210
rect 5112 800 5802 808
rect 6520 800 8548 808
use not  x1
timestamp 1696661316
transform -1 0 5462 0 1 4624
box 472 -578 1868 1036
use sky130_fd_pr__nfet_01v8_lvt_4833E6  XM1 ~/ColRO/mag
timestamp 1696133064
transform 1 0 6830 0 1 4780
box -1812 -4210 1812 4210
use sky130_fd_pr__pfet_01v8_lvt_RMWXAE  XM10 ~/ColRO/mag
timestamp 1696133064
transform 1 0 1735 0 -1 4788
box -1812 -4219 1812 4219
<< labels >>
flabel metal2 4202 7748 4402 7948 0 FreeSans 256 0 0 0 out
port 1 nsew
rlabel via1 4284 3282 4402 3404 1 toggle
port 6 nsew
rlabel metal1 -40 9086 8604 10274 1 VDD
port 4 nsew
flabel metal2 4238 1644 4438 1844 0 FreeSans 256 0 0 0 in
port 2 nsew
rlabel metal1 -30 -918 8632 430 1 GROUND
port 7 nsew
<< end >>
