magic
tech sky130A
magscale 1 2
timestamp 1695698273
<< error_p >>
rect 163778 19434 164168 19468
rect 163778 18936 163812 19434
rect 163992 19366 164039 19413
rect 163954 19332 164039 19366
rect 163881 19273 163926 19284
rect 164009 19273 164054 19284
rect 163892 19097 163926 19273
rect 164020 19097 164054 19273
rect 163992 19038 164039 19085
rect 163954 19004 164039 19038
rect 164134 18936 164168 19434
rect 163778 18902 164168 18936
rect 163760 18232 164182 18852
rect 172116 17882 172128 18164
rect 172150 17916 172162 18138
<< error_s >>
rect 77095 40320 77129 46278
rect 74349 40013 74383 40320
rect 74463 40109 74497 40143
rect 75121 40109 75155 40143
rect 75779 40109 75813 40143
rect 76437 40109 76471 40143
rect 77095 40109 77129 40143
rect 77753 40109 77807 40143
rect 74413 40075 74417 40109
rect 74429 40075 77807 40109
rect 74317 38203 74383 40013
rect 74459 40023 74463 40041
rect 74459 40007 74509 40023
rect 74520 40013 74538 40028
rect 74548 40013 74566 40026
rect 75061 40007 75108 40054
rect 75117 40023 75121 40041
rect 75117 40007 75167 40023
rect 75719 40013 75766 40054
rect 75710 40007 75766 40013
rect 75775 40023 75779 40041
rect 75775 40007 75825 40023
rect 75840 40013 75846 40016
rect 75868 40013 75874 40026
rect 76377 40007 76424 40054
rect 76433 40023 76437 40041
rect 76433 40007 76483 40023
rect 77035 40013 77082 40054
rect 77030 40007 77082 40013
rect 77091 40023 77095 40041
rect 77091 40007 77141 40023
rect 77693 40007 77740 40054
rect 74463 39973 75108 40007
rect 75121 39973 75766 40007
rect 75779 39973 76424 40007
rect 76437 39973 77082 40007
rect 77095 39973 77740 40007
rect 74463 39926 74509 39973
rect 74419 39914 74437 39926
rect 74463 39914 74497 39926
rect 74419 38302 74497 39914
rect 74520 38626 74538 39967
rect 74548 38598 74566 39967
rect 75121 39926 75167 39973
rect 75710 39967 75731 39973
rect 75738 39939 75759 39973
rect 75779 39926 75825 39973
rect 75078 39914 75109 39925
rect 75121 39914 75155 39926
rect 75736 39914 75767 39925
rect 75779 39914 75813 39926
rect 57080 34865 57336 34874
rect 57108 34837 57308 34846
rect 51612 34568 52178 34602
rect 51612 34280 51646 34568
rect 51983 34488 51994 34499
rect 51667 34426 51748 34473
rect 51807 34454 51994 34488
rect 51995 34426 52076 34473
rect 51714 34388 51748 34426
rect 51767 34388 52023 34394
rect 52042 34388 52076 34426
rect 51767 34374 52024 34388
rect 51983 34366 51994 34371
rect 51795 34360 51995 34366
rect 51795 34346 51996 34360
rect 52034 34346 52130 34360
rect 51807 34326 51994 34346
rect 52144 34332 52178 34568
rect 52006 34318 52178 34332
rect 51769 34288 52021 34291
rect 52144 34280 52178 34318
rect 51612 34257 52178 34280
rect 51612 34246 51646 34257
rect 52144 34246 52178 34257
rect 51612 34245 52178 34246
rect 51646 34231 52144 34245
rect 51612 34212 52178 34231
rect 52228 34194 52848 34616
rect 56702 34242 56718 34244
rect 56610 34133 57230 34242
rect 57342 34228 57784 34262
rect 57280 34201 57846 34228
rect 56610 34099 60480 34133
rect 56610 34063 57230 34099
rect 57280 33934 57314 34099
rect 57382 34065 57416 34068
rect 57710 34065 57744 34068
rect 57812 33934 57846 34099
rect 44606 30992 44640 33696
rect 44792 31012 52768 31026
rect 52920 30992 52954 33696
rect 74317 33341 74351 38203
rect 74419 38141 74465 38302
rect 75018 38249 75028 39648
rect 75046 38277 75056 39620
rect 75089 38302 75155 39914
rect 75747 38302 75813 39914
rect 75840 38614 75846 39967
rect 75868 38586 75874 39967
rect 76437 39926 76483 39973
rect 77030 39967 77047 39973
rect 77058 39939 77075 39973
rect 77095 39926 77141 39973
rect 76394 39914 76425 39925
rect 76437 39914 76471 39926
rect 77052 39914 77083 39925
rect 77095 39914 77129 39926
rect 75089 38290 75123 38302
rect 75747 38290 75781 38302
rect 75077 38277 75136 38290
rect 75046 38268 75136 38277
rect 75143 38268 75174 38277
rect 75077 38249 75136 38268
rect 75018 38243 75136 38249
rect 74525 38209 75136 38243
rect 75171 38243 75202 38249
rect 75735 38243 75794 38290
rect 76328 38249 76348 39654
rect 76356 38277 76376 39626
rect 76405 38302 76471 39914
rect 77063 38302 77129 39914
rect 77162 38592 77166 39967
rect 77190 38564 77194 39967
rect 77710 39914 77741 39925
rect 77753 39914 77787 40075
rect 76405 38290 76439 38302
rect 77063 38290 77097 38302
rect 76393 38277 76452 38290
rect 76356 38274 76452 38277
rect 76459 38274 76484 38277
rect 76393 38249 76452 38274
rect 76328 38246 76452 38249
rect 76487 38246 76512 38249
rect 76393 38243 76452 38246
rect 77051 38243 77110 38290
rect 77650 38249 77670 39624
rect 77678 38249 77698 39596
rect 77721 38302 77787 39914
rect 77835 40013 77853 40075
rect 77867 40013 77901 40320
rect 79420 40018 79454 40320
rect 79534 40114 79568 40148
rect 80192 40114 80226 40148
rect 80850 40114 80884 40148
rect 81508 40114 81542 40148
rect 82166 40114 82200 40148
rect 82824 40114 82878 40148
rect 79484 40080 79488 40114
rect 79500 40080 82878 40114
rect 77721 38290 77755 38302
rect 77709 38243 77767 38290
rect 75171 38240 75794 38243
rect 75183 38209 75794 38240
rect 75841 38209 76452 38243
rect 76499 38209 77110 38243
rect 77157 38209 77767 38243
rect 75077 38193 75123 38209
rect 75735 38193 75781 38209
rect 76393 38193 76439 38209
rect 77051 38193 77097 38209
rect 77709 38193 77755 38209
rect 77835 38203 77901 40013
rect 79388 38226 79454 40018
rect 79530 40028 79534 40046
rect 79530 40012 79580 40028
rect 80132 40012 80170 40050
rect 80188 40028 80192 40046
rect 80188 40012 80238 40028
rect 80790 40018 80828 40050
rect 80780 40012 80828 40018
rect 80846 40028 80850 40046
rect 80846 40012 80896 40028
rect 81448 40012 81486 40050
rect 81504 40028 81508 40046
rect 81504 40012 81554 40028
rect 82106 40012 82144 40050
rect 82162 40028 82166 40046
rect 82162 40012 82212 40028
rect 82764 40012 82802 40050
rect 79534 39978 80170 40012
rect 80192 40008 80828 40012
rect 80192 39978 80830 40008
rect 79534 39940 79580 39978
rect 80192 39940 80238 39978
rect 80780 39972 80802 39978
rect 80808 39944 80830 39978
rect 80850 39978 81486 40012
rect 81508 39978 82144 40012
rect 82166 39978 82802 40012
rect 80850 39940 80896 39978
rect 81508 39940 81554 39978
rect 82102 39972 82118 39978
rect 82130 39944 82146 39972
rect 82166 39940 82212 39978
rect 79490 39928 79508 39940
rect 79534 39928 79568 39940
rect 80149 39928 80180 39939
rect 80192 39928 80226 39940
rect 80807 39928 80838 39939
rect 80850 39928 80884 39940
rect 81465 39928 81496 39939
rect 81508 39928 81542 39940
rect 82123 39928 82154 39939
rect 82166 39928 82200 39940
rect 79490 38316 79568 39928
rect 77063 38141 77097 38193
rect 74419 38107 77767 38141
rect 74431 33437 74465 33471
rect 75089 33437 75123 33471
rect 75747 33437 75781 33471
rect 76405 33437 76439 33471
rect 77063 33437 77097 38107
rect 77721 33437 77755 33471
rect 74399 33403 77789 33437
rect 56504 30992 56538 33322
rect 64818 30992 64852 33322
rect 74303 31839 74351 33341
rect 74431 33351 74465 33403
rect 75089 33382 75123 33403
rect 75747 33382 75781 33403
rect 76405 33382 76439 33403
rect 77063 33382 77097 33403
rect 77721 33382 77755 33403
rect 75047 33351 75123 33382
rect 75705 33351 75781 33382
rect 76363 33351 76439 33382
rect 77021 33351 77097 33382
rect 74431 33254 74477 33351
rect 75047 33335 75135 33351
rect 75705 33335 75793 33351
rect 76363 33335 76451 33351
rect 77021 33335 77109 33351
rect 77679 33335 77755 33382
rect 77835 33341 77869 38203
rect 79388 36384 79422 38226
rect 79490 38164 79536 38316
rect 80088 38272 80114 39392
rect 80116 38272 80142 39364
rect 80160 38316 80226 39928
rect 80818 38316 80884 39928
rect 80160 38304 80194 38316
rect 80818 38304 80852 38316
rect 80148 38266 80198 38304
rect 80252 38272 80270 38288
rect 80806 38266 80856 38304
rect 81408 38272 81424 39374
rect 81436 38272 81452 39346
rect 81476 38316 81542 39928
rect 82134 38316 82200 39928
rect 82232 38570 82238 39972
rect 82260 38542 82266 39972
rect 82781 39928 82812 39939
rect 82824 39928 82858 40080
rect 81476 38304 81510 38316
rect 82134 38304 82168 38316
rect 81464 38266 81514 38304
rect 82122 38266 82172 38304
rect 82716 38272 82740 39376
rect 82744 38272 82768 39348
rect 82792 38316 82858 39928
rect 82906 40018 82924 40080
rect 82938 40018 82972 40320
rect 82792 38304 82826 38316
rect 82780 38266 82830 38304
rect 79596 38232 80198 38266
rect 80254 38232 80856 38266
rect 80912 38232 81514 38266
rect 81570 38232 82172 38266
rect 82228 38232 82830 38266
rect 80148 38216 80194 38232
rect 80806 38216 80852 38232
rect 81464 38216 81510 38232
rect 82122 38216 82168 38232
rect 82780 38216 82826 38232
rect 82906 38226 82972 40018
rect 80160 38164 80194 38216
rect 79490 38130 82838 38164
rect 80160 36384 80194 38130
rect 82128 36384 82150 36574
rect 82906 36384 82940 38226
rect 79388 36356 82940 36384
rect 79082 35914 79084 35962
rect 79054 35886 79084 35906
rect 79388 33346 79422 36356
rect 80160 36328 80194 36356
rect 82128 36328 82150 36356
rect 79460 36300 82878 36328
rect 79502 33442 79536 33476
rect 80160 33442 80194 36300
rect 82128 35906 82150 36300
rect 80852 33644 80858 34718
rect 80852 33476 80884 33644
rect 80818 33442 80884 33476
rect 80908 33442 80912 33672
rect 81476 33442 81510 33476
rect 82070 33442 82096 33636
rect 82128 33608 82152 34718
rect 82098 33476 82152 33608
rect 82098 33442 82168 33476
rect 82792 33442 82826 33476
rect 79470 33408 82860 33442
rect 74479 33301 75135 33335
rect 75137 33301 75793 33335
rect 75795 33301 76451 33335
rect 76453 33301 77109 33335
rect 77111 33301 77755 33335
rect 75055 33295 75059 33301
rect 75083 33267 75087 33301
rect 75089 33254 75135 33301
rect 75747 33254 75793 33301
rect 76371 33295 76375 33301
rect 76399 33267 76403 33301
rect 76405 33254 76451 33301
rect 77063 33254 77109 33301
rect 77687 33295 77691 33301
rect 77715 33267 77719 33301
rect 74431 33242 74465 33254
rect 75064 33242 75077 33253
rect 75089 33242 75123 33254
rect 75722 33242 75735 33253
rect 75747 33242 75781 33254
rect 76380 33242 76393 33253
rect 76405 33242 76439 33254
rect 77038 33242 77051 33253
rect 77063 33242 77097 33254
rect 77696 33242 77709 33253
rect 77721 33242 77755 33301
rect 74417 31938 74465 33242
rect 75075 31938 75123 33242
rect 75733 31938 75781 33242
rect 41408 30958 68008 30992
rect 44606 30890 44640 30958
rect 44708 30890 44742 30958
rect 45188 30890 45226 30928
rect 45946 30890 45984 30928
rect 46704 30890 46742 30928
rect 47462 30890 47500 30928
rect 48220 30890 48258 30928
rect 48978 30890 49016 30928
rect 49736 30890 49774 30928
rect 50494 30890 50532 30928
rect 51252 30890 51290 30928
rect 52010 30890 52048 30928
rect 52768 30890 52780 30928
rect 44606 30856 45226 30890
rect 45278 30856 45984 30890
rect 46036 30856 46742 30890
rect 46794 30856 47500 30890
rect 47552 30856 48258 30890
rect 48310 30856 49016 30890
rect 49068 30856 49774 30890
rect 49826 30856 50532 30890
rect 50584 30856 51290 30890
rect 51342 30856 52048 30890
rect 52100 30856 52780 30890
rect 42942 26258 42976 30806
rect 44606 30274 44640 30856
rect 44708 30416 44742 30856
rect 52820 30840 52852 30928
rect 52858 30856 52890 30890
rect 44780 30818 44781 30819
rect 52779 30818 52780 30819
rect 52820 30818 52864 30840
rect 44779 30817 44780 30818
rect 52780 30817 52781 30818
rect 45205 30806 45250 30817
rect 45963 30806 46008 30817
rect 46721 30806 46766 30817
rect 47479 30806 47524 30817
rect 48237 30806 48282 30817
rect 48995 30806 49040 30817
rect 49753 30806 49798 30817
rect 50511 30806 50556 30817
rect 51269 30806 51314 30817
rect 52027 30806 52072 30817
rect 45204 30400 45205 30401
rect 45203 30399 45204 30400
rect 45216 30388 45250 30806
rect 45261 30400 45262 30401
rect 45962 30400 45963 30401
rect 45262 30399 45263 30400
rect 45961 30399 45962 30400
rect 45974 30388 46008 30806
rect 46019 30400 46020 30401
rect 46720 30400 46721 30401
rect 46020 30399 46021 30400
rect 46719 30399 46720 30400
rect 46732 30388 46766 30806
rect 46777 30400 46778 30401
rect 47478 30400 47479 30401
rect 46778 30399 46779 30400
rect 47477 30399 47478 30400
rect 47490 30388 47524 30806
rect 47535 30400 47536 30401
rect 48236 30400 48237 30401
rect 47536 30399 47537 30400
rect 48235 30399 48236 30400
rect 48248 30388 48282 30806
rect 48293 30400 48294 30401
rect 48994 30400 48995 30401
rect 48294 30399 48295 30400
rect 48993 30399 48994 30400
rect 49006 30388 49040 30806
rect 49051 30400 49052 30401
rect 49752 30400 49753 30401
rect 49052 30399 49053 30400
rect 49751 30399 49752 30400
rect 49764 30388 49798 30806
rect 49809 30400 49810 30401
rect 50510 30400 50511 30401
rect 49810 30399 49811 30400
rect 50509 30399 50510 30400
rect 50522 30388 50556 30806
rect 50567 30400 50568 30401
rect 51268 30400 51269 30401
rect 50568 30399 50569 30400
rect 51267 30399 51268 30400
rect 51280 30388 51314 30806
rect 51325 30400 51326 30401
rect 52026 30400 52027 30401
rect 51326 30399 51327 30400
rect 52025 30399 52026 30400
rect 52038 30388 52072 30806
rect 52784 30416 52864 30818
rect 52083 30400 52084 30401
rect 52784 30400 52842 30416
rect 52084 30399 52085 30400
rect 52768 30388 52779 30399
rect 44792 30354 52784 30388
rect 45216 30274 45250 30354
rect 45974 30274 46008 30354
rect 46732 30274 46766 30354
rect 47490 30274 47524 30354
rect 48248 30274 48282 30354
rect 49006 30274 49040 30354
rect 49764 30274 49798 30354
rect 50522 30274 50556 30354
rect 51280 30274 51314 30354
rect 52038 30274 52072 30354
rect 52796 30320 52818 30400
rect 52796 30316 52806 30320
rect 52796 30274 52830 30308
rect 52920 30274 52954 30958
rect 56504 30890 56538 30958
rect 56590 30928 56616 30948
rect 55132 30856 56574 30890
rect 44606 30240 52954 30274
rect 48296 29824 48322 29986
rect 48324 29824 48350 29986
rect 48100 29362 48738 29824
rect 49006 29770 49040 29804
rect 49134 29770 49160 29948
rect 49162 29770 49188 29948
rect 48788 29736 49336 29770
rect 48788 29454 48822 29736
rect 49006 29656 49040 29736
rect 49134 29667 49160 29736
rect 49134 29662 49161 29667
rect 49162 29662 49188 29736
rect 49150 29656 49161 29662
rect 48852 29612 48924 29650
rect 48974 29622 49161 29656
rect 48890 29578 48924 29612
rect 48993 29610 48994 29611
rect 48994 29609 48995 29610
rect 48994 29580 48995 29581
rect 48993 29579 48994 29580
rect 49006 29568 49040 29622
rect 49162 29612 49234 29650
rect 49052 29610 49053 29611
rect 49051 29609 49052 29610
rect 49051 29580 49052 29581
rect 49052 29579 49053 29580
rect 49150 29568 49161 29579
rect 49200 29578 49234 29612
rect 48974 29534 49161 29568
rect 49006 29454 49040 29534
rect 49134 29454 49152 29528
rect 49162 29454 49180 29528
rect 49302 29454 49336 29736
rect 48788 29420 49336 29454
rect 48302 29212 48322 29362
rect 48330 29240 48350 29362
rect 49134 29338 49152 29420
rect 49162 29366 49180 29420
rect 49134 29240 49154 29338
rect 49162 29212 49182 29366
rect 45428 28757 45750 28788
rect 48474 28757 48796 28776
rect 44575 26036 53013 28757
rect 55828 26258 55862 30806
rect 56504 29900 56538 30856
rect 56590 30840 56640 30928
rect 57316 30890 57354 30928
rect 58074 30890 58112 30928
rect 58832 30890 58870 30928
rect 59590 30890 59628 30928
rect 60348 30890 60386 30928
rect 61106 30890 61144 30928
rect 61864 30890 61902 30928
rect 62622 30890 62660 30928
rect 63380 30890 63418 30928
rect 64138 30890 64176 30928
rect 64716 30890 64750 30958
rect 64818 30890 64852 30958
rect 56648 30856 57354 30890
rect 57406 30856 58112 30890
rect 58164 30856 58870 30890
rect 58922 30856 59628 30890
rect 59680 30856 60386 30890
rect 60438 30856 61144 30890
rect 61196 30856 61902 30890
rect 61954 30856 62660 30890
rect 62712 30856 63418 30890
rect 63470 30856 64176 30890
rect 64228 30856 64852 30890
rect 56590 30818 56654 30840
rect 56678 30818 56679 30819
rect 64677 30818 64678 30819
rect 56575 30803 56654 30818
rect 56677 30817 56678 30818
rect 64678 30817 64679 30818
rect 57333 30806 57378 30817
rect 58091 30806 58136 30817
rect 58849 30806 58894 30817
rect 59607 30806 59652 30817
rect 60365 30806 60410 30817
rect 61123 30806 61168 30817
rect 61881 30806 61926 30817
rect 62639 30806 62684 30817
rect 63397 30806 63442 30817
rect 64155 30806 64200 30817
rect 56590 30700 56654 30803
rect 56590 30684 56632 30700
rect 57332 30684 57333 30685
rect 57331 30683 57332 30684
rect 57344 30672 57378 30806
rect 57389 30684 57390 30685
rect 58090 30684 58091 30685
rect 57390 30683 57391 30684
rect 58089 30683 58090 30684
rect 58102 30672 58136 30806
rect 58147 30684 58148 30685
rect 58848 30684 58849 30685
rect 58148 30683 58149 30684
rect 58847 30683 58848 30684
rect 58860 30672 58894 30806
rect 58905 30684 58906 30685
rect 59606 30684 59607 30685
rect 58906 30683 58907 30684
rect 59605 30683 59606 30684
rect 59618 30672 59652 30806
rect 59663 30684 59664 30685
rect 60364 30684 60365 30685
rect 59664 30683 59665 30684
rect 60363 30683 60364 30684
rect 60376 30672 60410 30806
rect 60421 30684 60422 30685
rect 61122 30684 61123 30685
rect 60422 30683 60423 30684
rect 61121 30683 61122 30684
rect 61134 30672 61168 30806
rect 61179 30684 61180 30685
rect 61880 30684 61881 30685
rect 61180 30683 61181 30684
rect 61879 30683 61880 30684
rect 61892 30672 61926 30806
rect 61937 30684 61938 30685
rect 62638 30684 62639 30685
rect 61938 30683 61939 30684
rect 62637 30683 62638 30684
rect 62650 30672 62684 30806
rect 62695 30684 62696 30685
rect 63396 30684 63397 30685
rect 62696 30683 62697 30684
rect 63395 30683 63396 30684
rect 63408 30672 63442 30806
rect 63453 30684 63454 30685
rect 64154 30684 64155 30685
rect 63454 30683 63455 30684
rect 64153 30683 64154 30684
rect 64166 30672 64200 30806
rect 64716 30700 64750 30856
rect 64211 30684 64212 30685
rect 64212 30683 64213 30684
rect 64666 30672 64677 30683
rect 56582 30644 56640 30648
rect 56572 30610 56640 30644
rect 56690 30638 64677 30672
rect 57331 30626 57332 30627
rect 57332 30625 57333 30626
rect 56590 30042 56654 30610
rect 56590 30026 56632 30042
rect 57344 30036 57378 30638
rect 57390 30626 57391 30627
rect 58089 30626 58090 30627
rect 57389 30625 57390 30626
rect 58090 30625 58091 30626
rect 57408 30036 58062 30038
rect 57302 30014 58062 30036
rect 58090 30026 58091 30027
rect 58089 30025 58090 30026
rect 58102 30014 58136 30638
rect 58148 30626 58149 30627
rect 58847 30626 58848 30627
rect 58147 30625 58148 30626
rect 58848 30625 58849 30626
rect 58147 30026 58148 30027
rect 58848 30026 58849 30027
rect 58148 30025 58149 30026
rect 58847 30025 58848 30026
rect 58860 30014 58894 30638
rect 58906 30626 58907 30627
rect 59605 30626 59606 30627
rect 58905 30625 58906 30626
rect 59606 30625 59607 30626
rect 58905 30026 58906 30027
rect 59606 30026 59607 30027
rect 58906 30025 58907 30026
rect 59605 30025 59606 30026
rect 59618 30014 59652 30638
rect 60300 30632 60370 30638
rect 59664 30626 59665 30627
rect 60363 30626 60364 30627
rect 59663 30625 59664 30626
rect 60364 30625 60365 30626
rect 60328 30604 60370 30612
rect 60300 30074 60322 30112
rect 60328 30046 60350 30112
rect 59663 30026 59664 30027
rect 60364 30026 60365 30027
rect 59664 30025 59665 30026
rect 60363 30025 60364 30026
rect 60376 30014 60410 30638
rect 60416 30632 60480 30638
rect 60422 30626 60423 30627
rect 61121 30626 61122 30627
rect 60421 30625 60422 30626
rect 61122 30625 61123 30626
rect 60416 30604 60452 30612
rect 60421 30026 60422 30027
rect 61122 30026 61123 30027
rect 60422 30025 60423 30026
rect 61121 30025 61122 30026
rect 61134 30014 61168 30638
rect 61180 30626 61181 30627
rect 61879 30626 61880 30627
rect 61179 30625 61180 30626
rect 61880 30625 61881 30626
rect 61179 30026 61180 30027
rect 61880 30026 61881 30027
rect 61180 30025 61181 30026
rect 61879 30025 61880 30026
rect 61892 30014 61926 30638
rect 61938 30626 61939 30627
rect 62637 30626 62638 30627
rect 61937 30625 61938 30626
rect 62638 30625 62639 30626
rect 61937 30026 61938 30027
rect 62638 30026 62639 30027
rect 61938 30025 61939 30026
rect 62637 30025 62638 30026
rect 62650 30014 62684 30638
rect 62696 30626 62697 30627
rect 63395 30626 63396 30627
rect 62695 30625 62696 30626
rect 63396 30625 63397 30626
rect 63324 30594 63402 30618
rect 63352 30566 63402 30590
rect 62695 30026 62696 30027
rect 63396 30026 63397 30027
rect 62696 30025 62697 30026
rect 63395 30025 63396 30026
rect 63408 30014 63442 30638
rect 63454 30626 63455 30627
rect 64153 30626 64154 30627
rect 63453 30625 63454 30626
rect 64154 30625 64155 30626
rect 63448 30594 63504 30618
rect 63448 30566 63476 30590
rect 63453 30026 63454 30027
rect 64154 30026 64155 30027
rect 63454 30025 63455 30026
rect 64153 30025 64154 30026
rect 64166 30014 64200 30638
rect 64212 30626 64213 30627
rect 64211 30625 64212 30626
rect 64678 30610 64750 30648
rect 64716 30042 64750 30610
rect 64211 30026 64212 30027
rect 64212 30025 64213 30026
rect 64666 30014 64677 30025
rect 56690 29980 64677 30014
rect 57302 29964 58062 29980
rect 56566 29900 56586 29934
rect 57302 29900 57422 29964
rect 58102 29900 58136 29980
rect 58860 29900 58894 29980
rect 59618 29900 59652 29980
rect 60376 29900 60410 29980
rect 61134 29900 61168 29980
rect 61892 29900 61926 29980
rect 62650 29900 62684 29980
rect 63408 29900 63442 29980
rect 64166 29900 64200 29980
rect 64818 29900 64852 30856
rect 56504 29866 64852 29900
rect 60376 29396 60410 29430
rect 60122 29362 60670 29396
rect 60122 29080 60156 29362
rect 60186 29238 60258 29276
rect 60224 29204 60258 29238
rect 60268 29126 60270 29316
rect 60296 29242 60298 29288
rect 60376 29282 60410 29362
rect 60484 29282 60495 29293
rect 60308 29248 60495 29282
rect 60363 29236 60364 29237
rect 60364 29235 60365 29236
rect 60328 29222 60370 29228
rect 60364 29206 60365 29207
rect 60363 29205 60364 29206
rect 60296 29154 60298 29200
rect 60300 29194 60370 29200
rect 60376 29194 60410 29248
rect 60496 29238 60568 29276
rect 60422 29236 60423 29237
rect 60421 29235 60422 29236
rect 60416 29222 60452 29228
rect 60421 29206 60422 29207
rect 60422 29205 60423 29206
rect 60416 29194 60480 29200
rect 60484 29194 60495 29205
rect 60534 29204 60568 29238
rect 60308 29160 60495 29194
rect 60376 29080 60410 29160
rect 60636 29080 60670 29362
rect 60122 29046 60670 29080
rect 60720 28988 61358 29450
rect 60622 28383 60944 28794
rect 56445 26036 64883 28383
rect 66440 26258 66474 30806
rect 67308 26214 67316 30850
rect 67336 26214 67372 30850
rect 74303 25167 74337 31839
rect 74417 31777 74451 31938
rect 75075 31926 75109 31938
rect 75733 31926 75767 31938
rect 74453 31811 74457 31913
rect 74481 31879 74485 31885
rect 75061 31879 75109 31926
rect 75719 31879 75767 31926
rect 74477 31845 74485 31879
rect 74493 31845 75109 31879
rect 75135 31845 75143 31879
rect 75151 31845 75767 31879
rect 74481 31839 74485 31845
rect 75063 31829 75109 31845
rect 75721 31829 75767 31845
rect 75075 31777 75109 31829
rect 75733 31777 75767 31829
rect 75769 31811 75773 31913
rect 76314 31885 76316 32982
rect 76342 31885 76344 32954
rect 76391 31938 76439 33242
rect 77049 31938 77097 33242
rect 76391 31926 76425 31938
rect 77049 31926 77083 31938
rect 75797 31879 75801 31885
rect 76377 31879 76425 31926
rect 77035 31879 77083 31926
rect 75793 31845 75801 31879
rect 75809 31845 76425 31879
rect 76451 31845 76459 31879
rect 76467 31845 77083 31879
rect 75797 31839 75801 31845
rect 76314 31832 76316 31839
rect 76342 31804 76344 31839
rect 76379 31829 76425 31845
rect 77037 31829 77083 31845
rect 76391 31777 76425 31829
rect 77049 31777 77083 31829
rect 77085 31811 77089 31913
rect 77636 31885 77638 32952
rect 77664 31885 77666 32924
rect 77707 31938 77755 33242
rect 77707 31926 77741 31938
rect 77113 31879 77117 31885
rect 77693 31879 77741 31926
rect 77109 31845 77117 31879
rect 77125 31845 77741 31879
rect 77113 31839 77117 31845
rect 77636 31832 77638 31839
rect 77664 31804 77666 31839
rect 77695 31829 77741 31845
rect 77707 31777 77741 31829
rect 77821 31839 77869 33341
rect 79374 31862 79422 33346
rect 79502 33356 79536 33408
rect 80118 33374 80156 33378
rect 79502 33268 79548 33356
rect 80118 33340 80158 33374
rect 79550 33306 80158 33340
rect 80126 33300 80130 33306
rect 80154 33272 80158 33306
rect 80160 33356 80194 33408
rect 80160 33268 80206 33356
rect 80776 33340 80814 33378
rect 80208 33306 80814 33340
rect 80818 33346 80884 33408
rect 80908 33346 80912 33408
rect 80818 33300 80864 33346
rect 81434 33340 81472 33378
rect 80866 33306 81472 33340
rect 81476 33356 81510 33408
rect 82070 33378 82096 33408
rect 82098 33378 82168 33408
rect 82070 33356 82168 33378
rect 82750 33374 82788 33378
rect 79502 33256 79536 33268
rect 80135 33256 80148 33267
rect 80160 33256 80194 33268
rect 80793 33256 80806 33267
rect 80818 33256 80884 33300
rect 79488 31952 79536 33256
rect 74405 31743 77753 31777
rect 77821 25167 77855 31839
rect 79374 25190 79408 31862
rect 79488 31800 79522 31952
rect 79524 31834 79528 31936
rect 80074 31908 80082 32720
rect 80102 31908 80110 32692
rect 80146 31952 80194 33256
rect 80804 32242 80884 33256
rect 80146 31940 80180 31952
rect 80804 31940 80858 32242
rect 80908 32214 80912 33300
rect 81476 33268 81522 33356
rect 82070 33346 82180 33356
rect 82092 33340 82130 33346
rect 81524 33306 82130 33340
rect 82134 33300 82180 33346
rect 82750 33340 82790 33374
rect 82182 33306 82790 33340
rect 82758 33300 82762 33306
rect 81451 33256 81464 33267
rect 81476 33256 81510 33268
rect 81462 31952 81510 33256
rect 82070 32178 82096 33300
rect 82098 33268 82180 33300
rect 82786 33272 82790 33306
rect 82098 32206 82168 33268
rect 82767 33256 82780 33267
rect 82792 33256 82826 33408
rect 82906 33346 82940 36356
rect 83558 34992 91534 35026
rect 84140 34410 85244 34430
rect 82086 32132 82096 32178
rect 82114 32132 82168 32206
rect 82702 32132 82708 32704
rect 82730 32132 82736 32676
rect 82120 31994 82168 32132
rect 81462 31940 81496 31952
rect 79552 31902 79556 31908
rect 80132 31902 80180 31940
rect 80790 31908 80844 31940
rect 80790 31902 80838 31908
rect 79548 31868 79556 31902
rect 79564 31868 80180 31902
rect 80206 31868 80214 31902
rect 80222 31868 80838 31902
rect 79552 31862 79556 31868
rect 80074 31856 80082 31862
rect 80102 31828 80110 31862
rect 80134 31852 80180 31868
rect 80792 31862 80838 31868
rect 80840 31862 80844 31908
rect 80868 31902 80872 31908
rect 81448 31902 81496 31940
rect 82086 31908 82096 31994
rect 82114 31952 82168 31994
rect 82114 31940 82154 31952
rect 82106 31902 82154 31940
rect 80864 31868 80872 31902
rect 80880 31868 81496 31902
rect 81522 31868 81530 31902
rect 81538 31868 82154 31902
rect 80868 31862 80872 31868
rect 80792 31852 80844 31862
rect 81450 31852 81496 31868
rect 80146 31800 80180 31852
rect 80804 31806 80844 31852
rect 80804 31800 80838 31806
rect 81462 31800 81496 31852
rect 82086 31800 82096 31862
rect 82108 31852 82154 31868
rect 82114 31800 82154 31852
rect 82156 31834 82160 31936
rect 82702 31908 82708 31994
rect 82730 31908 82736 31994
rect 82778 31952 82826 33256
rect 82778 31940 82812 31952
rect 82184 31902 82188 31908
rect 82764 31902 82812 31940
rect 82180 31868 82188 31902
rect 82196 31868 82812 31902
rect 82184 31862 82188 31868
rect 82702 31850 82708 31862
rect 82730 31828 82736 31862
rect 82766 31852 82812 31868
rect 82778 31800 82812 31852
rect 82892 31862 82940 33346
rect 83336 33332 86647 33473
rect 83219 33301 86647 33332
rect 83336 33298 86647 33301
rect 83139 32920 83162 33282
rect 83185 33267 86647 33298
rect 83167 32920 83190 33254
rect 83336 32280 86647 33267
rect 88130 33408 91665 33442
rect 88130 33052 88164 33408
rect 88874 33340 88912 33378
rect 89532 33340 89570 33378
rect 90190 33340 90228 33378
rect 90848 33340 90886 33378
rect 91506 33340 91544 33378
rect 88306 33306 88912 33340
rect 88964 33306 89570 33340
rect 89622 33306 90228 33340
rect 90280 33306 90886 33340
rect 90938 33306 91544 33340
rect 91584 33296 91602 33306
rect 88233 33256 88278 33267
rect 88891 33256 88936 33267
rect 89549 33256 89594 33267
rect 90207 33256 90252 33267
rect 90865 33256 90910 33267
rect 88244 33052 88278 33256
rect 88289 33064 88290 33065
rect 88890 33064 88891 33065
rect 88290 33063 88291 33064
rect 88889 33063 88890 33064
rect 88902 33052 88936 33256
rect 88947 33064 88948 33065
rect 89548 33064 89549 33065
rect 88948 33063 88949 33064
rect 89547 33063 89548 33064
rect 89560 33052 89594 33256
rect 89605 33064 89606 33065
rect 90206 33064 90207 33065
rect 89606 33063 89607 33064
rect 90205 33063 90206 33064
rect 90218 33052 90252 33256
rect 90263 33064 90264 33065
rect 90864 33064 90865 33065
rect 90264 33063 90265 33064
rect 90863 33063 90864 33064
rect 90876 33052 90910 33256
rect 91500 33144 91518 33296
rect 91578 33294 91602 33296
rect 91550 33268 91568 33272
rect 91578 33268 91606 33294
rect 91528 33267 91606 33268
rect 91523 33256 91606 33267
rect 91528 33116 91606 33256
rect 91534 33080 91606 33116
rect 91534 33068 91602 33080
rect 90921 33064 90922 33065
rect 91522 33064 91523 33065
rect 90922 33063 90923 33064
rect 91521 33063 91522 33064
rect 91534 33052 91580 33068
rect 91584 33064 91602 33068
rect 91614 33064 91618 33408
rect 91648 33080 91665 33408
rect 88130 33049 91580 33052
rect 88130 33040 91574 33049
rect 88130 33030 91568 33040
rect 91648 33037 91652 33080
rect 88130 33028 91574 33030
rect 88130 33018 91580 33028
rect 88130 32394 88164 33018
rect 88244 32394 88278 33018
rect 88290 33006 88291 33007
rect 88889 33006 88890 33007
rect 88289 33005 88290 33006
rect 88890 33005 88891 33006
rect 88289 32406 88290 32407
rect 88890 32406 88891 32407
rect 88290 32405 88291 32406
rect 88889 32405 88890 32406
rect 88902 32394 88936 33018
rect 88948 33006 88949 33007
rect 89547 33006 89548 33007
rect 88947 33005 88948 33006
rect 89548 33005 89549 33006
rect 88947 32406 88948 32407
rect 89548 32406 89549 32407
rect 88948 32405 88949 32406
rect 89547 32405 89548 32406
rect 89560 32394 89594 33018
rect 89606 33006 89607 33007
rect 90205 33006 90206 33007
rect 89605 33005 89606 33006
rect 90206 33005 90207 33006
rect 89605 32406 89606 32407
rect 90206 32406 90207 32407
rect 89606 32405 89607 32406
rect 90205 32405 90206 32406
rect 90218 32394 90252 33018
rect 90264 33006 90265 33007
rect 90863 33006 90864 33007
rect 90263 33005 90264 33006
rect 90864 33005 90865 33006
rect 90263 32406 90264 32407
rect 90864 32406 90865 32407
rect 90264 32405 90265 32406
rect 90863 32405 90864 32406
rect 90876 32394 90910 33018
rect 90922 33006 90923 33007
rect 91521 33006 91522 33007
rect 90921 33005 90922 33006
rect 91522 33005 91523 33006
rect 91534 33002 91580 33018
rect 91584 33002 91602 33006
rect 91534 32990 91602 33002
rect 91534 32940 91606 32990
rect 90921 32406 90922 32407
rect 91522 32406 91523 32407
rect 90922 32405 90923 32406
rect 91521 32405 91522 32406
rect 91534 32394 91580 32940
rect 91584 32422 91606 32940
rect 91584 32406 91602 32422
rect 91614 32406 91618 33006
rect 91648 32422 91665 33037
rect 88130 32391 91580 32394
rect 88130 32360 91568 32391
rect 91648 32372 91652 32422
rect 88130 32280 88164 32360
rect 88244 32280 88278 32360
rect 88902 32280 88936 32360
rect 89560 32280 89594 32360
rect 90218 32280 90252 32360
rect 90876 32280 90910 32360
rect 91534 32280 91568 32360
rect 83336 32246 91580 32280
rect 91648 32246 91658 32314
rect 91686 32280 91720 33496
rect 113115 33045 113149 39409
rect 115197 35610 115243 37670
rect 115246 35610 115271 37670
rect 113229 33141 113263 33175
rect 113887 33141 113921 33175
rect 114545 33141 114579 33175
rect 115197 33141 115243 34422
rect 115246 33141 115271 34422
rect 115861 33141 115895 39310
rect 116476 37640 116492 37976
rect 116633 33437 116667 39409
rect 118958 33473 118992 39324
rect 121101 33478 121774 36685
rect 127606 35970 129070 35976
rect 127162 35185 127942 35196
rect 127200 35147 127904 35158
rect 127668 34594 129020 34610
rect 124686 34527 124744 34540
rect 128422 34527 128514 34540
rect 124720 34493 124744 34506
rect 128422 34493 128480 34506
rect 118150 33437 119557 33473
rect 121101 33442 124628 33478
rect 115969 33403 119557 33437
rect 115969 33141 116003 33403
rect 116098 33335 116565 33382
rect 116145 33301 116565 33335
rect 116507 33254 116565 33301
rect 116072 33242 116128 33253
rect 116083 33141 116128 33242
rect 116519 33175 116564 33254
rect 116519 33141 116573 33175
rect 116633 33141 116667 33403
rect 117370 33310 117383 33341
rect 117337 33295 117383 33310
rect 118107 33310 118130 33341
rect 118150 33310 119557 33403
rect 118107 33295 119557 33310
rect 118150 33182 119557 33295
rect 113179 33107 113183 33141
rect 113195 33107 116667 33141
rect 83336 32210 86647 32246
rect 79476 31766 82824 31800
rect 80146 25280 80180 31766
rect 82086 31398 82096 31766
rect 82114 31398 82152 31766
rect 81528 30892 82120 30906
rect 82154 30892 82308 30906
rect 81562 30858 82120 30872
rect 82154 30858 82308 30872
rect 82086 27438 82096 30210
rect 82114 27438 82152 30210
rect 80846 26512 80870 26972
rect 80852 25570 80870 26512
rect 80804 25280 80844 25292
rect 80798 25268 80844 25280
rect 82086 25240 82096 25534
rect 82114 25292 82152 25534
rect 82246 25478 82248 26992
rect 82114 25280 82154 25292
rect 82114 25268 82160 25280
rect 82892 25190 82926 31862
rect 83135 31790 83136 31876
rect 83173 31752 83174 31914
rect 83342 31872 83764 32210
rect 83831 30727 83865 30761
rect 84489 30727 84523 30761
rect 85147 30727 85181 30761
rect 85805 30727 85839 30761
rect 86463 30727 86497 30761
rect 86577 30727 86611 32210
rect 86612 31830 86647 32084
rect 86866 31368 86901 31830
rect 87322 31658 87424 31670
rect 88130 30763 88164 32246
rect 88206 32018 88220 32104
rect 88244 31980 88258 32142
rect 113083 31235 113149 33045
rect 113225 33055 113229 33073
rect 113225 33039 113275 33055
rect 113286 33045 113304 33060
rect 113314 33045 113332 33058
rect 113827 33039 113874 33086
rect 113883 33055 113887 33073
rect 113883 33039 113933 33055
rect 114485 33045 114532 33086
rect 114476 33039 114532 33045
rect 114541 33055 114545 33073
rect 114541 33039 114591 33055
rect 114606 33045 114612 33048
rect 114634 33045 114640 33058
rect 115143 33039 115190 33086
rect 115197 33055 115243 33107
rect 115246 33055 115271 33107
rect 115197 33045 115271 33055
rect 115199 33039 115249 33045
rect 115801 33039 115848 33086
rect 115861 33073 115895 33107
rect 115857 33055 115895 33073
rect 115857 33039 115907 33055
rect 115969 33039 116003 33107
rect 116083 33104 116128 33107
rect 116519 33104 116564 33107
rect 116083 33086 116117 33104
rect 116083 33039 116130 33086
rect 116459 33039 116506 33086
rect 113229 33005 113874 33039
rect 113887 33005 114532 33039
rect 114545 33005 115190 33039
rect 115203 33005 115848 33039
rect 115861 33005 116506 33039
rect 113229 32958 113275 33005
rect 113185 32946 113203 32958
rect 113229 32946 113263 32958
rect 113185 31322 113263 32946
rect 113286 31658 113304 32999
rect 113314 31630 113332 32999
rect 113887 32958 113933 33005
rect 114476 32999 114497 33005
rect 114504 32971 114525 33005
rect 114545 32958 114591 33005
rect 115203 32999 115249 33005
rect 113844 32946 113875 32957
rect 113887 32946 113921 32958
rect 114502 32946 114533 32957
rect 114545 32946 114579 32958
rect 113784 31322 113794 32680
rect 113812 31322 113822 32652
rect 113855 31322 113921 32946
rect 114513 31322 114579 32946
rect 114606 31646 114612 32999
rect 114634 31618 114640 32999
rect 115197 32958 115271 32999
rect 115190 32957 115243 32958
rect 115160 32946 115243 32957
rect 115066 31322 115114 32714
rect 115171 32658 115243 32946
rect 115246 32658 115271 32958
rect 115861 32958 115907 33005
rect 115818 32946 115849 32957
rect 115861 32946 115895 32958
rect 115122 31322 115142 32658
rect 115171 31322 115237 32658
rect 115829 31334 115895 32946
rect 115829 31322 115863 31334
rect 113185 31318 115550 31322
rect 113185 31308 113231 31318
rect 113244 31308 115550 31318
rect 113185 31284 115550 31308
rect 113083 30832 113117 31235
rect 113185 31173 113231 31284
rect 113244 31275 115550 31284
rect 115817 31275 115876 31322
rect 115969 31275 116003 33005
rect 116083 31322 116117 33005
rect 116519 32957 116553 33104
rect 116476 32946 116553 32957
rect 116487 31334 116553 32946
rect 116487 31322 116532 31334
rect 116083 31275 116130 31322
rect 116475 31275 116534 31322
rect 113291 31241 113902 31275
rect 113937 31272 114560 31275
rect 113949 31241 114560 31272
rect 114607 31241 115218 31275
rect 115265 31241 115876 31275
rect 115907 31241 116534 31275
rect 113843 31225 113889 31241
rect 114501 31225 114547 31241
rect 115159 31225 115211 31241
rect 115817 31225 115863 31241
rect 115190 31173 115211 31225
rect 115829 31173 115863 31225
rect 115969 31173 116003 31241
rect 116083 31173 116117 31241
rect 116475 31225 116521 31241
rect 116487 31173 116521 31225
rect 116601 31173 116667 33107
rect 118118 33146 119557 33182
rect 121040 33408 124628 33442
rect 119616 33146 119650 33180
rect 120274 33146 120308 33180
rect 120932 33146 120966 33180
rect 121040 33146 121074 33408
rect 121101 33146 124628 33408
rect 118118 33131 124628 33146
rect 124725 33403 128277 33437
rect 124725 33245 124759 33403
rect 125469 33335 125516 33382
rect 126127 33335 126174 33382
rect 126785 33335 126832 33382
rect 127443 33335 127490 33382
rect 128101 33335 128148 33382
rect 124901 33301 125516 33335
rect 125559 33301 126174 33335
rect 126217 33301 126832 33335
rect 126875 33301 127490 33335
rect 127533 33301 128148 33335
rect 128046 33295 128113 33301
rect 128046 33267 128141 33288
rect 124885 33254 125485 33257
rect 125543 33254 126143 33257
rect 126201 33254 126801 33257
rect 126859 33254 127459 33257
rect 127517 33254 128117 33257
rect 128243 33245 128277 33403
rect 132016 33346 132032 33366
rect 124725 33211 128277 33245
rect 124725 33131 124759 33211
rect 124839 33131 124873 33211
rect 125497 33131 125531 33211
rect 126155 33131 126189 33211
rect 126813 33131 126847 33211
rect 127471 33131 127505 33211
rect 128129 33131 128163 33211
rect 128243 33131 128277 33211
rect 118118 33112 129407 33131
rect 118118 33082 119557 33112
rect 118118 33040 119594 33082
rect 119604 33060 119624 33106
rect 119604 33050 119662 33060
rect 119612 33044 119662 33050
rect 120214 33044 120252 33082
rect 120270 33060 120274 33078
rect 120270 33044 120320 33060
rect 120872 33044 120910 33082
rect 120928 33060 120932 33078
rect 120970 33060 120972 33112
rect 120928 33044 120978 33060
rect 121026 33050 121028 33076
rect 121040 33044 121074 33112
rect 121101 33097 129407 33112
rect 121101 33061 124628 33097
rect 121154 33044 121192 33061
rect 121530 33044 121568 33061
rect 118118 33010 119596 33040
rect 118118 33004 119568 33010
rect 116698 31596 116704 32948
rect 118118 32460 119557 33004
rect 119574 32976 119596 33010
rect 119616 33010 120252 33044
rect 120274 33010 120910 33044
rect 120932 33010 121568 33044
rect 119574 32971 119588 32976
rect 119616 32972 119662 33010
rect 120274 32972 120320 33010
rect 120932 33004 120978 33010
rect 121040 33004 121074 33010
rect 120932 32972 121004 33004
rect 119573 32960 119604 32971
rect 119616 32960 119650 32972
rect 120231 32960 120262 32971
rect 120274 32960 120308 32972
rect 120889 32960 120920 32971
rect 120932 32960 120966 32972
rect 118100 31602 119557 32460
rect 119574 31638 119650 32960
rect 113185 31139 116667 31173
rect 118118 31298 119557 31602
rect 119578 31348 119650 31638
rect 120242 31580 120308 32960
rect 120900 31580 120966 32960
rect 120970 31828 121004 32972
rect 121026 31828 121074 33004
rect 121040 31690 121074 31828
rect 120970 31602 121004 31690
rect 120970 31580 120972 31602
rect 120242 31348 120319 31580
rect 120900 31348 120977 31580
rect 121026 31546 121074 31690
rect 119578 31336 119618 31348
rect 120242 31336 120276 31348
rect 120900 31336 120972 31348
rect 121026 31336 121028 31546
rect 121040 31336 121074 31546
rect 121154 31580 121188 33010
rect 121590 32971 121624 33061
rect 121547 32960 121624 32971
rect 121154 31578 121199 31580
rect 121558 31578 121624 32960
rect 121672 31578 121738 33061
rect 121774 32692 121790 32694
rect 121768 31828 121790 32692
rect 121812 32596 121846 33061
rect 121812 32514 121912 32596
rect 121768 31588 121790 31690
rect 121812 31578 121846 32514
rect 122122 31902 122584 32540
rect 122176 31818 122526 31852
rect 121904 31690 121938 31702
rect 121904 31662 121938 31674
rect 122176 31578 122210 31818
rect 122492 31790 122526 31818
rect 122368 31750 122406 31788
rect 122458 31756 122526 31790
rect 122334 31716 122406 31750
rect 122386 31696 122446 31706
rect 122492 31696 122538 31756
rect 122386 31690 122464 31696
rect 122492 31690 122596 31696
rect 122386 31677 122418 31678
rect 122279 31666 122324 31677
rect 122367 31668 122418 31677
rect 122492 31668 122538 31690
rect 122367 31666 122464 31668
rect 122290 31578 122324 31666
rect 122378 31662 122464 31666
rect 122492 31662 122596 31668
rect 122378 31578 122412 31662
rect 122492 31612 122538 31662
rect 122470 31578 122538 31612
rect 123128 31578 123162 31612
rect 123786 31578 123820 31612
rect 124444 31578 124478 31612
rect 124558 31578 124592 33061
rect 124725 32434 124759 33097
rect 125426 32838 125440 32976
rect 125426 32578 125434 32838
rect 125454 32810 125468 32948
rect 125454 32578 125462 32810
rect 124839 32434 124852 32436
rect 124600 31664 124626 32402
rect 124725 32012 125362 32434
rect 125474 32426 125497 32454
rect 125474 32420 125550 32426
rect 125576 32420 125582 32480
rect 125604 32420 125610 32480
rect 125412 32386 125978 32420
rect 125412 32064 125446 32386
rect 125480 32270 125550 32386
rect 125576 32340 125582 32386
rect 125474 32244 125550 32270
rect 125474 32206 125565 32244
rect 125567 32238 125582 32340
rect 125604 32312 125610 32386
rect 125595 32306 125610 32312
rect 125783 32306 125794 32317
rect 125595 32272 125794 32306
rect 125595 32266 125610 32272
rect 125795 32244 125876 32291
rect 125567 32206 125582 32212
rect 125842 32206 125876 32244
rect 125474 32180 125550 32206
rect 125480 32098 125550 32180
rect 125474 32064 125550 32098
rect 125566 32064 125582 32206
rect 125595 32178 125610 32184
rect 125783 32178 125794 32189
rect 125594 32144 125794 32178
rect 125594 32064 125610 32144
rect 125944 32064 125978 32386
rect 125412 32030 125978 32064
rect 124725 31614 124759 32012
rect 124805 31664 124818 32012
rect 124839 31630 124852 32012
rect 125480 31970 125550 32030
rect 125426 31682 125452 31882
rect 125454 31654 125480 31910
rect 125566 31618 125582 32030
rect 125594 31646 125610 32030
rect 128243 31614 128277 33097
rect 124689 31578 128313 31614
rect 121154 31544 128313 31578
rect 121154 31516 121199 31544
rect 121126 31482 121199 31516
rect 121154 31336 121222 31482
rect 121558 31464 121624 31544
rect 121672 31464 121738 31544
rect 121812 31464 121846 31544
rect 122176 31464 122210 31544
rect 122290 31474 122324 31544
rect 122336 31474 122366 31476
rect 122378 31474 122412 31544
rect 122300 31468 122402 31474
rect 122296 31464 122406 31468
rect 122470 31464 122538 31544
rect 123128 31464 123162 31544
rect 123786 31464 123820 31544
rect 124444 31464 124478 31544
rect 124558 31464 124592 31544
rect 121224 31402 121296 31440
rect 121346 31430 124592 31464
rect 119572 31298 119622 31336
rect 120098 31298 120280 31336
rect 120298 31304 120940 31336
rect 120298 31298 120938 31304
rect 120956 31298 121222 31336
rect 121262 31298 121296 31402
rect 121558 31348 121624 31430
rect 121558 31332 121603 31348
rect 121558 31298 121596 31332
rect 118118 31264 119622 31298
rect 119678 31264 120280 31298
rect 120336 31264 120938 31298
rect 120982 31264 121596 31298
rect 118118 31196 119557 31264
rect 119572 31248 119618 31264
rect 120230 31248 120276 31264
rect 120888 31258 120934 31264
rect 120982 31258 120996 31264
rect 120888 31248 120940 31258
rect 120900 31202 120940 31248
rect 120900 31196 120934 31202
rect 121040 31196 121074 31264
rect 121154 31196 121222 31264
rect 121262 31200 121296 31264
rect 121558 31200 121592 31264
rect 121262 31196 121334 31200
rect 121558 31196 121603 31200
rect 121672 31196 121738 31430
rect 121799 31418 121800 31419
rect 121800 31417 121801 31418
rect 118118 31162 121738 31196
rect 121812 31344 121846 31430
rect 121858 31418 121859 31419
rect 121857 31417 121858 31418
rect 121812 31272 121857 31344
rect 122176 31338 122210 31430
rect 122318 31418 122406 31430
rect 122457 31418 122458 31419
rect 122334 31406 122406 31418
rect 122458 31417 122459 31418
rect 122470 31400 122538 31430
rect 123115 31418 123116 31419
rect 123116 31417 123117 31418
rect 122470 31338 122526 31400
rect 122176 31304 122526 31338
rect 121812 31186 121884 31272
rect 115190 30832 115211 31139
rect 111898 30798 115354 30832
rect 88094 30727 91718 30763
rect 83377 30693 91718 30727
rect 83377 27209 83411 30693
rect 83831 30692 83865 30693
rect 83831 30619 83871 30692
rect 83890 30619 83899 30664
rect 83831 30613 83865 30619
rect 84489 30613 84523 30693
rect 85147 30613 85181 30693
rect 85805 30613 85839 30693
rect 86463 30613 86497 30693
rect 86577 30613 86611 30693
rect 83432 30551 83513 30598
rect 83572 30579 86611 30613
rect 83831 30573 83865 30579
rect 83818 30567 83819 30568
rect 83819 30566 83820 30567
rect 83479 29983 83513 30551
rect 83831 30508 83871 30573
rect 83877 30567 83878 30568
rect 83876 30566 83877 30567
rect 83890 30536 83899 30573
rect 84476 30567 84477 30568
rect 84477 30566 84478 30567
rect 83819 29967 83820 29968
rect 83818 29966 83819 29967
rect 83831 29955 83865 30508
rect 83876 29967 83877 29968
rect 84477 29967 84478 29968
rect 83877 29966 83878 29967
rect 84476 29966 84477 29967
rect 84489 29955 84523 30579
rect 84535 30567 84536 30568
rect 85134 30567 85135 30568
rect 84534 30566 84535 30567
rect 85135 30566 85136 30567
rect 84534 29967 84535 29968
rect 85135 29967 85136 29968
rect 84535 29966 84536 29967
rect 85134 29966 85135 29967
rect 85147 29955 85181 30579
rect 85193 30567 85194 30568
rect 85792 30567 85793 30568
rect 85192 30566 85193 30567
rect 85793 30566 85794 30567
rect 85192 29967 85193 29968
rect 85793 29967 85794 29968
rect 85193 29966 85194 29967
rect 85792 29966 85793 29967
rect 85805 29955 85839 30579
rect 85851 30567 85852 30568
rect 86450 30567 86451 30568
rect 85850 30566 85851 30567
rect 86451 30566 86452 30567
rect 85850 29967 85851 29968
rect 86451 29967 86452 29968
rect 85851 29966 85852 29967
rect 86450 29966 86451 29967
rect 86463 29955 86497 30579
rect 86577 29955 86611 30579
rect 88094 29955 91736 30693
rect 104936 30668 104940 30673
rect 104866 30640 104912 30645
rect 104866 30633 104934 30640
rect 104872 30630 104934 30633
rect 83432 29893 83513 29940
rect 83572 29921 91736 29955
rect 83818 29909 83819 29910
rect 83819 29908 83820 29909
rect 83479 29325 83513 29893
rect 83819 29309 83820 29310
rect 83818 29308 83819 29309
rect 83831 29297 83865 29921
rect 83877 29909 83878 29910
rect 84476 29909 84477 29910
rect 83876 29908 83877 29909
rect 84477 29908 84478 29909
rect 84489 29312 84523 29921
rect 84535 29909 84536 29910
rect 85134 29909 85135 29910
rect 84534 29908 84535 29909
rect 85135 29908 85136 29909
rect 84714 29312 84926 29444
rect 83876 29309 83877 29310
rect 83877 29308 83878 29309
rect 84404 29297 84926 29312
rect 85135 29309 85136 29310
rect 85134 29308 85135 29309
rect 85147 29297 85181 29921
rect 85193 29909 85194 29910
rect 85792 29909 85793 29910
rect 85192 29908 85193 29909
rect 85793 29908 85794 29909
rect 85192 29309 85193 29310
rect 85793 29309 85794 29310
rect 85193 29308 85194 29309
rect 85792 29308 85793 29309
rect 85805 29297 85839 29921
rect 85851 29909 85852 29910
rect 86450 29909 86451 29910
rect 85850 29908 85851 29909
rect 86451 29908 86452 29909
rect 85850 29309 85851 29310
rect 86451 29309 86452 29310
rect 85851 29308 85852 29309
rect 86450 29308 86451 29309
rect 86463 29297 86497 29921
rect 86577 29297 86611 29921
rect 87288 29878 87678 29912
rect 86642 29396 86898 29402
rect 87288 29380 87322 29878
rect 87502 29810 87549 29857
rect 87464 29776 87549 29810
rect 87391 29717 87436 29728
rect 87519 29717 87564 29728
rect 87402 29541 87436 29717
rect 87530 29541 87564 29717
rect 87502 29482 87549 29529
rect 87464 29448 87549 29482
rect 87644 29380 87678 29878
rect 87798 29396 88054 29414
rect 86670 29368 86870 29374
rect 87288 29346 87678 29380
rect 87826 29368 88026 29386
rect 83432 29235 83513 29282
rect 83572 29263 86611 29297
rect 83818 29251 83819 29252
rect 83819 29250 83820 29251
rect 83479 28667 83513 29235
rect 83819 28651 83820 28652
rect 83818 28650 83819 28651
rect 83831 28639 83865 29263
rect 83877 29251 83878 29252
rect 83876 29250 83877 29251
rect 84404 29242 84926 29263
rect 85134 29251 85135 29252
rect 85135 29250 85136 29251
rect 83876 28651 83877 28652
rect 84477 28651 84478 28652
rect 83877 28650 83878 28651
rect 84476 28650 84477 28651
rect 84489 28639 84523 29242
rect 84714 28996 84926 29242
rect 84534 28651 84535 28652
rect 85135 28651 85136 28652
rect 84535 28650 84536 28651
rect 85134 28650 85135 28651
rect 85147 28639 85181 29263
rect 85193 29251 85194 29252
rect 85792 29251 85793 29252
rect 85192 29250 85193 29251
rect 85793 29250 85794 29251
rect 85192 28651 85193 28652
rect 85793 28651 85794 28652
rect 85193 28650 85194 28651
rect 85792 28650 85793 28651
rect 85805 28639 85839 29263
rect 85851 29251 85852 29252
rect 86450 29251 86451 29252
rect 85850 29250 85851 29251
rect 86451 29250 86452 29251
rect 85850 28651 85851 28652
rect 86451 28651 86452 28652
rect 85851 28650 85852 28651
rect 86450 28650 86451 28651
rect 86463 28639 86497 29263
rect 86577 28639 86611 29263
rect 86870 29182 87130 29202
rect 86870 29154 87130 29174
rect 87274 28676 87696 29296
rect 87826 29186 88026 29202
rect 87798 29158 88054 29174
rect 88094 28639 91736 29921
rect 102714 29219 103150 29242
rect 102748 29185 103116 29208
rect 103621 29120 103655 30587
rect 104880 30448 104934 30630
rect 104880 30160 104912 30448
rect 104872 30157 104912 30160
rect 104866 30145 104912 30157
rect 104936 30420 104962 30668
rect 106182 30642 106228 30645
rect 106164 30633 106228 30642
rect 112610 30644 112614 30649
rect 106164 30630 106222 30633
rect 106164 30456 106180 30630
rect 112610 30458 112638 30644
rect 104936 30117 104940 30420
rect 106182 30157 106222 30160
rect 106182 30145 106228 30157
rect 104934 30064 105502 30098
rect 107706 29798 107930 29818
rect 109898 29802 110118 29822
rect 107726 29646 107727 29798
rect 107910 29646 107930 29798
rect 109918 29646 109919 29802
rect 110098 29646 110118 29802
rect 112610 29606 112614 30458
rect 83432 28577 83513 28624
rect 83572 28605 91736 28639
rect 83818 28593 83819 28594
rect 83819 28592 83820 28593
rect 83479 28009 83513 28577
rect 83819 27993 83820 27994
rect 83818 27992 83819 27993
rect 83831 27981 83865 28605
rect 83877 28593 83878 28594
rect 84476 28593 84477 28594
rect 83876 28592 83877 28593
rect 84477 28592 84478 28593
rect 83876 27993 83877 27994
rect 84477 27993 84478 27994
rect 83877 27992 83878 27993
rect 84476 27992 84477 27993
rect 84489 27981 84523 28605
rect 84535 28593 84536 28594
rect 85134 28593 85135 28594
rect 84534 28592 84535 28593
rect 85135 28592 85136 28593
rect 84534 27993 84535 27994
rect 85135 27993 85136 27994
rect 84535 27992 84536 27993
rect 85134 27992 85135 27993
rect 85147 27981 85181 28605
rect 85193 28593 85194 28594
rect 85792 28593 85793 28594
rect 85192 28592 85193 28593
rect 85793 28592 85794 28593
rect 85192 27993 85193 27994
rect 85793 27993 85794 27994
rect 85193 27992 85194 27993
rect 85792 27992 85793 27993
rect 85805 27981 85839 28605
rect 85851 28593 85852 28594
rect 86450 28593 86451 28594
rect 85850 28592 85851 28593
rect 86451 28592 86452 28593
rect 85850 27993 85851 27994
rect 86451 27993 86452 27994
rect 85851 27992 85852 27993
rect 86450 27992 86451 27993
rect 86463 27981 86497 28605
rect 86577 27981 86611 28605
rect 87838 28534 87880 28540
rect 88018 28534 88046 28540
rect 87810 28506 87880 28512
rect 88018 28506 88074 28512
rect 83432 27919 83513 27966
rect 83572 27947 86611 27981
rect 83818 27935 83819 27936
rect 83819 27934 83820 27935
rect 83479 27351 83513 27919
rect 83819 27335 83820 27336
rect 83818 27334 83819 27335
rect 83831 27323 83865 27947
rect 83877 27935 83878 27936
rect 84476 27935 84477 27936
rect 83876 27934 83877 27935
rect 84477 27934 84478 27935
rect 83876 27335 83877 27336
rect 84477 27335 84478 27336
rect 83877 27334 83878 27335
rect 84476 27334 84477 27335
rect 84489 27323 84523 27947
rect 84535 27935 84536 27936
rect 85134 27935 85135 27936
rect 84534 27934 84535 27935
rect 85135 27934 85136 27935
rect 84534 27335 84535 27336
rect 85135 27335 85136 27336
rect 84535 27334 84536 27335
rect 85134 27334 85135 27335
rect 85147 27323 85181 27947
rect 85193 27935 85194 27936
rect 85792 27935 85793 27936
rect 85192 27934 85193 27935
rect 85793 27934 85794 27935
rect 85192 27335 85193 27336
rect 85793 27335 85794 27336
rect 85193 27334 85194 27335
rect 85792 27334 85793 27335
rect 85805 27323 85839 27947
rect 85851 27935 85852 27936
rect 86450 27935 86451 27936
rect 85850 27934 85851 27935
rect 86451 27934 86452 27935
rect 85850 27335 85851 27336
rect 86451 27335 86452 27336
rect 85851 27334 85852 27335
rect 86450 27334 86451 27335
rect 86463 27323 86497 27947
rect 86577 27323 86611 27947
rect 87276 27941 87532 27960
rect 87304 27913 87504 27932
rect 83572 27289 86611 27323
rect 83831 27209 83865 27289
rect 84489 27209 84523 27289
rect 85147 27209 85181 27289
rect 85805 27209 85839 27289
rect 86463 27209 86497 27289
rect 86577 27209 86611 27289
rect 88094 27209 91736 28605
rect 103078 29086 105218 29120
rect 103078 28595 103112 29086
rect 103519 29018 103553 29086
rect 103621 29018 103655 29086
rect 103254 28984 103655 29018
rect 103471 28937 103472 28938
rect 103472 28936 103473 28937
rect 103181 28925 103226 28936
rect 103192 28595 103226 28925
rect 103519 28623 103553 28984
rect 103237 28607 103238 28608
rect 103238 28606 103239 28607
rect 103460 28595 103471 28606
rect 103078 28561 103471 28595
rect 95846 27897 96102 27906
rect 95874 27869 96074 27878
rect 103078 27788 103112 28561
rect 103192 27949 103226 28561
rect 103238 28549 103239 28550
rect 103237 28548 103238 28549
rect 103472 28533 103553 28580
rect 103237 27949 103238 27950
rect 103238 27948 103239 27949
rect 103256 27948 103258 27971
rect 103519 27965 103553 28533
rect 103256 27937 103286 27943
rect 103460 27937 103471 27948
rect 103154 27924 103472 27937
rect 103154 27911 103476 27924
rect 103204 27903 103476 27911
rect 103214 27897 103472 27903
rect 103238 27891 103472 27897
rect 103242 27890 103294 27891
rect 103621 27890 103655 28984
rect 106396 28728 106420 28938
rect 104550 28212 104574 28220
rect 104550 27960 104576 28212
rect 104550 27948 104574 27960
rect 103238 27869 103655 27890
rect 103254 27856 103655 27869
rect 103519 27788 103553 27856
rect 103621 27788 103655 27856
rect 83377 27175 91718 27209
rect 86577 26860 86611 27175
rect 88094 27139 91718 27175
rect 83336 26824 86647 26860
rect 88130 26824 88164 27139
rect 90248 26874 90252 27036
rect 90286 26912 90290 26998
rect 88244 26824 88278 26858
rect 88902 26824 88936 26858
rect 89560 26824 89594 26858
rect 90218 26824 90252 26858
rect 90876 26824 90910 26858
rect 91534 26824 91568 26858
rect 83336 26790 91580 26824
rect 91648 26790 91658 26858
rect 83336 25820 86647 26790
rect 88130 26710 88164 26790
rect 88244 26710 88278 26790
rect 88902 26710 88936 26790
rect 89560 26710 89594 26790
rect 90218 26710 90252 26790
rect 90876 26710 90910 26790
rect 91534 26710 91568 26790
rect 91652 26728 91682 26762
rect 88130 26688 91568 26710
rect 91648 26695 91652 26698
rect 88130 26686 91574 26688
rect 88130 26676 91580 26686
rect 87416 26306 87864 26468
rect 87340 26256 87864 26306
rect 87340 26152 87494 26256
rect 83328 25200 86647 25820
rect 56720 24759 57340 25144
rect 57390 25096 57956 25130
rect 57390 24964 57424 25096
rect 57545 25026 57582 25050
rect 57762 25027 57801 25050
rect 57761 25026 57801 25027
rect 57761 25022 57772 25026
rect 57445 24964 57526 25001
rect 57573 24998 57582 25022
rect 57761 25016 57773 25022
rect 57585 25001 57773 25016
rect 57585 24998 57854 25001
rect 57585 24982 57772 24998
rect 57773 24964 57854 24998
rect 57922 24964 57956 25096
rect 83336 25035 86647 25200
rect 88130 26052 88164 26676
rect 88244 26052 88278 26676
rect 88290 26664 88291 26665
rect 88889 26664 88890 26665
rect 88289 26663 88290 26664
rect 88890 26663 88891 26664
rect 88289 26064 88290 26065
rect 88890 26064 88891 26065
rect 88290 26063 88291 26064
rect 88889 26063 88890 26064
rect 88902 26052 88936 26676
rect 88948 26664 88949 26665
rect 89547 26664 89548 26665
rect 88947 26663 88948 26664
rect 89548 26663 89549 26664
rect 88947 26064 88948 26065
rect 89548 26064 89549 26065
rect 88948 26063 88949 26064
rect 89547 26063 89548 26064
rect 89560 26052 89594 26676
rect 89606 26664 89607 26665
rect 90205 26664 90206 26665
rect 89605 26663 89606 26664
rect 90206 26663 90207 26664
rect 89605 26064 89606 26065
rect 90206 26064 90207 26065
rect 89606 26063 89607 26064
rect 90205 26063 90206 26064
rect 90218 26052 90252 26676
rect 90264 26664 90265 26665
rect 90863 26664 90864 26665
rect 90263 26663 90264 26664
rect 90864 26663 90865 26664
rect 90858 26065 90864 26086
rect 90263 26064 90264 26065
rect 90858 26064 90865 26065
rect 90264 26063 90265 26064
rect 90858 26052 90864 26064
rect 90876 26052 90910 26676
rect 90922 26664 90923 26665
rect 91521 26664 91522 26665
rect 90921 26663 90922 26664
rect 91522 26663 91523 26664
rect 91534 26660 91580 26676
rect 91584 26660 91602 26664
rect 91534 26648 91602 26660
rect 91534 26592 91606 26648
rect 91534 26144 91580 26592
rect 91584 26144 91606 26592
rect 91534 26080 91606 26144
rect 91534 26068 91602 26080
rect 90921 26064 90922 26065
rect 91522 26064 91523 26065
rect 90922 26063 90923 26064
rect 91521 26063 91522 26064
rect 91534 26052 91580 26068
rect 91584 26064 91602 26068
rect 91614 26064 91618 26664
rect 91648 26080 91665 26695
rect 88130 26049 91580 26052
rect 88130 26040 91574 26049
rect 88130 26030 91568 26040
rect 91648 26037 91652 26080
rect 88130 26028 91574 26030
rect 88130 26018 91580 26028
rect 88130 25394 88164 26018
rect 88244 25394 88278 26018
rect 88290 26006 88291 26007
rect 88889 26006 88890 26007
rect 88289 26005 88290 26006
rect 88890 26005 88891 26006
rect 88289 25406 88290 25407
rect 88890 25406 88891 25407
rect 88290 25405 88291 25406
rect 88889 25405 88890 25406
rect 88902 25394 88936 26018
rect 88948 26006 88949 26007
rect 89547 26006 89548 26007
rect 88947 26005 88948 26006
rect 89548 26005 89549 26006
rect 88947 25406 88948 25407
rect 89548 25406 89549 25407
rect 88948 25405 88949 25406
rect 89547 25405 89548 25406
rect 89560 25394 89594 26018
rect 89606 26006 89607 26007
rect 90205 26006 90206 26007
rect 89605 26005 89606 26006
rect 90206 26005 90207 26006
rect 89605 25406 89606 25407
rect 90206 25406 90207 25407
rect 89606 25405 89607 25406
rect 90205 25405 90206 25406
rect 90218 25394 90252 26018
rect 90264 26006 90265 26007
rect 90858 26006 90864 26018
rect 90263 26005 90264 26006
rect 90858 26005 90865 26006
rect 90858 26000 90864 26005
rect 90263 25406 90264 25407
rect 90864 25406 90865 25407
rect 90264 25405 90265 25406
rect 90863 25405 90864 25406
rect 90876 25394 90910 26018
rect 90922 26006 90923 26007
rect 91521 26006 91522 26007
rect 90921 26005 90922 26006
rect 91522 26005 91523 26006
rect 91534 26002 91580 26018
rect 91584 26002 91602 26006
rect 91534 25990 91602 26002
rect 91534 25940 91606 25990
rect 91534 25492 91580 25940
rect 91584 25492 91606 25940
rect 91534 25422 91606 25492
rect 91534 25410 91602 25422
rect 90921 25406 90922 25407
rect 91522 25406 91523 25407
rect 90922 25405 90923 25406
rect 91521 25405 91522 25406
rect 91534 25394 91580 25410
rect 91584 25406 91602 25410
rect 91614 25406 91618 26006
rect 91648 25422 91665 26037
rect 88130 25391 91580 25394
rect 88130 25382 91574 25391
rect 88130 25372 91568 25382
rect 91648 25379 91652 25422
rect 88130 25370 91574 25372
rect 88130 25360 91580 25370
rect 88130 25128 88164 25360
rect 88244 25280 88278 25360
rect 88290 25348 88291 25349
rect 88889 25348 88890 25349
rect 88289 25347 88290 25348
rect 88890 25347 88891 25348
rect 88902 25280 88936 25360
rect 88948 25348 88949 25349
rect 89547 25348 89548 25349
rect 88947 25347 88948 25348
rect 89548 25347 89549 25348
rect 89028 25296 89476 25304
rect 89560 25280 89594 25360
rect 89606 25348 89607 25349
rect 90205 25348 90206 25349
rect 89605 25347 89606 25348
rect 90206 25347 90207 25348
rect 90218 25280 90252 25360
rect 90264 25348 90265 25349
rect 90863 25348 90864 25349
rect 90263 25347 90264 25348
rect 90864 25347 90865 25348
rect 90876 25280 90910 25360
rect 90922 25348 90923 25349
rect 91521 25348 91522 25349
rect 90921 25347 90922 25348
rect 91522 25347 91523 25348
rect 91534 25344 91580 25360
rect 91584 25344 91602 25348
rect 91534 25332 91602 25344
rect 91534 25280 91606 25332
rect 91546 25276 91606 25280
rect 89000 25268 89504 25276
rect 91546 25268 91580 25276
rect 88874 25230 88912 25268
rect 89532 25230 89570 25268
rect 90190 25230 90228 25268
rect 90848 25230 90886 25268
rect 91506 25230 91544 25268
rect 91550 25264 91568 25268
rect 91584 25242 91606 25276
rect 91584 25230 91602 25242
rect 88306 25196 88912 25230
rect 88964 25196 89570 25230
rect 89622 25196 90228 25230
rect 90280 25196 90886 25230
rect 90938 25196 91544 25230
rect 91614 25132 91618 25348
rect 91648 25128 91665 25379
rect 88130 25094 91665 25128
rect 91686 25094 91720 26790
rect 92292 26436 92326 27762
rect 103078 27754 105218 27788
rect 103621 27570 103655 27754
rect 95468 27274 95484 27276
rect 95376 27165 95996 27274
rect 96108 27260 96550 27294
rect 96046 27233 96612 27260
rect 95376 27131 100800 27165
rect 95376 27095 95996 27131
rect 96046 26966 96080 27131
rect 96148 27097 96182 27100
rect 96476 27097 96510 27100
rect 96578 26966 96612 27131
rect 103066 27095 103691 27570
rect 92406 26436 92430 26470
rect 95888 26450 95922 26590
rect 96064 26550 100800 26584
rect 95968 26522 96070 26540
rect 95996 26494 96042 26512
rect 96002 26450 96036 26484
rect 101060 26450 101094 26484
rect 101174 26450 101208 26590
rect 103102 26450 103136 27095
rect 104446 27074 104466 27356
rect 103216 26450 103250 26484
rect 92198 26402 92492 26436
rect 95366 26416 103618 26450
rect 92292 26368 92326 26402
rect 92292 26300 92350 26368
rect 92424 26340 92440 26374
rect 92292 26040 92326 26300
rect 92344 26065 92360 26241
rect 92368 26065 92378 26241
rect 92394 26053 92444 26307
rect 92292 25972 92350 26040
rect 92406 26027 92416 26053
rect 92292 25904 92326 25972
rect 92406 25904 92430 25938
rect 92458 25904 92492 26402
rect 92198 25870 92492 25904
rect 92292 25820 92326 25870
rect 92256 25456 92506 25820
rect 92436 25270 92470 25282
rect 92214 25236 92470 25270
rect 95270 25228 95304 26354
rect 95888 26336 95922 26416
rect 96002 26336 96036 26416
rect 101060 26336 101094 26416
rect 101174 26336 101208 26416
rect 95888 26302 101208 26336
rect 95888 25572 95922 26302
rect 96002 25724 96036 26302
rect 96048 26290 96049 26291
rect 101047 26290 101048 26291
rect 96047 26289 96048 26290
rect 101048 26289 101049 26290
rect 96002 25708 96036 25712
rect 97072 25708 97112 25716
rect 97128 25708 97140 25744
rect 101060 25724 101094 26302
rect 101060 25708 101094 25712
rect 96030 25682 101066 25708
rect 96026 25678 101070 25682
rect 95968 25674 101128 25678
rect 96026 25644 101070 25674
rect 96048 25640 101070 25644
rect 96048 25632 101048 25640
rect 97072 25608 97112 25632
rect 97128 25618 97140 25632
rect 101174 25572 101208 26302
rect 103102 26220 103136 26416
rect 103204 26360 103262 26402
rect 103216 26356 103250 26360
rect 103244 26348 103432 26356
rect 103244 26342 103444 26348
rect 103182 26336 103444 26342
rect 103178 26334 103444 26336
rect 103182 26322 103444 26334
rect 103240 26312 103444 26322
rect 103240 26302 103554 26312
rect 103262 26290 103554 26302
rect 103278 26288 103554 26290
rect 103482 26220 103516 26274
rect 103584 26220 103618 26416
rect 103102 26186 103926 26220
rect 103482 25726 103516 26186
rect 103584 25726 103618 26186
rect 106368 25980 106370 27368
rect 106344 25774 106370 25980
rect 106368 25768 106370 25774
rect 106694 26500 112614 29242
rect 113083 26500 113117 30798
rect 115190 30794 115211 30798
rect 113197 30761 113244 30777
rect 113185 30696 113244 30761
rect 113855 30746 113902 30777
rect 114513 30746 114560 30777
rect 115171 30746 115218 30777
rect 113843 30730 113902 30746
rect 114501 30730 114560 30746
rect 115159 30730 115218 30746
rect 113294 30696 113902 30730
rect 113952 30696 114560 30730
rect 114610 30696 115218 30730
rect 113185 30687 113220 30696
rect 113843 30687 113878 30696
rect 114501 30687 114536 30696
rect 115159 30687 115194 30696
rect 113185 30649 113231 30687
rect 113136 26608 113162 26724
rect 113164 26649 113190 26696
rect 113197 26649 113231 30649
rect 113232 30648 113265 30653
rect 113843 30649 113889 30687
rect 113232 28284 113266 30648
rect 113232 26661 113277 28284
rect 113286 26652 113290 26864
rect 113314 26649 113318 26892
rect 113855 26649 113889 30649
rect 113890 30648 113923 30653
rect 114501 30649 114547 30687
rect 113890 28284 113924 30648
rect 114513 29606 114547 30649
rect 114479 28938 114490 29606
rect 114507 28938 114547 29606
rect 113890 26661 113935 28284
rect 114513 27750 114547 28938
rect 114479 26684 114490 27750
rect 114507 26684 114547 27750
rect 114513 26649 114547 26684
rect 114548 30648 114581 30653
rect 115159 30649 115205 30687
rect 114548 28284 114582 30648
rect 115109 28938 115140 29606
rect 115165 28938 115168 29606
rect 114548 26661 114593 28284
rect 114606 26654 114616 26862
rect 114634 26649 114644 26890
rect 115109 26649 115140 27750
rect 115165 26649 115168 27750
rect 115171 26649 115205 30649
rect 115206 30648 115239 30653
rect 115206 28284 115240 30648
rect 115206 26661 115251 28284
rect 113164 26608 113244 26649
rect 113185 26568 113244 26608
rect 113247 26602 113902 26649
rect 113905 26602 114560 26649
rect 114563 26602 115218 26649
rect 113185 26552 113220 26568
rect 113185 26537 113200 26552
rect 113254 26534 113272 26602
rect 113282 26568 113902 26602
rect 113952 26568 114560 26602
rect 113282 26562 113300 26568
rect 113843 26552 113878 26568
rect 114501 26552 114536 26568
rect 114570 26534 114580 26602
rect 114598 26562 114608 26602
rect 114610 26568 115218 26602
rect 115159 26552 115211 26568
rect 115190 26500 115211 26552
rect 115320 26500 115354 30798
rect 106694 26469 115354 26500
rect 115829 26469 115863 31139
rect 115969 26469 116003 31139
rect 116083 28284 116117 31139
rect 116302 28996 116304 29152
rect 116487 28284 116521 31139
rect 116083 26469 116128 28284
rect 116487 26469 116532 28284
rect 116601 26469 116635 31139
rect 117374 29616 117433 29650
rect 118019 29626 118034 29708
rect 117312 29582 117702 29616
rect 118057 29588 118072 29746
rect 116638 28938 116648 29134
rect 117312 29084 117346 29582
rect 117399 29421 117433 29582
rect 117526 29514 117573 29561
rect 117488 29480 117573 29514
rect 117445 29421 117460 29432
rect 117543 29421 117588 29432
rect 117399 29245 117460 29421
rect 117554 29245 117588 29421
rect 117399 29118 117433 29245
rect 117526 29186 117573 29233
rect 117488 29152 117573 29186
rect 117374 29084 117433 29118
rect 117668 29084 117702 29582
rect 116694 28938 116704 29078
rect 117312 29050 117702 29084
rect 117298 28380 117720 29000
rect 118023 28938 118050 29090
rect 118051 28938 118097 29146
rect 117300 27408 117306 27664
rect 117328 27436 117334 27636
rect 106694 26466 116635 26469
rect 106694 26126 112614 26466
rect 113083 26373 113117 26466
rect 113165 26435 116635 26466
rect 106694 25906 112624 26126
rect 103404 25712 103796 25726
rect 103340 25700 103796 25712
rect 103404 25684 103796 25700
rect 104470 25690 105016 25726
rect 105566 25696 105892 25726
rect 106228 25696 106558 25726
rect 103312 25678 103796 25684
rect 103312 25672 103444 25678
rect 103584 25670 103618 25678
rect 103404 25622 103852 25670
rect 104442 25662 105044 25670
rect 105538 25668 105892 25670
rect 106228 25668 106586 25670
rect 95888 25538 101208 25572
rect 92364 25194 102616 25228
rect 95270 25114 95304 25194
rect 102582 25138 102616 25194
rect 95341 25118 95444 25126
rect 95334 25114 95444 25118
rect 102430 25114 102441 25125
rect 102442 25118 102616 25138
rect 95236 25080 102441 25114
rect 57390 24943 58046 24964
rect 57356 24909 58046 24943
rect 68386 24920 70026 24940
rect 57390 24897 58046 24909
rect 57392 24890 58046 24897
rect 57569 24875 57777 24888
rect 57573 24863 57773 24875
rect 57390 24836 57424 24863
rect 57569 24854 57777 24863
rect 57573 24842 57773 24854
rect 57922 24836 57956 24863
rect 57535 24828 57811 24829
rect 57424 24795 57922 24828
rect 57424 24761 57922 24774
rect 45246 24271 45280 24305
rect 48304 24271 48338 24305
rect 51362 24271 51396 24305
rect 51476 24271 51510 24516
rect 43719 24237 51989 24271
rect 43719 23658 43753 24237
rect 45246 24157 45280 24237
rect 48304 24157 48338 24237
rect 51362 24157 51396 24237
rect 51476 24157 51510 24237
rect 43774 24095 43855 24142
rect 43914 24123 51510 24157
rect 45233 24111 45234 24112
rect 45234 24110 45235 24111
rect 43821 23658 43855 24095
rect 44902 24082 44958 24096
rect 45246 23658 45280 24123
rect 45292 24111 45293 24112
rect 48291 24111 48292 24112
rect 45291 24110 45292 24111
rect 48292 24110 48293 24111
rect 45476 24082 45532 24096
rect 48304 23658 48338 24123
rect 48350 24111 48351 24112
rect 51349 24111 51350 24112
rect 48349 24110 48350 24111
rect 51350 24110 51351 24111
rect 51362 23658 51396 24123
rect 51476 23658 51510 24123
rect 41160 23594 57474 23658
rect 43719 23578 43753 23594
rect 43821 23578 43855 23594
rect 45246 23578 45280 23594
rect 48304 23578 48338 23594
rect 51054 23592 51110 23594
rect 51362 23578 51396 23594
rect 51476 23578 51510 23594
rect 41160 23514 57554 23578
rect 43719 20753 43753 23514
rect 45234 23511 45235 23512
rect 45233 23510 45234 23511
rect 45246 23499 45280 23514
rect 45291 23511 45292 23512
rect 48292 23511 48293 23512
rect 45292 23510 45293 23511
rect 48291 23510 48292 23511
rect 48304 23499 48338 23514
rect 48349 23511 48350 23512
rect 51350 23511 51351 23512
rect 48350 23510 48351 23511
rect 51349 23510 51350 23511
rect 51362 23499 51396 23514
rect 51476 23499 51510 23514
rect 43774 23437 43855 23484
rect 43914 23465 51510 23499
rect 45233 23453 45234 23454
rect 45234 23452 45235 23453
rect 43821 22869 43855 23437
rect 45246 23246 45280 23465
rect 45292 23453 45293 23454
rect 48291 23453 48292 23454
rect 45291 23452 45292 23453
rect 48292 23452 48293 23453
rect 44902 22934 44958 22938
rect 44902 22878 44958 22882
rect 45132 22862 45340 23246
rect 45476 22934 45532 22938
rect 45476 22878 45532 22882
rect 44630 22858 45340 22862
rect 44630 22841 45284 22858
rect 45291 22853 45292 22854
rect 48292 22853 48293 22854
rect 45292 22852 45293 22853
rect 48291 22852 48292 22853
rect 48304 22841 48338 23465
rect 48350 23453 48351 23454
rect 51349 23453 51350 23454
rect 48349 23452 48350 23453
rect 51350 23452 51351 23453
rect 51054 23414 51110 23438
rect 51054 23358 51110 23382
rect 48349 22853 48350 22854
rect 51350 22853 51351 22854
rect 48350 22852 48351 22853
rect 51349 22852 51350 22853
rect 51362 22841 51396 23465
rect 51476 22841 51510 23465
rect 60482 23240 60930 23320
rect 60480 23108 60930 23240
rect 60480 23012 60600 23108
rect 43774 22779 43855 22826
rect 43914 22807 51510 22841
rect 44630 22788 45284 22807
rect 45292 22795 45293 22796
rect 48291 22795 48292 22796
rect 45291 22794 45292 22795
rect 48292 22794 48293 22795
rect 43821 22211 43855 22779
rect 44902 22774 44958 22776
rect 44902 22718 44958 22720
rect 45084 22208 45240 22217
rect 45234 22195 45235 22196
rect 45233 22194 45234 22195
rect 45056 22183 45240 22189
rect 45246 22183 45280 22788
rect 45476 22774 45532 22776
rect 45476 22718 45532 22720
rect 45286 22208 45380 22217
rect 45291 22195 45292 22196
rect 48292 22195 48293 22196
rect 45292 22194 45293 22195
rect 48291 22194 48292 22195
rect 45286 22183 45408 22189
rect 48304 22183 48338 22807
rect 48350 22795 48351 22796
rect 51349 22795 51350 22796
rect 48349 22794 48350 22795
rect 51350 22794 51351 22795
rect 51054 22272 51110 22288
rect 51256 22242 51356 22260
rect 51054 22216 51110 22232
rect 51228 22214 51356 22232
rect 48349 22195 48350 22196
rect 51350 22195 51351 22196
rect 48350 22194 48351 22195
rect 51349 22194 51350 22195
rect 51362 22183 51396 22807
rect 51476 22260 51510 22807
rect 51402 22242 51510 22260
rect 51476 22232 51510 22242
rect 51402 22214 51510 22232
rect 51476 22183 51510 22214
rect 43774 22121 43855 22168
rect 43914 22149 51510 22183
rect 45233 22137 45234 22138
rect 45234 22136 45235 22137
rect 43821 21553 43855 22121
rect 44902 21602 44958 21618
rect 44902 21546 44958 21562
rect 45234 21537 45235 21538
rect 45233 21536 45234 21537
rect 45246 21525 45280 22149
rect 45292 22137 45293 22138
rect 48291 22137 48292 22138
rect 45291 22136 45292 22137
rect 48292 22136 48293 22137
rect 45476 21602 45532 21618
rect 45476 21546 45532 21562
rect 45291 21537 45292 21538
rect 48292 21537 48293 21538
rect 45292 21536 45293 21537
rect 48291 21536 48292 21537
rect 48304 21525 48338 22149
rect 48350 22137 48351 22138
rect 51349 22137 51350 22138
rect 48349 22136 48350 22137
rect 51350 22136 51351 22137
rect 51054 22104 51110 22106
rect 51054 22048 51110 22050
rect 48349 21537 48350 21538
rect 51350 21537 51351 21538
rect 48350 21536 48351 21537
rect 51349 21536 51350 21537
rect 51362 21525 51396 22149
rect 51476 21525 51510 22149
rect 43774 21463 43855 21510
rect 43914 21491 51510 21525
rect 45233 21479 45234 21480
rect 45234 21478 45235 21479
rect 43821 20895 43855 21463
rect 45234 20879 45235 20880
rect 45233 20878 45234 20879
rect 45246 20867 45280 21491
rect 45292 21479 45293 21480
rect 48291 21479 48292 21480
rect 45291 21478 45292 21479
rect 48292 21478 48293 21479
rect 45291 20879 45292 20880
rect 48292 20879 48293 20880
rect 45292 20878 45293 20879
rect 48291 20878 48292 20879
rect 48304 20867 48338 21491
rect 48350 21479 48351 21480
rect 51349 21479 51350 21480
rect 48349 21478 48350 21479
rect 51350 21478 51351 21479
rect 51054 20950 51110 20966
rect 51054 20894 51110 20910
rect 48349 20879 48350 20880
rect 51350 20879 51351 20880
rect 48350 20878 48351 20879
rect 51349 20878 51350 20879
rect 51362 20867 51396 21491
rect 51476 20867 51510 21491
rect 64928 21006 64962 24224
rect 68406 23578 68407 24920
rect 70006 23578 70026 24920
rect 83490 24782 83514 24798
rect 83468 24752 83514 24782
rect 83440 24724 83542 24726
rect 95270 24656 95304 25080
rect 95356 25068 95444 25080
rect 95372 25048 95406 25068
rect 102442 25052 102514 25090
rect 102480 25032 102514 25052
rect 102442 25020 102530 25032
rect 95334 24958 95406 24996
rect 95456 24986 102530 25020
rect 102442 24974 102530 24986
rect 95372 24668 95406 24958
rect 102480 24684 102514 24974
rect 95356 24660 95444 24668
rect 95334 24656 95444 24660
rect 102430 24656 102441 24667
rect 95236 24622 102441 24656
rect 95270 24542 95304 24622
rect 95341 24610 95444 24622
rect 102582 24542 102616 25118
rect 92364 24508 102616 24542
rect 68406 23308 70006 23328
rect 68406 23231 68407 23308
rect 70006 23231 70026 23308
rect 68406 23230 70026 23231
rect 95270 22994 95304 24508
rect 103584 22994 103618 25622
rect 106694 25322 112614 25906
rect 106694 25306 112654 25322
rect 106694 25058 112614 25306
rect 112654 25242 112670 25306
rect 112902 25242 112906 25322
rect 106694 24955 112615 25058
rect 112653 24994 112654 24995
rect 112654 24993 112655 24994
rect 112668 24955 112695 24998
rect 106694 24954 112614 24955
rect 106694 24634 112838 24954
rect 113069 24871 113117 26373
rect 113197 26383 113231 26435
rect 113855 26414 113889 26435
rect 114513 26414 114547 26435
rect 115171 26414 115211 26435
rect 115829 26414 115863 26435
rect 113813 26383 113889 26414
rect 114471 26383 114547 26414
rect 115129 26383 115211 26414
rect 115787 26383 115863 26414
rect 113197 26286 113243 26383
rect 113813 26367 113901 26383
rect 114471 26367 114559 26383
rect 115129 26367 115217 26383
rect 115787 26367 115875 26383
rect 115969 26367 116003 26435
rect 116083 26432 116128 26435
rect 116487 26432 116532 26435
rect 116083 26414 116117 26432
rect 116487 26414 116521 26432
rect 116083 26367 116130 26414
rect 116445 26367 116521 26414
rect 113245 26333 113901 26367
rect 113903 26333 114559 26367
rect 114561 26333 115217 26367
rect 115219 26333 115875 26367
rect 115877 26333 116521 26367
rect 113821 26327 113825 26333
rect 113849 26299 113853 26333
rect 113855 26286 113901 26333
rect 114513 26286 114559 26333
rect 115137 26327 115141 26333
rect 115165 26299 115169 26333
rect 115171 26286 115217 26333
rect 115829 26286 115875 26333
rect 113197 26274 113231 26286
rect 113830 26274 113843 26285
rect 113855 26274 113889 26286
rect 114488 26274 114501 26285
rect 114513 26274 114547 26286
rect 115146 26274 115159 26285
rect 115171 26274 115211 26286
rect 115804 26274 115817 26285
rect 115829 26274 115863 26286
rect 113183 24970 113231 26274
rect 113841 24970 113889 26274
rect 114499 24970 114547 26274
rect 113183 24898 113217 24970
rect 113841 24958 113875 24970
rect 114499 24958 114533 24970
rect 113219 24898 113223 24945
rect 113247 24911 113251 24917
rect 113827 24911 113875 24958
rect 114485 24911 114533 24958
rect 106694 24633 112614 24634
rect 106694 24526 112615 24633
rect 112654 24594 112655 24595
rect 112653 24593 112654 24594
rect 112668 24586 112695 24633
rect 106694 23322 112614 24526
rect 99486 22020 100124 22263
rect 96584 21894 96772 21920
rect 96556 21866 96744 21892
rect 95006 21819 95021 21859
rect 103155 21379 103189 21877
rect 95247 21345 103517 21379
rect 95006 21161 95021 21207
rect 43914 20833 51510 20867
rect 45246 20753 45280 20833
rect 48304 20753 48338 20833
rect 51362 20753 51396 20833
rect 51476 20753 51510 20833
rect 64438 20972 66690 21006
rect 64438 20916 64472 20972
rect 64826 20928 64860 20972
rect 64438 20892 64776 20916
rect 64928 20892 64962 20972
rect 64438 20882 64962 20892
rect 64438 20802 64472 20882
rect 64624 20858 64962 20882
rect 64540 20830 64574 20836
rect 64928 20802 64962 20858
rect 60480 20768 64962 20802
rect 43719 20719 51989 20753
rect 51476 20160 51510 20719
rect 59224 20144 59480 20170
rect 59252 20116 59452 20142
rect 47324 19634 47944 20056
rect 48304 20042 48338 20076
rect 47994 20008 48560 20042
rect 47994 19686 48028 20008
rect 48049 19906 48130 19913
rect 48049 19866 48138 19906
rect 48096 19828 48138 19866
rect 48116 19786 48138 19828
rect 48144 19758 48166 19934
rect 48304 19928 48338 20008
rect 48365 19928 48376 19939
rect 48189 19894 48376 19928
rect 48291 19882 48292 19883
rect 48292 19881 48293 19882
rect 48292 19812 48293 19813
rect 48291 19811 48292 19812
rect 48304 19800 48338 19894
rect 48350 19882 48351 19883
rect 48349 19881 48350 19882
rect 48377 19866 48458 19913
rect 48424 19828 48458 19866
rect 48349 19812 48350 19813
rect 48350 19811 48351 19812
rect 48365 19800 48376 19811
rect 48189 19766 48376 19800
rect 48304 19686 48338 19766
rect 48526 19686 48560 20008
rect 60196 19912 60550 20334
rect 64438 20160 64472 20768
rect 95247 20640 95281 21345
rect 101292 21299 101748 21327
rect 95402 21294 96584 21299
rect 96784 21294 101748 21299
rect 103100 21294 103106 21299
rect 95430 21266 96584 21271
rect 96784 21266 101748 21271
rect 102108 21265 102564 21286
rect 103006 21271 103118 21277
rect 103006 21266 103134 21271
rect 103006 21265 103118 21266
rect 95442 21262 103118 21265
rect 95302 21213 95383 21250
rect 95442 21235 103103 21262
rect 95426 21231 103103 21235
rect 95430 21225 96584 21231
rect 96784 21225 101348 21231
rect 102108 21218 102564 21231
rect 103006 21219 103103 21231
rect 101722 21216 102564 21218
rect 95302 21207 95430 21213
rect 95302 21201 96584 21207
rect 96784 21201 101348 21207
rect 101722 21201 102178 21216
rect 102994 21201 103005 21212
rect 95302 21197 103010 21201
rect 95302 21176 103005 21197
rect 103006 21176 103087 21186
rect 95302 21167 103087 21176
rect 95308 21161 96584 21167
rect 96784 21161 101348 21167
rect 95333 21155 95430 21161
rect 95336 21133 95343 21148
rect 95349 20669 95383 21155
rect 101722 21148 102178 21167
rect 102700 21161 103087 21167
rect 103006 21148 103087 21161
rect 95389 21133 96584 21148
rect 96784 21133 101348 21148
rect 102700 21139 103087 21148
rect 102700 21133 103034 21139
rect 99164 20964 99612 21036
rect 98740 20824 99612 20964
rect 98740 20752 99188 20824
rect 95349 20640 95732 20669
rect 95247 20636 95732 20640
rect 97134 20636 103047 20641
rect 95006 20503 95021 20549
rect 47994 19652 48560 19686
rect 54554 19576 54610 19588
rect 55002 19576 55058 19588
rect 56246 19576 56302 19588
rect 54554 19520 54610 19532
rect 55002 19520 55058 19532
rect 56246 19520 56302 19532
rect 60480 19249 60514 19912
rect 64402 19249 64993 19285
rect 56591 19238 60439 19249
rect 43706 18382 51546 19236
rect 56591 19226 60428 19238
rect 56591 19215 60439 19226
rect 60480 19215 64993 19249
rect 56591 18930 56625 19215
rect 60331 19135 60443 19147
rect 56786 19132 60443 19135
rect 56646 19073 56727 19120
rect 56786 19101 60428 19132
rect 60331 19089 60428 19101
rect 54554 18916 54610 18930
rect 55002 18916 55058 18930
rect 56246 18916 56302 18930
rect 56591 18916 56680 18930
rect 54554 18860 54610 18874
rect 55002 18860 55058 18874
rect 56246 18860 56302 18874
rect 56591 18868 56625 18916
rect 56693 18881 56727 19073
rect 60378 18896 60412 19089
rect 56557 18834 56625 18868
rect 56646 18880 56727 18881
rect 56646 18868 56774 18880
rect 60319 18868 60330 18879
rect 56646 18834 60330 18868
rect 42250 18348 51546 18382
rect 43706 18210 51546 18348
rect 54554 18256 54610 18272
rect 55002 18256 55058 18272
rect 56246 18256 56302 18272
rect 56591 18216 56625 18834
rect 56677 18822 56774 18834
rect 56693 18505 56727 18822
rect 60331 18806 60412 18853
rect 60378 18490 60412 18806
rect 60331 18489 60412 18490
rect 60331 18477 60428 18489
rect 56646 18415 56727 18462
rect 56786 18443 60428 18477
rect 60331 18431 60428 18443
rect 56693 18223 56727 18415
rect 60378 18238 60412 18431
rect 56646 18222 56727 18223
rect 56646 18216 56774 18222
rect 54554 18200 54610 18216
rect 55002 18200 55058 18216
rect 56246 18200 56302 18216
rect 56591 18210 56774 18216
rect 60319 18210 60330 18221
rect 56557 18200 60330 18210
rect 56557 18176 56625 18200
rect 56646 18176 60330 18200
rect 56591 18096 56625 18176
rect 56662 18164 56774 18176
rect 60480 18096 60514 19215
rect 54244 18062 60514 18096
rect 56591 17668 56625 18062
rect 43706 15612 51582 17662
rect 54244 17634 60514 17668
rect 56591 17554 56625 17634
rect 56557 17520 56625 17554
rect 56646 17554 56774 17566
rect 60319 17554 60330 17565
rect 56646 17520 60330 17554
rect 56591 17518 56625 17520
rect 56677 17518 56774 17520
rect 54554 17514 54610 17518
rect 55002 17514 55058 17518
rect 56246 17514 56302 17518
rect 56591 17514 56774 17518
rect 54554 17458 54610 17462
rect 55002 17458 55058 17462
rect 56246 17458 56302 17462
rect 56591 16958 56625 17514
rect 56677 17508 56774 17514
rect 56693 17189 56727 17508
rect 60331 17492 60412 17539
rect 60378 17174 60412 17492
rect 60331 17173 60412 17174
rect 60331 17161 60428 17173
rect 56646 17099 56727 17146
rect 56786 17127 60428 17161
rect 60331 17115 60428 17127
rect 54554 16956 54610 16958
rect 55002 16956 55058 16958
rect 56246 16956 56302 16958
rect 56591 16956 56664 16958
rect 56591 16902 56625 16956
rect 56693 16909 56727 17099
rect 60378 16924 60412 17115
rect 56646 16908 56727 16909
rect 56646 16902 56774 16908
rect 54554 16900 54610 16902
rect 55002 16900 55058 16902
rect 56246 16900 56302 16902
rect 56591 16900 56774 16902
rect 56591 16896 56625 16900
rect 56557 16862 56625 16896
rect 56646 16896 56774 16900
rect 60319 16896 60330 16907
rect 56646 16862 60330 16896
rect 55002 16292 55058 16300
rect 56246 16292 56302 16300
rect 56591 16244 56625 16862
rect 56677 16850 56774 16862
rect 56693 16531 56727 16850
rect 60331 16834 60412 16881
rect 60378 16516 60412 16834
rect 60331 16515 60412 16516
rect 60331 16503 60428 16515
rect 56646 16441 56727 16488
rect 56786 16469 60428 16503
rect 60331 16457 60428 16469
rect 56693 16251 56727 16441
rect 60378 16266 60412 16457
rect 56646 16250 56727 16251
rect 56646 16244 56774 16250
rect 54554 16236 54610 16244
rect 55002 16236 55058 16244
rect 56246 16236 56302 16244
rect 56591 16238 56774 16244
rect 60319 16238 60330 16249
rect 56557 16236 60330 16238
rect 56557 16204 56625 16236
rect 56646 16204 60330 16236
rect 56591 16150 56625 16204
rect 56677 16192 56774 16204
rect 54554 16142 54610 16150
rect 55002 16142 55058 16150
rect 56246 16142 56302 16150
rect 56591 16142 56680 16150
rect 56591 15731 56625 16142
rect 56693 15873 56727 16192
rect 60331 16176 60412 16223
rect 60378 15858 60412 16176
rect 60331 15857 60412 15858
rect 60331 15845 60428 15857
rect 56786 15814 60428 15845
rect 56786 15811 60443 15814
rect 60331 15799 60443 15811
rect 60480 15731 60514 17634
rect 64402 15731 64993 19215
rect 66650 18876 66684 20160
rect 95006 19845 95021 19891
rect 95247 19320 95281 20636
rect 95343 20623 95389 20636
rect 95430 20608 95732 20613
rect 96138 20607 96792 20626
rect 103053 20620 103087 21139
rect 103006 20619 103087 20620
rect 103006 20613 103103 20619
rect 97134 20608 103103 20613
rect 101292 20607 102756 20608
rect 103006 20607 103103 20608
rect 95302 20555 95383 20592
rect 95442 20577 103103 20607
rect 95426 20573 103103 20577
rect 96138 20564 96792 20573
rect 97134 20567 103103 20573
rect 95302 20543 95430 20555
rect 95734 20552 96792 20564
rect 103006 20561 103103 20567
rect 95734 20543 96388 20552
rect 102994 20549 103005 20554
rect 97134 20543 103006 20549
rect 95302 20539 103010 20543
rect 95302 20528 103006 20539
rect 95302 20509 103087 20528
rect 95333 20497 95430 20509
rect 95349 19977 95383 20497
rect 95734 20490 96388 20509
rect 96732 20503 103087 20509
rect 103006 20496 103087 20503
rect 96732 20481 103087 20496
rect 96732 20475 103034 20481
rect 96732 20447 97190 20475
rect 99164 20318 99612 20390
rect 98748 20178 99612 20318
rect 98748 20160 99196 20178
rect 101298 19983 101778 20011
rect 95402 19974 101778 19983
rect 95430 19949 101778 19955
rect 102130 19949 102586 19964
rect 103053 19962 103087 20481
rect 103006 19961 103087 19962
rect 103006 19949 103103 19961
rect 103155 19949 103189 21345
rect 113069 20160 113103 24871
rect 113183 24809 113223 24898
rect 113243 24898 113251 24911
rect 113259 24898 113875 24911
rect 113243 24877 113875 24898
rect 113901 24877 113909 24911
rect 113917 24877 114533 24911
rect 113247 24871 113300 24877
rect 113242 24843 113300 24870
rect 113829 24861 113875 24877
rect 114487 24861 114533 24877
rect 113242 24809 113251 24843
rect 113841 24809 113875 24861
rect 114499 24809 114533 24861
rect 114535 24843 114539 24945
rect 115080 24917 115082 26014
rect 115157 25986 115211 26274
rect 115108 24917 115110 25986
rect 115157 24958 115236 25986
rect 115143 24917 115236 24958
rect 115246 24917 115264 26014
rect 115815 24970 115863 26274
rect 115969 25105 116003 26333
rect 116083 25266 116117 26333
rect 116487 26285 116521 26333
rect 116462 26274 116521 26285
rect 116473 25254 116521 26274
rect 116473 25207 116533 25254
rect 116145 25173 116533 25207
rect 116402 25105 116404 25160
rect 116430 25105 116460 25160
rect 116473 25142 116533 25173
rect 116473 25105 116521 25142
rect 116587 25105 116635 26435
rect 117302 26036 117306 27036
rect 117378 26010 117452 26636
rect 117364 25856 117518 26010
rect 117282 25780 117306 25836
rect 117302 25522 117306 25780
rect 118023 25226 118042 27750
rect 118051 25254 118097 27750
rect 118118 26510 119557 31162
rect 120900 30004 120934 31162
rect 120162 29310 120624 29948
rect 120834 29922 120934 30004
rect 120252 29260 120276 29310
rect 120286 29260 120310 29310
rect 120220 29226 120570 29260
rect 120220 28752 120276 29226
rect 120286 28752 120310 29226
rect 120340 29158 120450 29196
rect 120378 29124 120450 29158
rect 120323 29074 120379 29085
rect 120411 29074 120467 29085
rect 120334 28898 120379 29074
rect 120422 28898 120467 29074
rect 120340 28848 120450 28886
rect 120378 28814 120450 28848
rect 120220 28746 120254 28752
rect 120536 28746 120570 29226
rect 120220 28712 120570 28746
rect 120862 28594 120898 28680
rect 120252 28406 120276 28534
rect 120286 28406 120310 28534
rect 118104 26474 119557 26510
rect 119584 26474 119618 26508
rect 120242 26474 120276 26508
rect 120900 26474 120934 29922
rect 120970 29528 120972 29606
rect 121026 29472 121028 29606
rect 120970 26474 120972 26640
rect 121026 26474 121028 26696
rect 121040 26474 121074 31162
rect 121154 28122 121222 31162
rect 121262 30834 121334 31162
rect 121558 30817 121603 31162
rect 121672 30817 121706 31162
rect 121812 31126 121857 31186
rect 122470 31126 122515 31304
rect 121800 30818 121801 30819
rect 121799 30817 121800 30818
rect 121335 30806 121752 30817
rect 121812 30806 121846 31126
rect 121857 30818 121858 30819
rect 122458 30818 122459 30819
rect 121858 30817 121859 30818
rect 122457 30817 122458 30818
rect 122470 30806 122504 31126
rect 122515 30818 122516 30819
rect 123116 30818 123117 30819
rect 122516 30817 122517 30818
rect 123115 30817 123116 30818
rect 123128 30806 123162 31430
rect 123174 31418 123175 31419
rect 123773 31418 123774 31419
rect 123173 31417 123174 31418
rect 123774 31417 123775 31418
rect 123173 30818 123174 30819
rect 123774 30818 123775 30819
rect 123174 30817 123175 30818
rect 123773 30817 123774 30818
rect 123786 30806 123820 31430
rect 123832 31418 123833 31419
rect 124431 31418 124432 31419
rect 123831 31417 123832 31418
rect 124432 31417 124433 31418
rect 123831 30818 123832 30819
rect 124432 30818 124433 30819
rect 123832 30817 123833 30818
rect 124431 30817 124432 30818
rect 124444 30806 124478 31430
rect 124558 30806 124592 31430
rect 121224 30744 121334 30782
rect 121346 30772 124592 30806
rect 121262 30288 121334 30744
rect 121262 30176 121296 30288
rect 121558 30262 121603 30772
rect 121558 30148 121592 30262
rect 121672 30148 121706 30772
rect 121799 30760 121800 30761
rect 121800 30759 121801 30760
rect 121734 30232 121790 30246
rect 121734 30176 121790 30190
rect 121800 30160 121801 30161
rect 121799 30159 121800 30160
rect 121812 30148 121846 30772
rect 121858 30760 121859 30761
rect 122457 30760 122458 30761
rect 121857 30759 121858 30760
rect 122458 30759 122459 30760
rect 121857 30160 121858 30161
rect 122458 30160 122459 30161
rect 121858 30159 121859 30160
rect 122457 30159 122458 30160
rect 122470 30148 122504 30772
rect 122516 30760 122517 30761
rect 123115 30760 123116 30761
rect 122515 30759 122516 30760
rect 123116 30759 123117 30760
rect 122515 30160 122516 30161
rect 123116 30160 123117 30161
rect 122516 30159 122517 30160
rect 123115 30159 123116 30160
rect 123128 30148 123162 30772
rect 123174 30760 123175 30761
rect 123773 30760 123774 30761
rect 123173 30759 123174 30760
rect 123774 30759 123775 30760
rect 123173 30160 123174 30161
rect 123774 30160 123775 30161
rect 123174 30159 123175 30160
rect 123773 30159 123774 30160
rect 123786 30148 123820 30772
rect 123832 30760 123833 30761
rect 124431 30760 124432 30761
rect 123831 30759 123832 30760
rect 124432 30759 124433 30760
rect 123831 30160 123832 30161
rect 124432 30160 124433 30161
rect 123832 30159 123833 30160
rect 124431 30159 124432 30160
rect 124444 30148 124478 30772
rect 124558 30148 124592 30772
rect 121224 30086 121296 30124
rect 121346 30114 124592 30148
rect 121262 29518 121296 30086
rect 121558 29490 121592 30114
rect 121672 29490 121706 30114
rect 121799 30102 121800 30103
rect 121800 30101 121801 30102
rect 121800 29502 121801 29503
rect 121799 29501 121800 29502
rect 121812 29490 121846 30114
rect 121858 30102 121859 30103
rect 122457 30102 122458 30103
rect 121857 30101 121858 30102
rect 122458 30101 122459 30102
rect 121857 29502 121858 29503
rect 122458 29502 122459 29503
rect 121858 29501 121859 29502
rect 122457 29501 122458 29502
rect 122470 29490 122504 30114
rect 122516 30102 122517 30103
rect 123115 30102 123116 30103
rect 122515 30101 122516 30102
rect 123116 30101 123117 30102
rect 122515 29502 122516 29503
rect 123116 29502 123117 29503
rect 122516 29501 122517 29502
rect 123115 29501 123116 29502
rect 123128 29490 123162 30114
rect 123174 30102 123175 30103
rect 123773 30102 123774 30103
rect 123173 30101 123174 30102
rect 123774 30101 123775 30102
rect 123173 29502 123174 29503
rect 123774 29502 123775 29503
rect 123174 29501 123175 29502
rect 123773 29501 123774 29502
rect 123786 29490 123820 30114
rect 123832 30102 123833 30103
rect 124431 30102 124432 30103
rect 123831 30101 123832 30102
rect 124432 30101 124433 30102
rect 123831 29502 123832 29503
rect 124432 29502 124433 29503
rect 123832 29501 123833 29502
rect 124431 29501 124432 29502
rect 124444 29490 124478 30114
rect 124558 29490 124592 30114
rect 121224 29428 121296 29466
rect 121346 29456 124592 29490
rect 121262 28860 121296 29428
rect 121558 28832 121592 29456
rect 121672 28832 121706 29456
rect 121799 29444 121800 29445
rect 121800 29443 121801 29444
rect 121734 28910 121798 28924
rect 121734 28854 121790 28868
rect 121800 28844 121801 28845
rect 121799 28843 121800 28844
rect 121812 28832 121846 29456
rect 121858 29444 121859 29445
rect 122457 29444 122458 29445
rect 121857 29443 121858 29444
rect 122458 29443 122459 29444
rect 121857 28844 121858 28845
rect 122458 28844 122459 28845
rect 121858 28843 121859 28844
rect 122457 28843 122458 28844
rect 122470 28832 122504 29456
rect 122516 29444 122517 29445
rect 123115 29444 123116 29445
rect 122515 29443 122516 29444
rect 123116 29443 123117 29444
rect 122515 28844 122516 28845
rect 123116 28844 123117 28845
rect 122516 28843 122517 28844
rect 123115 28843 123116 28844
rect 123128 28832 123162 29456
rect 123174 29444 123175 29445
rect 123773 29444 123774 29445
rect 123173 29443 123174 29444
rect 123774 29443 123775 29444
rect 123173 28844 123174 28845
rect 123774 28844 123775 28845
rect 123174 28843 123175 28844
rect 123773 28843 123774 28844
rect 123786 28832 123820 29456
rect 123832 29444 123833 29445
rect 124431 29444 124432 29445
rect 123831 29443 123832 29444
rect 124432 29443 124433 29444
rect 123831 28844 123832 28845
rect 124432 28844 124433 28845
rect 123832 28843 123833 28844
rect 124431 28843 124432 28844
rect 124444 28832 124478 29456
rect 124558 28832 124592 29456
rect 121224 28770 121296 28808
rect 121346 28798 124592 28832
rect 121262 28202 121296 28770
rect 121558 28174 121592 28798
rect 121672 28174 121706 28798
rect 121799 28786 121800 28787
rect 121800 28785 121801 28786
rect 121734 28760 121798 28762
rect 121734 28704 121790 28706
rect 121812 28284 121846 28798
rect 121858 28786 121859 28787
rect 122457 28786 122458 28787
rect 121857 28785 121858 28786
rect 122458 28785 122459 28786
rect 122470 28284 122504 28798
rect 122516 28786 122517 28787
rect 123115 28786 123116 28787
rect 122515 28785 122516 28786
rect 123116 28785 123117 28786
rect 123128 28284 123162 28798
rect 123174 28786 123175 28787
rect 123773 28786 123774 28787
rect 123173 28785 123174 28786
rect 123774 28785 123775 28786
rect 123786 28284 123820 28798
rect 123832 28786 123833 28787
rect 124431 28786 124432 28787
rect 123831 28785 123832 28786
rect 124432 28785 124433 28786
rect 124444 28284 124478 28798
rect 121812 28187 121857 28284
rect 122470 28187 122515 28284
rect 123128 28187 123173 28284
rect 123786 28187 123831 28284
rect 121800 28186 121801 28187
rect 121812 28186 121858 28187
rect 122458 28186 122459 28187
rect 122470 28186 122516 28187
rect 123116 28186 123117 28187
rect 123128 28186 123174 28187
rect 123774 28186 123775 28187
rect 123786 28186 123832 28187
rect 124432 28186 124433 28187
rect 124444 28186 124489 28284
rect 121799 28185 121800 28186
rect 121812 28174 121846 28186
rect 121858 28185 121859 28186
rect 122457 28185 122458 28186
rect 121858 28174 122458 28185
rect 122470 28174 122504 28186
rect 122516 28185 122517 28186
rect 123115 28185 123116 28186
rect 122516 28174 123116 28185
rect 123128 28174 123162 28186
rect 123174 28185 123175 28186
rect 123773 28185 123774 28186
rect 123174 28174 123774 28185
rect 123786 28174 123820 28186
rect 123832 28185 123833 28186
rect 124431 28185 124432 28186
rect 123832 28174 124432 28185
rect 124444 28174 124478 28186
rect 124558 28174 124592 28798
rect 124689 29514 128313 31544
rect 128922 30114 129338 30136
rect 128956 30080 129372 30102
rect 124689 29422 128364 29514
rect 124689 29414 128313 29422
rect 124689 29402 128336 29414
rect 124689 29396 128564 29402
rect 124689 29394 128740 29396
rect 124689 28174 128313 29394
rect 128336 29368 128536 29374
rect 128336 29366 128768 29368
rect 128918 29310 129380 29948
rect 128976 29226 129326 29260
rect 128976 28746 129010 29226
rect 129168 29158 129206 29196
rect 129134 29124 129206 29158
rect 129079 29074 129124 29085
rect 129167 29074 129212 29085
rect 129090 28898 129124 29074
rect 129178 28898 129212 29074
rect 129168 28866 129206 28886
rect 129134 28844 129206 28866
rect 129118 28832 129206 28844
rect 129118 28798 129184 28832
rect 129292 28746 129326 29226
rect 128976 28712 129326 28746
rect 121346 28140 128313 28174
rect 121154 28060 121199 28122
rect 121558 28060 121592 28140
rect 121672 28060 121706 28140
rect 121812 28060 121846 28140
rect 122470 28060 122504 28140
rect 123128 28060 123162 28140
rect 123786 28060 123820 28140
rect 124444 28060 124478 28140
rect 124558 28060 124592 28140
rect 124689 28060 128313 28140
rect 121154 28026 128313 28060
rect 121154 28012 121199 28026
rect 121154 27972 121188 28012
rect 121154 27916 121199 27972
rect 121154 27830 121270 27916
rect 121154 27691 121199 27830
rect 121558 27691 121592 28026
rect 121672 27691 121706 28026
rect 121776 27754 121790 27954
rect 122474 27814 122504 27976
rect 122512 27852 122542 27938
rect 121720 27698 121734 27754
rect 124444 27691 124478 28026
rect 124558 27691 124592 28026
rect 124689 27990 128313 28026
rect 121119 27655 124628 27691
rect 124725 27655 124759 27990
rect 124839 27655 124873 27990
rect 125497 27655 125531 27689
rect 126155 27655 126189 27689
rect 126779 27655 126782 27750
rect 126807 27655 126810 27750
rect 126813 27655 126847 27689
rect 127471 27655 127505 27689
rect 128129 27655 128163 27689
rect 128243 27655 128277 27990
rect 121119 27621 129425 27655
rect 121119 26474 124628 27621
rect 118104 26469 124628 26474
rect 124725 27541 124759 27621
rect 124839 27541 124873 27621
rect 124885 27541 125485 27552
rect 125497 27541 125531 27621
rect 126155 27541 126189 27621
rect 126779 27547 126782 27621
rect 126807 27547 126810 27621
rect 126813 27541 126847 27621
rect 127471 27541 127505 27621
rect 128129 27541 128163 27621
rect 128243 27541 128277 27621
rect 124725 27507 128277 27541
rect 124725 26883 124759 27507
rect 124839 27495 124873 27507
rect 124885 27495 124886 27496
rect 125484 27495 125485 27496
rect 125497 27495 125531 27507
rect 125543 27495 125544 27496
rect 126142 27495 126143 27496
rect 124839 27494 124885 27495
rect 125485 27494 125486 27495
rect 125497 27494 125543 27495
rect 126143 27494 126144 27495
rect 124839 26896 124884 27494
rect 125497 26896 125542 27494
rect 124839 26895 124885 26896
rect 125485 26895 125486 26896
rect 125497 26895 125543 26896
rect 126143 26895 126144 26896
rect 124839 26883 124873 26895
rect 124885 26894 124886 26895
rect 125484 26894 125485 26895
rect 124885 26883 125485 26894
rect 125497 26883 125531 26895
rect 125543 26894 125544 26895
rect 126142 26894 126143 26895
rect 125543 26883 125580 26894
rect 126155 26883 126189 27507
rect 126201 27495 126202 27496
rect 126200 27494 126201 27495
rect 126779 27424 126782 27501
rect 126800 27495 126801 27496
rect 126801 27494 126802 27495
rect 126807 27424 126810 27501
rect 126200 26895 126201 26896
rect 126201 26894 126202 26895
rect 126779 26889 126782 26976
rect 126801 26895 126802 26896
rect 126800 26894 126801 26895
rect 126807 26889 126810 26976
rect 126813 26883 126847 27507
rect 126859 27495 126860 27496
rect 127458 27495 127459 27496
rect 126858 27494 126859 27495
rect 127459 27494 127460 27495
rect 127406 26976 127465 26986
rect 127434 26948 127465 26958
rect 126858 26895 126859 26896
rect 127459 26895 127460 26896
rect 126859 26894 126860 26895
rect 127458 26894 127459 26895
rect 127471 26883 127505 27507
rect 127517 27495 127518 27496
rect 128116 27495 128117 27496
rect 127516 27494 127517 27495
rect 128117 27494 128118 27495
rect 127511 26976 127570 26986
rect 127511 26948 127542 26958
rect 127516 26895 127517 26896
rect 128117 26895 128118 26896
rect 127517 26894 127518 26895
rect 128116 26894 128117 26895
rect 128129 26883 128163 27507
rect 128243 26883 128277 27507
rect 124725 26849 128277 26883
rect 124725 26469 124759 26849
rect 124839 26837 124873 26849
rect 124885 26837 124886 26838
rect 125484 26837 125485 26838
rect 125497 26837 125531 26849
rect 125543 26837 125544 26838
rect 126142 26837 126143 26838
rect 124839 26836 124885 26837
rect 125485 26836 125486 26837
rect 125497 26836 125543 26837
rect 126143 26836 126144 26837
rect 124839 26469 124884 26836
rect 118104 26440 125377 26469
rect 118104 26410 119557 26440
rect 118104 26338 119580 26410
rect 119584 26388 119618 26440
rect 117337 25198 117383 25213
rect 117370 25167 117383 25198
rect 118104 25105 119557 26338
rect 119584 26300 119630 26388
rect 120200 26372 120238 26410
rect 119632 26338 120238 26372
rect 120242 26388 120276 26440
rect 120242 26300 120288 26388
rect 120858 26372 120896 26410
rect 120290 26338 120896 26372
rect 120900 26388 120934 26440
rect 120900 26300 120946 26388
rect 120956 26378 120972 26440
rect 121026 26404 121028 26440
rect 121012 26378 121028 26404
rect 121040 26372 121074 26440
rect 121119 26436 125377 26440
rect 121119 26435 125402 26436
rect 121119 26372 124628 26435
rect 120948 26338 124628 26372
rect 124725 26367 124759 26435
rect 124839 26414 124884 26435
rect 124839 26367 124886 26414
rect 125012 26402 125402 26435
rect 125012 26367 125046 26402
rect 125201 26381 125248 26402
rect 125201 26367 125273 26381
rect 119559 26288 119572 26299
rect 119584 26288 119618 26300
rect 120217 26288 120230 26299
rect 120242 26288 120276 26300
rect 120875 26288 120888 26299
rect 120900 26288 120934 26300
rect 115969 25071 119557 25105
rect 115815 24958 115849 24970
rect 114563 24911 114567 24917
rect 115143 24911 115191 24917
rect 115801 24911 115849 24958
rect 116402 24917 116404 25071
rect 116430 24958 116460 25071
rect 116473 24970 116521 25071
rect 116473 24958 116507 24970
rect 116430 24917 116507 24958
rect 116459 24911 116507 24917
rect 114559 24877 114567 24911
rect 114575 24877 115191 24911
rect 115217 24877 115225 24911
rect 115233 24877 115849 24911
rect 115875 24877 115883 24911
rect 115891 24877 116507 24911
rect 114563 24871 114567 24877
rect 115145 24871 115191 24877
rect 115080 24864 115082 24871
rect 115108 24836 115110 24871
rect 115145 24861 115236 24871
rect 115157 24809 115236 24861
rect 115246 24809 115264 24871
rect 115803 24861 115849 24877
rect 116402 24864 116404 24871
rect 115815 24809 115849 24861
rect 116430 24809 116460 24871
rect 116461 24861 116507 24877
rect 116473 24809 116507 24861
rect 116587 24871 116635 25071
rect 118104 25035 119557 25071
rect 118140 24894 118188 25035
rect 118254 24984 118302 25035
rect 113171 24775 116519 24809
rect 113214 24642 113223 24775
rect 113242 24670 113251 24775
rect 115190 24634 115236 24775
rect 115190 24430 115197 24634
rect 115246 24606 115264 24775
rect 116430 24726 116446 24775
rect 95302 19897 95383 19934
rect 95430 19919 103103 19949
rect 95426 19915 103103 19919
rect 103121 19915 103223 19949
rect 95430 19909 101354 19915
rect 102110 19906 102586 19915
rect 95302 19891 95430 19897
rect 101706 19894 102586 19906
rect 103006 19903 103103 19915
rect 95302 19885 101354 19891
rect 101706 19885 102162 19894
rect 102994 19885 103005 19896
rect 95302 19881 103010 19885
rect 95302 19854 103005 19881
rect 103006 19854 103087 19870
rect 95302 19851 103087 19854
rect 95308 19845 101354 19851
rect 95333 19839 95430 19845
rect 95336 19817 95343 19826
rect 95349 19353 95383 19839
rect 101706 19836 102162 19851
rect 102706 19845 103087 19851
rect 103006 19835 103087 19845
rect 103006 19826 103093 19835
rect 103155 19826 103189 19915
rect 95389 19817 101354 19826
rect 102706 19810 103189 19826
rect 115190 19822 115197 23242
rect 116587 20160 116621 24871
rect 118140 20210 118174 24894
rect 118254 24832 118288 24984
rect 118358 24940 118374 25035
rect 118386 24940 118402 25035
rect 118840 24940 118848 25035
rect 118868 24940 118876 25035
rect 118912 24984 118960 25035
rect 119570 24984 119618 26288
rect 120228 24984 120276 26288
rect 120886 24984 120934 26288
rect 120956 25238 120972 26332
rect 121012 25196 121028 26332
rect 121040 25128 121074 26338
rect 121119 26314 124628 26338
rect 124633 26333 125273 26367
rect 121119 26231 124639 26314
rect 121119 26225 124628 26231
rect 124725 26225 124759 26333
rect 124839 26225 124873 26333
rect 125012 26225 125046 26333
rect 125188 26300 125273 26333
rect 125229 26285 125263 26290
rect 125218 26274 125263 26285
rect 125229 26257 125263 26274
rect 125229 26252 125274 26257
rect 125115 26241 125160 26252
rect 125126 26225 125160 26241
rect 125229 26225 125288 26252
rect 125343 26225 125402 26402
rect 125497 26432 125542 26836
rect 125485 26237 125486 26238
rect 125484 26236 125485 26237
rect 125497 26225 125531 26432
rect 125542 26237 125543 26238
rect 126143 26237 126144 26238
rect 125543 26236 125544 26237
rect 126142 26236 126143 26237
rect 126155 26225 126189 26849
rect 126201 26837 126202 26838
rect 126200 26836 126201 26837
rect 126779 26766 126782 26843
rect 126800 26837 126801 26838
rect 126801 26836 126802 26837
rect 126807 26766 126810 26843
rect 126200 26237 126201 26238
rect 126201 26236 126202 26237
rect 126779 26231 126782 26318
rect 126801 26237 126802 26238
rect 126800 26236 126801 26237
rect 126807 26231 126810 26318
rect 126813 26225 126847 26849
rect 126859 26837 126860 26838
rect 127458 26837 127459 26838
rect 126858 26836 126859 26837
rect 127459 26836 127460 26837
rect 127471 26510 127505 26849
rect 127517 26837 127518 26838
rect 128116 26837 128117 26838
rect 127516 26836 127517 26837
rect 128117 26836 128118 26837
rect 128046 26798 128123 26822
rect 128129 26510 128163 26849
rect 128243 26822 128277 26849
rect 128169 26798 128298 26822
rect 128243 26510 128277 26798
rect 126860 26474 129557 26510
rect 129796 26474 129830 33346
rect 132016 32730 132032 33300
rect 130638 31830 130660 32692
rect 130638 31588 130660 31692
rect 132016 31514 132036 32730
rect 132016 27738 132032 31514
rect 129910 26474 129944 26508
rect 126860 26440 130448 26474
rect 126858 26237 126859 26238
rect 126860 26237 129557 26440
rect 129664 26304 129684 26406
rect 129692 26332 129712 26378
rect 126859 26236 129557 26237
rect 126860 26225 129557 26236
rect 121119 26191 129557 26225
rect 121119 26185 124628 26191
rect 121119 26104 124639 26185
rect 121119 25662 124628 26104
rect 121119 25656 124698 25662
rect 121119 25567 124628 25656
rect 124644 25600 124698 25606
rect 124725 25567 124759 26191
rect 124839 25567 124873 26191
rect 125012 25904 125046 26191
rect 125126 26065 125160 26191
rect 125229 26065 125288 26191
rect 125229 26053 125274 26065
rect 125226 26049 125274 26053
rect 125226 26006 125273 26049
rect 125188 26000 125273 26006
rect 125343 26000 125402 26191
rect 125484 26179 125485 26180
rect 125485 26178 125486 26179
rect 125497 26000 125531 26191
rect 125543 26179 125544 26180
rect 126142 26179 126143 26180
rect 125542 26178 125543 26179
rect 126143 26178 126144 26179
rect 125080 25904 125531 26000
rect 125012 25870 125531 25904
rect 125080 25820 125531 25870
rect 124994 25788 125531 25820
rect 124994 25567 125416 25788
rect 125485 25579 125486 25580
rect 125484 25578 125485 25579
rect 125497 25567 125531 25788
rect 125542 25579 125543 25580
rect 125543 25578 125544 25579
rect 125614 25573 125616 25656
rect 126114 25578 126149 25601
rect 126086 25567 126149 25573
rect 126155 25567 126189 26191
rect 126201 26179 126202 26180
rect 126200 26178 126201 26179
rect 126779 26104 126782 26185
rect 126800 26179 126801 26180
rect 126801 26178 126802 26179
rect 126807 26104 126810 26185
rect 126195 25578 126222 25601
rect 126779 25573 126782 25656
rect 126801 25579 126802 25580
rect 126800 25578 126801 25579
rect 126807 25573 126810 25656
rect 126195 25567 126250 25573
rect 126813 25567 126847 26191
rect 126860 26180 129557 26191
rect 126859 26179 129557 26180
rect 126858 26178 126859 26179
rect 126858 25579 126859 25580
rect 126860 25579 129557 26179
rect 126859 25578 129557 25579
rect 126860 25567 129557 25578
rect 121119 25533 129557 25567
rect 121119 25128 124628 25533
rect 121040 25094 124628 25128
rect 121119 25058 124628 25094
rect 124725 25105 124759 25533
rect 124839 25276 124873 25533
rect 124994 25304 125416 25533
rect 125484 25521 125485 25522
rect 125485 25520 125486 25521
rect 125497 25304 125531 25533
rect 125543 25521 125544 25522
rect 125542 25520 125543 25521
rect 125614 25434 125616 25527
rect 126142 25521 126143 25522
rect 126143 25520 126144 25521
rect 124839 25266 124884 25276
rect 124994 25266 125531 25304
rect 126155 25266 126189 25533
rect 126201 25521 126202 25522
rect 126200 25520 126201 25521
rect 126779 25434 126782 25527
rect 126800 25521 126801 25522
rect 126801 25520 126802 25521
rect 126807 25434 126810 25527
rect 126813 25266 126847 25533
rect 126860 25522 129557 25533
rect 126859 25521 129557 25522
rect 126858 25520 126859 25521
rect 124994 25254 125520 25266
rect 124854 25207 125520 25254
rect 126127 25207 126174 25254
rect 126785 25207 126832 25254
rect 124901 25173 125520 25207
rect 125559 25173 126174 25207
rect 126217 25173 126832 25207
rect 125072 25105 125520 25173
rect 126860 25105 129557 25521
rect 124725 25071 129557 25105
rect 129796 25128 129830 26440
rect 129898 26338 130310 26410
rect 129898 26300 129956 26338
rect 129910 25280 129955 26300
rect 130289 26288 130345 26299
rect 130300 25268 130345 26288
rect 129934 25230 130346 25268
rect 129972 25196 130346 25230
rect 130288 25180 130346 25196
rect 130331 25165 130346 25180
rect 130414 25128 130448 26440
rect 131988 25236 131990 27682
rect 132016 25236 132046 27738
rect 130832 25196 131198 25218
rect 130870 25128 131242 25180
rect 131988 25144 131990 25190
rect 132016 25172 132046 25190
rect 129796 25094 133252 25128
rect 118912 24972 118946 24984
rect 119570 24972 119604 24984
rect 120228 24972 120262 24984
rect 120886 24972 120920 24984
rect 121119 24972 121742 25058
rect 118898 24934 118946 24972
rect 119556 24934 119610 24972
rect 118314 24900 118322 24934
rect 118330 24900 118946 24934
rect 118972 24900 118980 24934
rect 118988 24900 119610 24934
rect 118358 24832 118374 24894
rect 118386 24832 118402 24894
rect 118840 24888 118848 24894
rect 118868 24860 118876 24894
rect 118900 24884 118946 24900
rect 119558 24884 119610 24900
rect 118912 24832 118946 24884
rect 119566 24832 119610 24884
rect 119622 24832 119638 24972
rect 120214 24934 120262 24972
rect 120872 24934 120920 24972
rect 119646 24900 120262 24934
rect 120288 24900 120296 24934
rect 120304 24900 120920 24934
rect 120216 24884 120262 24900
rect 120874 24884 120920 24900
rect 120228 24832 120262 24884
rect 120886 24832 120920 24884
rect 120922 24866 120928 24968
rect 121038 24946 121742 24972
rect 120950 24934 120996 24940
rect 121038 24934 121758 24946
rect 120946 24930 121758 24934
rect 120946 24909 121742 24930
rect 121825 24909 121859 25058
rect 121939 24946 121984 25058
rect 122108 24946 122530 25058
rect 121939 24930 122056 24946
rect 122108 24930 122554 24946
rect 121939 24922 121984 24930
rect 121939 24921 121985 24922
rect 121939 24909 121973 24921
rect 121985 24920 121986 24921
rect 122108 24920 122530 24930
rect 122597 24922 122642 25058
rect 122682 24930 122714 24946
rect 123255 24922 123300 25058
rect 123913 24922 123958 25058
rect 124571 24922 124616 25058
rect 125214 24964 125284 25071
rect 122585 24921 122586 24922
rect 122597 24921 122643 24922
rect 123243 24921 123244 24922
rect 123255 24921 123301 24922
rect 123901 24921 123902 24922
rect 123913 24921 123959 24922
rect 124559 24921 124560 24922
rect 124571 24921 124617 24922
rect 125217 24921 125218 24922
rect 122584 24920 122585 24921
rect 121985 24909 122585 24920
rect 122597 24909 122631 24921
rect 122643 24920 122644 24921
rect 123242 24920 123243 24921
rect 122643 24909 123243 24920
rect 123255 24909 123289 24921
rect 123301 24920 123302 24921
rect 123900 24920 123901 24921
rect 123301 24909 123901 24920
rect 123913 24909 123947 24921
rect 123959 24920 123960 24921
rect 124558 24920 124559 24921
rect 123959 24909 124559 24920
rect 124571 24909 124605 24921
rect 124617 24920 124618 24921
rect 125216 24920 125217 24921
rect 125229 24909 125263 24964
rect 125343 24909 125377 25071
rect 120946 24900 125377 24909
rect 120950 24894 120984 24900
rect 121119 24875 125377 24900
rect 121119 24832 121742 24875
rect 118242 24798 121742 24832
rect 118358 24726 118374 24798
rect 118386 24726 118402 24798
rect 118358 22344 118374 23242
rect 118386 22344 118402 23242
rect 118358 21944 118374 22144
rect 118386 21944 118402 22144
rect 118358 20592 118374 21744
rect 118386 20564 118402 21744
rect 102706 19789 103087 19810
rect 99172 19622 99620 19694
rect 98740 19482 99620 19622
rect 98740 19410 99188 19482
rect 95349 19320 95754 19353
rect 95247 19304 95754 19320
rect 95006 19187 95021 19233
rect 66306 18172 66684 18876
rect 95006 18535 95021 18575
rect 95247 18455 95281 19304
rect 95430 19291 95754 19297
rect 96158 19291 96812 19310
rect 97156 19304 103047 19325
rect 103053 19304 103087 19789
rect 103093 19304 103106 19325
rect 103006 19303 103087 19304
rect 103006 19297 103103 19303
rect 97156 19291 103134 19297
rect 103155 19291 103189 19810
rect 95430 19276 103223 19291
rect 95302 19239 95383 19276
rect 95442 19261 103103 19276
rect 95426 19257 103103 19261
rect 103121 19257 103223 19276
rect 96158 19248 96812 19257
rect 97156 19251 103103 19257
rect 95302 19227 95430 19239
rect 95714 19236 96812 19248
rect 103006 19245 103103 19251
rect 95714 19227 96368 19236
rect 102994 19233 103005 19238
rect 97156 19227 103006 19233
rect 95302 19223 103010 19227
rect 95302 19220 103005 19223
rect 95302 19212 103006 19220
rect 95302 19193 103087 19212
rect 95333 19181 95430 19193
rect 95349 18661 95383 19181
rect 95714 19174 96368 19193
rect 101716 19192 103087 19193
rect 96710 19187 103087 19192
rect 103006 19165 103087 19187
rect 96710 19159 103034 19164
rect 96710 19131 97212 19159
rect 99164 18976 99612 19048
rect 98740 18836 99612 18976
rect 98740 18764 99188 18836
rect 95402 18652 95984 18667
rect 96184 18652 101772 18667
rect 103053 18646 103087 19165
rect 103006 18645 103087 18646
rect 95430 18633 95984 18639
rect 96184 18633 101772 18639
rect 103006 18633 103103 18645
rect 103155 18633 103189 19257
rect 113244 18634 113258 19822
rect 95302 18581 95383 18618
rect 95430 18603 103103 18633
rect 95426 18599 103103 18603
rect 103121 18599 103223 18633
rect 95430 18593 95992 18599
rect 95302 18575 95430 18581
rect 95984 18580 95992 18593
rect 96178 18593 101324 18599
rect 96178 18580 96184 18593
rect 102146 18582 102152 18596
rect 103006 18587 103103 18599
rect 95302 18569 95992 18575
rect 96178 18569 101324 18575
rect 102994 18569 103005 18580
rect 95302 18565 103010 18569
rect 95302 18535 103005 18565
rect 95318 18534 95430 18535
rect 95308 18529 95992 18534
rect 96178 18529 101324 18534
rect 102676 18529 103006 18534
rect 95318 18523 95430 18529
rect 103155 18506 103189 18599
rect 95336 18501 95343 18506
rect 95389 18501 95992 18506
rect 96178 18501 101324 18506
rect 102676 18500 103189 18506
rect 102676 18473 103062 18500
rect 103155 18455 103189 18500
rect 94919 18421 103189 18455
rect 66650 17862 66684 18172
rect 95247 17923 95281 18421
rect 115190 18301 115197 18634
rect 115157 18298 115197 18301
rect 116473 18298 116507 20160
rect 118012 19892 118028 20066
rect 118040 19918 118056 20038
rect 118104 19912 118220 20210
rect 118270 20118 118818 20152
rect 118270 20090 118304 20118
rect 118236 20056 118304 20090
rect 118038 19908 118220 19912
rect 118104 19748 118220 19908
rect 118270 19898 118322 20056
rect 118632 20038 118643 20049
rect 118334 19994 118406 20032
rect 118456 20004 118643 20038
rect 118644 19994 118716 20032
rect 118372 19960 118406 19994
rect 118632 19950 118643 19961
rect 118682 19960 118716 19994
rect 118456 19916 118643 19950
rect 118270 19836 118304 19898
rect 118784 19836 118818 20118
rect 118270 19802 118818 19836
rect 118238 19610 118312 19684
rect 118186 19538 118312 19610
rect 118912 19560 118946 24798
rect 119566 24726 119610 24798
rect 119622 24726 119638 24798
rect 121119 24762 121742 24798
rect 121119 24251 121728 24762
rect 121825 24289 121859 24875
rect 121901 24822 121902 24875
rect 121939 24863 121973 24875
rect 121985 24863 121986 24864
rect 122584 24863 122585 24864
rect 122597 24863 122631 24875
rect 122643 24863 122644 24864
rect 123242 24863 123243 24864
rect 123255 24863 123289 24875
rect 123301 24863 123302 24864
rect 123900 24863 123901 24864
rect 123913 24863 123947 24875
rect 123959 24863 123960 24864
rect 124558 24863 124559 24864
rect 124571 24863 124605 24875
rect 124617 24863 124618 24864
rect 125216 24863 125217 24864
rect 121939 24862 121985 24863
rect 122585 24862 122586 24863
rect 122597 24862 122643 24863
rect 123243 24862 123244 24863
rect 123255 24862 123301 24863
rect 123901 24862 123902 24863
rect 123913 24862 123959 24863
rect 124559 24862 124560 24863
rect 124571 24862 124617 24863
rect 125217 24862 125218 24863
rect 121939 24289 121984 24862
rect 121744 24284 122186 24289
rect 121825 24251 121859 24284
rect 121939 24264 121984 24284
rect 122597 24264 122642 24862
rect 123255 24264 123300 24862
rect 123913 24264 123958 24862
rect 124494 24288 124516 24313
rect 124571 24264 124616 24862
rect 121939 24263 121985 24264
rect 122585 24263 122586 24264
rect 122597 24263 122643 24264
rect 123243 24263 123244 24264
rect 123255 24263 123301 24264
rect 123901 24263 123902 24264
rect 123913 24263 123959 24264
rect 124559 24263 124560 24264
rect 124571 24263 124617 24264
rect 121939 24251 121973 24263
rect 121985 24262 121986 24263
rect 122584 24262 122585 24263
rect 121985 24251 122585 24262
rect 122597 24251 122631 24263
rect 122643 24262 122644 24263
rect 123242 24262 123243 24263
rect 122643 24251 123243 24262
rect 123255 24251 123289 24263
rect 123301 24262 123302 24263
rect 123900 24262 123901 24263
rect 123301 24251 123901 24262
rect 123913 24251 123947 24263
rect 123959 24262 123960 24263
rect 124558 24262 124559 24263
rect 123959 24251 124559 24262
rect 124571 24257 124611 24263
rect 124617 24262 124618 24263
rect 124571 24251 124605 24257
rect 124617 24251 124620 24262
rect 124628 24257 124639 24334
rect 125217 24263 125218 24264
rect 125216 24262 125217 24263
rect 125229 24251 125263 24875
rect 125343 24251 125377 24875
rect 121119 24246 125377 24251
rect 121119 24137 121728 24246
rect 121825 24217 125377 24246
rect 121825 24137 121859 24217
rect 121939 24137 121973 24217
rect 122597 24137 122631 24217
rect 123255 24137 123289 24217
rect 123913 24137 123947 24217
rect 124494 24211 124605 24217
rect 124565 24137 124611 24211
rect 124628 24137 124639 24211
rect 125229 24137 125263 24217
rect 125343 24137 125377 24217
rect 126860 24137 129557 25071
rect 121119 24103 129557 24137
rect 121119 24067 121728 24103
rect 119472 19822 119486 20060
rect 119566 20004 119610 23242
rect 119622 20004 119638 23242
rect 121544 22584 121578 22618
rect 121658 22584 121692 24067
rect 121720 24032 121768 24040
rect 121720 23998 121734 24006
rect 121825 22620 121859 24103
rect 124565 23482 124611 24103
rect 124628 23538 124639 24103
rect 124584 22904 124605 23442
rect 125343 23440 125377 24103
rect 126860 24067 129557 24103
rect 124584 22834 124611 22904
rect 124584 22696 124605 22834
rect 124584 22640 124611 22696
rect 124618 22668 124639 23408
rect 124760 23018 125380 23440
rect 125430 23036 125431 23426
rect 125764 23000 126032 23234
rect 125242 22660 125269 22916
rect 125270 22688 125297 22888
rect 126180 22774 126186 22876
rect 126214 22808 126220 22842
rect 124584 22636 124605 22640
rect 121789 22584 125413 22620
rect 121178 22550 125413 22584
rect 120850 19822 120866 19968
rect 120956 19822 120958 19844
rect 117350 19234 117504 19338
rect 117242 18934 117738 19234
rect 118238 19030 118312 19538
rect 118850 19474 118946 19560
rect 116556 18730 118198 18750
rect 116556 18674 118198 18694
rect 118912 18312 118946 19474
rect 120254 19396 120262 19446
rect 120244 18970 120262 19396
rect 120288 19362 120296 19412
rect 120278 19004 120296 19362
rect 121178 19066 121212 22550
rect 121544 22470 121578 22550
rect 121658 22470 121692 22550
rect 121242 22408 121314 22446
rect 121364 22436 121692 22470
rect 121531 22424 121532 22425
rect 121532 22423 121533 22424
rect 121280 21840 121314 22408
rect 121532 21824 121533 21825
rect 121531 21823 121532 21824
rect 121544 21812 121578 22436
rect 121658 21812 121692 22436
rect 121242 21750 121314 21788
rect 121364 21778 121692 21812
rect 121531 21766 121532 21767
rect 121532 21765 121533 21766
rect 121280 21182 121314 21750
rect 121532 21166 121533 21167
rect 121531 21165 121532 21166
rect 121544 21154 121578 21778
rect 121658 21154 121692 21778
rect 121242 21092 121314 21130
rect 121364 21120 121692 21154
rect 121531 21108 121532 21109
rect 121532 21107 121533 21108
rect 121280 20524 121314 21092
rect 121532 20508 121533 20509
rect 121531 20507 121532 20508
rect 121544 20496 121578 21120
rect 121658 20496 121692 21120
rect 121242 20434 121314 20472
rect 121364 20462 121692 20496
rect 121531 20450 121532 20451
rect 121532 20449 121533 20450
rect 121280 19866 121314 20434
rect 121544 19930 121578 20462
rect 121658 19930 121692 20462
rect 121789 22434 125413 22550
rect 126018 22584 126480 22620
rect 126896 22584 126930 24067
rect 127010 22584 127044 22618
rect 127668 22584 127702 22618
rect 128326 22584 128360 22618
rect 128984 22584 129018 22618
rect 126018 22550 129526 22584
rect 121789 22430 125664 22434
rect 121789 19930 125413 22430
rect 125436 22402 125636 22406
rect 126018 22342 126480 22550
rect 126896 22470 126930 22550
rect 127010 22470 127044 22550
rect 127668 22470 127702 22550
rect 128326 22470 128360 22550
rect 128984 22470 129018 22550
rect 129340 22470 129351 22481
rect 126564 22430 126820 22446
rect 126896 22436 129351 22470
rect 126592 22402 126792 22418
rect 126076 22258 126426 22292
rect 126076 21778 126110 22258
rect 126268 22190 126306 22228
rect 126234 22156 126306 22190
rect 126179 22106 126224 22117
rect 126267 22106 126312 22117
rect 126190 21930 126224 22106
rect 126278 21930 126312 22106
rect 126268 21916 126306 21918
rect 126190 21890 126312 21916
rect 126268 21888 126306 21890
rect 126218 21862 126306 21888
rect 126234 21846 126306 21862
rect 126218 21830 126284 21846
rect 126190 21802 126312 21818
rect 126330 21778 126364 21812
rect 126392 21778 126426 22258
rect 126076 21744 126426 21778
rect 126896 21812 126930 22436
rect 127010 21812 127044 22436
rect 127056 22424 127057 22425
rect 127655 22424 127656 22425
rect 127055 22423 127056 22424
rect 127656 22423 127657 22424
rect 127055 21824 127056 21825
rect 127656 21824 127657 21825
rect 127056 21823 127057 21824
rect 127655 21823 127656 21824
rect 127668 21812 127702 22436
rect 127714 22424 127715 22425
rect 128313 22424 128314 22425
rect 127713 22423 127714 22424
rect 128314 22423 128315 22424
rect 127713 21824 127714 21825
rect 128314 21824 128315 21825
rect 127714 21823 127715 21824
rect 128313 21823 128314 21824
rect 128326 21812 128360 22436
rect 128372 22424 128373 22425
rect 128971 22424 128972 22425
rect 128371 22423 128372 22424
rect 128972 22423 128973 22424
rect 128371 21824 128372 21825
rect 128972 21824 128973 21825
rect 128372 21823 128373 21824
rect 128971 21823 128972 21824
rect 128984 21812 129018 22436
rect 129030 22424 129031 22425
rect 129029 22423 129030 22424
rect 129352 22408 129424 22446
rect 129390 21840 129424 22408
rect 129029 21824 129030 21825
rect 129030 21823 129031 21824
rect 129340 21812 129351 21823
rect 126896 21778 129351 21812
rect 121544 19916 125413 19930
rect 121532 19850 121533 19851
rect 121531 19849 121532 19850
rect 121544 19844 121584 19916
rect 121544 19838 121578 19844
rect 121658 19838 121692 19916
rect 121242 19776 121314 19814
rect 121364 19804 121692 19838
rect 121531 19792 121532 19793
rect 121532 19791 121533 19792
rect 121280 19208 121314 19776
rect 121532 19192 121533 19193
rect 121531 19191 121532 19192
rect 121544 19180 121578 19804
rect 121658 19180 121692 19804
rect 121364 19146 121692 19180
rect 121544 19066 121578 19146
rect 121658 19066 121692 19146
rect 121789 19066 125413 19916
rect 126896 21154 126930 21778
rect 127010 21154 127044 21778
rect 127056 21766 127057 21767
rect 127655 21766 127656 21767
rect 127055 21765 127056 21766
rect 127656 21765 127657 21766
rect 127055 21166 127056 21167
rect 127656 21166 127657 21167
rect 127056 21165 127057 21166
rect 127655 21165 127656 21166
rect 127668 21154 127702 21778
rect 127714 21766 127715 21767
rect 128313 21766 128314 21767
rect 127713 21765 127714 21766
rect 128314 21765 128315 21766
rect 127713 21166 127714 21167
rect 128314 21166 128315 21167
rect 127714 21165 127715 21166
rect 128313 21165 128314 21166
rect 128326 21154 128360 21778
rect 128372 21766 128373 21767
rect 128971 21766 128972 21767
rect 128371 21765 128372 21766
rect 128972 21765 128973 21766
rect 128371 21166 128372 21167
rect 128972 21166 128973 21167
rect 128372 21165 128373 21166
rect 128971 21165 128972 21166
rect 128984 21154 129018 21778
rect 129030 21766 129031 21767
rect 129029 21765 129030 21766
rect 129352 21750 129424 21788
rect 129390 21182 129424 21750
rect 129029 21166 129030 21167
rect 129030 21165 129031 21166
rect 129340 21154 129351 21165
rect 126896 21120 129351 21154
rect 126896 20496 126930 21120
rect 127010 20496 127044 21120
rect 127056 21108 127057 21109
rect 127655 21108 127656 21109
rect 127055 21107 127056 21108
rect 127656 21107 127657 21108
rect 127055 20508 127056 20509
rect 127656 20508 127657 20509
rect 127056 20507 127057 20508
rect 127655 20507 127656 20508
rect 127668 20496 127702 21120
rect 127714 21108 127715 21109
rect 128313 21108 128314 21109
rect 127713 21107 127714 21108
rect 128314 21107 128315 21108
rect 127713 20508 127714 20509
rect 128314 20508 128315 20509
rect 127714 20507 127715 20508
rect 128313 20507 128314 20508
rect 128326 20496 128360 21120
rect 128372 21108 128373 21109
rect 128971 21108 128972 21109
rect 128371 21107 128372 21108
rect 128972 21107 128973 21108
rect 128371 20508 128372 20509
rect 128972 20508 128973 20509
rect 128372 20507 128373 20508
rect 128971 20507 128972 20508
rect 128984 20496 129018 21120
rect 129030 21108 129031 21109
rect 129029 21107 129030 21108
rect 129352 21092 129424 21130
rect 129390 20524 129424 21092
rect 129029 20508 129030 20509
rect 129030 20507 129031 20508
rect 129340 20496 129351 20507
rect 126896 20462 129351 20496
rect 126896 19838 126930 20462
rect 127010 19838 127044 20462
rect 127056 20450 127057 20451
rect 127655 20450 127656 20451
rect 127055 20449 127056 20450
rect 127656 20449 127657 20450
rect 127055 19850 127056 19851
rect 127656 19850 127657 19851
rect 127056 19849 127057 19850
rect 127655 19849 127656 19850
rect 127668 19838 127702 20462
rect 127714 20450 127715 20451
rect 128313 20450 128314 20451
rect 127713 20449 127714 20450
rect 128314 20449 128315 20450
rect 127713 19850 127714 19851
rect 128314 19850 128315 19851
rect 127714 19849 127715 19850
rect 128313 19849 128314 19850
rect 128326 19838 128360 20462
rect 128372 20450 128373 20451
rect 128971 20450 128972 20451
rect 128371 20449 128372 20450
rect 128972 20449 128973 20450
rect 128371 19850 128372 19851
rect 128972 19850 128973 19851
rect 128372 19849 128373 19850
rect 128971 19849 128972 19850
rect 128984 19838 129018 20462
rect 129030 20450 129031 20451
rect 129029 20449 129030 20450
rect 129352 20434 129424 20472
rect 129390 19866 129424 20434
rect 129029 19850 129030 19851
rect 129030 19849 129031 19850
rect 129340 19838 129351 19849
rect 126896 19804 129351 19838
rect 126896 19180 126930 19804
rect 127010 19180 127044 19804
rect 127056 19792 127057 19793
rect 127655 19792 127656 19793
rect 127055 19791 127056 19792
rect 127656 19791 127657 19792
rect 127055 19192 127056 19193
rect 127656 19192 127657 19193
rect 127056 19191 127057 19192
rect 127655 19191 127656 19192
rect 127668 19180 127702 19804
rect 127714 19792 127715 19793
rect 128313 19792 128314 19793
rect 127713 19791 127714 19792
rect 128314 19791 128315 19792
rect 128326 19656 128360 19804
rect 128372 19792 128373 19793
rect 128971 19792 128972 19793
rect 128371 19791 128372 19792
rect 128972 19791 128973 19792
rect 128308 19204 128382 19656
rect 127713 19192 127714 19193
rect 127714 19191 127715 19192
rect 127912 19180 128382 19204
rect 128972 19192 128973 19193
rect 128971 19191 128972 19192
rect 128984 19180 129018 19804
rect 129030 19792 129031 19793
rect 129029 19791 129030 19792
rect 129352 19776 129424 19814
rect 129390 19208 129424 19776
rect 129029 19192 129030 19193
rect 129030 19191 129031 19192
rect 129340 19180 129351 19191
rect 126896 19146 129351 19180
rect 126896 19066 126930 19146
rect 127010 19066 127044 19146
rect 127668 19066 127702 19146
rect 127912 19112 128382 19146
rect 128308 19066 128382 19112
rect 128984 19066 129018 19146
rect 129492 19066 129526 22550
rect 130414 20160 130448 25094
rect 130870 24604 131242 25094
rect 133350 24850 133362 25132
rect 133384 24884 133396 25106
rect 130500 24476 131242 24604
rect 130500 24284 130942 24476
rect 142468 23482 142668 23504
rect 129606 19822 129620 19844
rect 131058 19468 131092 20160
rect 131172 19468 131196 19502
rect 130964 19434 131258 19468
rect 131058 19400 131092 19434
rect 131058 19332 131116 19400
rect 131190 19339 131206 19434
rect 131058 19076 131092 19332
rect 131110 19081 131126 19289
rect 131138 19273 131144 19289
rect 131134 19097 131144 19273
rect 131138 19081 131144 19097
rect 131160 19085 131210 19339
rect 131032 19072 131096 19076
rect 131032 19066 131116 19072
rect 121178 19032 129526 19066
rect 119590 18602 119636 18634
rect 119590 18300 119610 18602
rect 119646 18574 119664 18634
rect 120850 18566 120864 18634
rect 121544 18594 121578 18628
rect 121658 18594 121692 19032
rect 121789 18996 125413 19032
rect 122112 18936 122146 18996
rect 122468 18936 122502 18996
rect 122597 18944 122631 18996
rect 122112 18902 122502 18936
rect 121866 18858 121938 18900
rect 122530 18858 122631 18944
rect 121866 18824 121952 18858
rect 121876 18786 121952 18824
rect 122094 18660 122516 18852
rect 122094 18634 122562 18660
rect 122094 18632 122516 18634
rect 121320 18560 121772 18594
rect 115151 18286 115197 18298
rect 121320 18278 121354 18560
rect 121544 18480 121578 18560
rect 121658 18486 121692 18560
rect 121658 18480 121694 18486
rect 121384 18436 121456 18474
rect 121506 18466 121694 18480
rect 121506 18446 121692 18466
rect 121422 18402 121456 18436
rect 121531 18434 121532 18435
rect 121532 18433 121533 18434
rect 121532 18404 121533 18405
rect 121531 18403 121532 18404
rect 121544 18392 121578 18446
rect 121658 18392 121692 18446
rect 121506 18358 121692 18392
rect 121544 18332 121578 18358
rect 121532 18300 121590 18332
rect 121544 18296 121578 18300
rect 121416 18278 121550 18296
rect 121658 18278 121692 18358
rect 121320 18244 121772 18278
rect 121658 18222 121692 18244
rect 121789 18208 121904 18630
rect 122094 18612 122562 18632
rect 121954 18578 122562 18612
rect 121954 18550 121988 18578
rect 121920 18516 121988 18550
rect 121954 18318 122007 18516
rect 122009 18436 122090 18483
rect 122056 18398 122090 18436
rect 121954 18256 121988 18318
rect 122094 18273 122520 18578
rect 122597 18298 122631 18858
rect 125229 18298 125263 18996
rect 126896 18750 126930 19032
rect 128308 19002 128382 19032
rect 131058 19004 131116 19066
rect 131172 19059 131182 19085
rect 131172 19047 131178 19059
rect 131058 18946 131092 19004
rect 131118 18950 131122 19038
rect 131146 18970 131178 19038
rect 131190 18970 131206 19085
rect 131058 18936 131096 18946
rect 131146 18936 131206 18970
rect 131224 18936 131258 19434
rect 130964 18902 131258 18936
rect 131396 18924 131416 19038
rect 131058 18852 131096 18902
rect 131146 18894 131178 18902
rect 131146 18852 131150 18894
rect 131022 18750 131272 18852
rect 125312 18730 126954 18750
rect 131022 18744 131404 18750
rect 131758 18744 133120 18750
rect 126896 18694 126930 18730
rect 131022 18694 131272 18744
rect 131396 18694 131416 18738
rect 125312 18674 126954 18694
rect 131022 18688 131416 18694
rect 131758 18688 133064 18694
rect 122050 18256 122520 18273
rect 121954 18222 122520 18256
rect 126896 18222 126930 18674
rect 128228 18546 128242 18634
rect 128978 18566 128992 18634
rect 129768 18566 129792 18634
rect 131022 18488 131272 18688
rect 131396 18666 131416 18688
rect 131396 18554 131416 18620
rect 131088 18438 131122 18448
rect 131104 18404 131156 18414
rect 131070 18370 131094 18404
rect 131104 18336 131128 18404
rect 131202 18302 131236 18314
rect 130980 18268 131236 18302
rect 95486 17791 96106 18176
rect 96156 18128 96722 18162
rect 96156 17996 96190 18128
rect 96311 18058 96348 18082
rect 96528 18059 96567 18082
rect 96527 18058 96567 18059
rect 96527 18054 96538 18058
rect 96211 17996 96292 18033
rect 96339 18030 96348 18054
rect 96527 18048 96539 18054
rect 96351 18033 96539 18048
rect 96351 18030 96620 18033
rect 96351 18014 96538 18030
rect 96539 17996 96620 18030
rect 96688 17996 96722 18128
rect 96156 17975 96812 17996
rect 96122 17941 96812 17975
rect 96156 17929 96812 17941
rect 96158 17922 96812 17929
rect 96335 17907 96543 17920
rect 96339 17895 96539 17907
rect 96156 17868 96190 17895
rect 96335 17886 96543 17895
rect 96339 17874 96539 17886
rect 96688 17868 96722 17895
rect 96301 17860 96577 17861
rect 96190 17827 96688 17860
rect 96190 17793 96688 17806
rect 98808 17791 99954 18034
rect 92032 17672 92060 17728
rect 98464 17372 99012 17406
rect 99098 17388 99132 17406
rect 99630 17388 99664 17406
rect 98504 17338 99046 17352
rect 99062 17318 99700 17388
rect 121370 17320 121516 17338
rect 130126 17320 130272 17338
rect 95380 16902 95414 17256
rect 98258 17198 98640 17222
rect 121460 17216 121522 17262
rect 121588 17216 121672 17262
rect 98286 17170 98640 17194
rect 121460 17188 121550 17212
rect 121560 17188 121616 17212
rect 101858 17156 102962 17182
rect 101830 17128 102990 17154
rect 94942 16868 103194 16902
rect 94992 16720 95012 16822
rect 95020 16748 95068 16794
rect 94992 16062 95012 16164
rect 95020 16090 95068 16136
rect 95380 16004 95414 16868
rect 95451 16792 95554 16800
rect 95444 16788 95554 16792
rect 103008 16788 103019 16799
rect 95444 16754 103019 16788
rect 95466 16742 95554 16754
rect 95464 16672 95476 16712
rect 95436 16644 95476 16656
rect 95482 16608 95516 16742
rect 103020 16726 103092 16764
rect 95522 16672 98464 16712
rect 98664 16672 98864 16712
rect 99064 16672 103052 16712
rect 95522 16644 98464 16656
rect 98664 16644 98864 16656
rect 99064 16644 103052 16656
rect 103058 16592 103092 16726
rect 103160 16712 103194 16868
rect 103098 16672 103194 16712
rect 103098 16644 103130 16656
rect 103020 16580 103108 16592
rect 103160 16580 103194 16672
rect 95444 16518 95516 16556
rect 95566 16546 103108 16580
rect 103126 16546 103194 16580
rect 121608 16570 121616 17188
rect 103020 16534 103108 16546
rect 95482 16142 95516 16518
rect 103058 16158 103092 16534
rect 95466 16134 95554 16142
rect 95444 16130 95554 16134
rect 103008 16130 103019 16141
rect 95444 16096 103019 16130
rect 95466 16084 95554 16096
rect 95458 16020 95476 16060
rect 56591 15720 60439 15731
rect 56591 15708 60428 15720
rect 56591 15697 60439 15708
rect 60480 15697 64993 15731
rect 55110 15614 55800 15624
rect 43848 14824 44468 15246
rect 44518 15194 45084 15228
rect 44518 14872 44552 15194
rect 44889 15114 44900 15125
rect 44573 15052 44654 15099
rect 44713 15080 44900 15114
rect 44901 15052 44982 15099
rect 44620 15014 44654 15052
rect 44948 15014 44982 15052
rect 44889 14986 44900 14997
rect 44713 14952 44900 14986
rect 45050 14872 45084 15194
rect 44518 14838 45084 14872
rect 45248 14840 45274 15612
rect 45282 14806 45308 15612
rect 42576 14078 45888 14116
rect 42632 14022 45832 14060
rect 45282 13973 45316 14007
rect 48340 13973 48374 14007
rect 51398 13973 51432 14007
rect 51512 13973 51546 15612
rect 55058 15600 56246 15614
rect 55138 15586 55772 15596
rect 55002 15544 56302 15586
rect 60480 15528 60514 15697
rect 64402 15661 64993 15697
rect 95048 15556 95068 16004
rect 95380 15964 95476 16004
rect 94992 15404 95012 15506
rect 95020 15432 95068 15478
rect 95380 15346 95414 15964
rect 95482 15950 95516 16084
rect 103020 16068 103092 16106
rect 95522 16020 103052 16060
rect 95522 15964 103052 16004
rect 103058 15934 103092 16068
rect 103160 16060 103194 16546
rect 103098 16020 103194 16060
rect 103098 15964 103134 16004
rect 103020 15922 103108 15934
rect 103160 15922 103194 16020
rect 95444 15860 95516 15898
rect 95566 15888 103108 15922
rect 103126 15888 103194 15922
rect 103020 15876 103108 15888
rect 95482 15484 95516 15860
rect 103058 15500 103092 15876
rect 95466 15476 95554 15484
rect 95444 15472 95554 15476
rect 103008 15472 103019 15483
rect 95444 15438 103019 15472
rect 95466 15426 95554 15438
rect 95470 15356 95476 15374
rect 95380 15300 95476 15346
rect 94992 14746 95012 14848
rect 95020 14774 95068 14820
rect 94992 14088 95012 14190
rect 95020 14116 95068 14162
rect 95380 14030 95414 15300
rect 95482 15292 95516 15426
rect 103020 15410 103092 15448
rect 95526 15374 103052 15402
rect 95522 15356 103052 15374
rect 95522 15300 103052 15346
rect 103058 15276 103092 15410
rect 103160 15402 103194 15888
rect 103098 15356 103194 15402
rect 103098 15300 103130 15346
rect 103020 15264 103108 15276
rect 103160 15264 103194 15356
rect 95444 15202 95516 15240
rect 95566 15230 103108 15264
rect 103126 15230 103194 15264
rect 103020 15218 103108 15230
rect 95482 14826 95516 15202
rect 103058 14842 103092 15218
rect 95466 14818 95554 14826
rect 95444 14814 95554 14818
rect 103008 14814 103019 14825
rect 95444 14780 103019 14814
rect 95466 14768 95554 14780
rect 95482 14634 95516 14768
rect 103020 14752 103092 14790
rect 95582 14698 103052 14738
rect 95526 14642 103052 14682
rect 103058 14618 103092 14752
rect 103160 14738 103194 15230
rect 103098 14698 103194 14738
rect 103098 14642 103118 14682
rect 103020 14606 103108 14618
rect 103160 14606 103194 14698
rect 95444 14544 95516 14582
rect 95566 14572 103108 14606
rect 103126 14572 103194 14606
rect 103020 14560 103108 14572
rect 95482 14168 95516 14544
rect 103058 14184 103092 14560
rect 95466 14160 95554 14168
rect 95444 14156 95554 14160
rect 103008 14156 103019 14167
rect 95444 14122 103019 14156
rect 95466 14110 95554 14122
rect 95470 14046 95476 14058
rect 95380 13990 95476 14030
rect 43619 13939 51889 13973
rect 43619 11396 43653 13939
rect 45282 13859 45316 13939
rect 48340 13859 48374 13939
rect 51398 13859 51432 13939
rect 51512 13859 51546 13939
rect 43674 13797 43755 13844
rect 43814 13825 51546 13859
rect 45269 13813 45270 13814
rect 45270 13812 45271 13813
rect 43721 13229 43755 13797
rect 44980 13784 45036 13798
rect 44980 13728 45036 13742
rect 45270 13213 45271 13214
rect 45269 13212 45270 13213
rect 45282 13201 45316 13825
rect 45328 13813 45329 13814
rect 48327 13813 48328 13814
rect 45327 13812 45328 13813
rect 48328 13812 48329 13813
rect 45327 13213 45328 13214
rect 48328 13213 48329 13214
rect 45328 13212 45329 13213
rect 48327 13212 48328 13213
rect 48340 13201 48374 13825
rect 48386 13813 48387 13814
rect 51385 13813 51386 13814
rect 48385 13812 48386 13813
rect 51386 13812 51387 13813
rect 51114 13294 51170 13300
rect 51114 13238 51170 13244
rect 48385 13213 48386 13214
rect 51386 13213 51387 13214
rect 48386 13212 48387 13213
rect 51385 13212 51386 13213
rect 51398 13201 51432 13825
rect 51512 13201 51546 13825
rect 95380 13834 95414 13990
rect 95482 13976 95516 14110
rect 103020 14094 103092 14132
rect 95522 14046 98998 14058
rect 99198 14046 99398 14058
rect 99598 14046 103052 14058
rect 95522 13990 98998 14030
rect 99198 13990 99398 14030
rect 99598 13990 103052 14030
rect 103058 13960 103092 14094
rect 103098 14046 103152 14058
rect 103098 13990 103124 14030
rect 103020 13948 103108 13960
rect 103160 13948 103194 14572
rect 95566 13917 103108 13948
rect 95566 13914 103123 13917
rect 103126 13914 103194 13948
rect 103020 13902 103123 13914
rect 99458 13834 99464 13872
rect 103160 13834 103194 13914
rect 95380 13800 103632 13834
rect 94992 13430 95012 13532
rect 98820 13508 99174 13532
rect 95020 13458 95068 13504
rect 98792 13480 99174 13504
rect 99458 13490 99464 13800
rect 101296 13548 102456 13574
rect 101324 13520 102428 13546
rect 103160 13446 103194 13800
rect 43674 13139 43755 13186
rect 43814 13167 51546 13201
rect 44980 13161 45084 13162
rect 45269 13155 45270 13156
rect 45270 13154 45271 13155
rect 43721 12571 43755 13139
rect 44980 13105 45028 13106
rect 44980 12636 45036 12640
rect 44980 12580 45036 12584
rect 45270 12555 45271 12556
rect 45269 12554 45270 12555
rect 45282 12543 45316 13167
rect 45328 13155 45329 13156
rect 48327 13155 48328 13156
rect 45327 13154 45328 13155
rect 48328 13154 48329 13155
rect 45327 12555 45328 12556
rect 48328 12555 48329 12556
rect 45328 12554 45329 12555
rect 48327 12554 48328 12555
rect 48340 12543 48374 13167
rect 48386 13155 48387 13156
rect 51385 13155 51386 13156
rect 48385 13154 48386 13155
rect 51386 13154 51387 13155
rect 51114 13116 51170 13140
rect 51114 13060 51170 13084
rect 48385 12555 48386 12556
rect 51386 12555 51387 12556
rect 48386 12554 48387 12555
rect 51385 12554 51386 12555
rect 51398 12543 51432 13167
rect 51512 12543 51546 13167
rect 93276 13076 93320 13426
rect 93332 13076 93376 13426
rect 98944 13350 100252 13384
rect 99038 13316 99546 13330
rect 99596 13314 100234 13350
rect 98998 13015 99032 13033
rect 99512 13015 99546 13033
rect 98962 12979 99582 13015
rect 99728 12979 100102 12992
rect 94937 12945 100800 12979
rect 43674 12481 43755 12528
rect 43814 12509 51546 12543
rect 94952 12526 95572 12945
rect 98962 12944 99582 12945
rect 95622 12911 96156 12930
rect 95656 12896 96154 12911
rect 95622 12871 96188 12877
rect 95622 12868 95656 12871
rect 96154 12868 96188 12871
rect 95588 12865 95690 12868
rect 96120 12865 96222 12868
rect 95588 12862 96222 12865
rect 95588 12831 95656 12862
rect 95779 12850 96031 12854
rect 95767 12831 96043 12850
rect 96120 12831 96222 12862
rect 95622 12574 95656 12831
rect 95993 12816 96004 12819
rect 95801 12801 96009 12816
rect 96016 12801 96124 12808
rect 95677 12754 95758 12801
rect 95801 12797 96124 12801
rect 95817 12782 96004 12797
rect 96005 12790 96124 12797
rect 96005 12780 96086 12790
rect 96005 12762 96096 12780
rect 96005 12754 96086 12762
rect 95724 12716 95758 12754
rect 96052 12716 96086 12754
rect 95993 12688 96004 12699
rect 95817 12654 96004 12688
rect 96154 12574 96188 12831
rect 95622 12540 96188 12574
rect 45269 12497 45270 12498
rect 45270 12496 45271 12497
rect 43721 11913 43755 12481
rect 44980 12476 45036 12478
rect 44980 12420 45036 12422
rect 45270 11897 45271 11898
rect 45269 11896 45270 11897
rect 45282 11885 45316 12509
rect 45328 12497 45329 12498
rect 48327 12497 48328 12498
rect 45327 12496 45328 12497
rect 48328 12496 48329 12497
rect 45327 11897 45328 11898
rect 48328 11897 48329 11898
rect 45328 11896 45329 11897
rect 48327 11896 48328 11897
rect 48340 11885 48374 12509
rect 48386 12497 48387 12498
rect 51385 12497 51386 12498
rect 48385 12496 48386 12497
rect 51386 12496 51387 12497
rect 51114 11974 51170 11990
rect 51114 11918 51170 11934
rect 48385 11897 48386 11898
rect 51386 11897 51387 11898
rect 48386 11896 48387 11897
rect 51385 11896 51386 11897
rect 51398 11885 51432 12509
rect 51512 11885 51546 12509
rect 99414 12281 99436 12570
rect 99442 12281 99492 12542
rect 101802 12300 102774 12306
rect 103173 12281 103207 12883
rect 95357 12247 103627 12281
rect 94996 12139 95012 12241
rect 95024 12167 95068 12213
rect 43674 11823 43755 11870
rect 43814 11851 51546 11885
rect 45269 11839 45270 11840
rect 45270 11838 45271 11839
rect 43721 11396 43755 11823
rect 45282 11455 45316 11851
rect 45328 11839 45329 11840
rect 48327 11839 48328 11840
rect 45327 11838 45328 11839
rect 48328 11838 48329 11839
rect 48340 11455 48374 11851
rect 48386 11839 48387 11840
rect 51385 11839 51386 11840
rect 48385 11838 48386 11839
rect 51386 11838 51387 11839
rect 51114 11750 51170 11752
rect 51398 11455 51432 11851
rect 43801 11443 43802 11444
rect 43802 11442 43803 11443
rect 45254 11396 45301 11443
rect 48312 11396 48359 11443
rect 51370 11396 51417 11443
rect 43619 11362 45301 11396
rect 45344 11362 48359 11396
rect 48402 11362 51417 11396
rect 43619 11294 43653 11362
rect 43721 11294 43755 11362
rect 51512 11294 51546 11851
rect 94996 11481 95012 11583
rect 95024 11509 95068 11555
rect 65052 11334 65110 11396
rect 65112 11334 65170 11336
rect 42206 11260 51546 11294
rect 43619 10517 43653 11260
rect 44104 11248 45036 11260
rect 94996 10823 95012 10925
rect 95024 10851 95068 10897
rect 94996 10165 95012 10267
rect 95024 10193 95068 10239
rect 56078 9680 56998 9684
rect 57268 9680 58188 9684
rect 58578 9672 59498 9684
rect 47858 9630 48496 9666
rect 59746 9664 60666 9684
rect 60906 9660 64458 9684
rect 41360 9596 48496 9630
rect 60872 9626 64492 9630
rect 42780 5370 42782 5672
rect 42836 5426 42838 5672
rect 42894 4896 42928 9444
rect 47260 9406 47294 9596
rect 47362 9530 47396 9580
rect 47406 9528 47426 9534
rect 47434 9528 47452 9562
rect 47504 9532 47656 9554
rect 47488 9528 47656 9532
rect 47672 9530 47706 9580
rect 47324 9494 47426 9528
rect 47430 9520 47464 9528
rect 47434 9510 47454 9520
rect 47488 9510 47744 9528
rect 47434 9494 47744 9510
rect 47406 9488 47426 9494
rect 47430 9486 47634 9494
rect 47434 9474 47634 9486
rect 47436 9460 47454 9474
rect 47442 9452 47476 9460
rect 47442 9406 47476 9440
rect 47774 9406 47808 9596
rect 47260 9372 47808 9406
rect 47858 9318 48496 9596
rect 50784 9554 50984 9566
rect 50756 9526 51012 9538
rect 44410 8902 44444 8936
rect 45168 8902 45202 8936
rect 45926 8902 45960 8936
rect 46684 8902 46718 8936
rect 47442 8902 47476 8936
rect 48200 8902 48234 8936
rect 48958 8902 48992 8936
rect 49716 8902 49750 8936
rect 50474 8902 50508 8936
rect 51232 8902 51266 8936
rect 43642 8868 51990 8902
rect 43642 8840 43676 8868
rect 43642 8766 43710 8840
rect 44410 8788 44444 8868
rect 45168 8788 45202 8868
rect 45926 8788 45960 8868
rect 46684 8788 46718 8868
rect 47442 8788 47476 8868
rect 48200 8788 48234 8868
rect 48958 8788 48992 8868
rect 49716 8788 49750 8868
rect 50474 8788 50508 8868
rect 51232 8788 51266 8868
rect 51804 8788 51815 8799
rect 43642 8764 43732 8766
rect 43642 8738 43778 8764
rect 43642 8726 43784 8738
rect 43642 8656 43732 8726
rect 43738 8656 43784 8726
rect 43790 8656 43812 8766
rect 43828 8754 51815 8788
rect 44397 8742 44398 8743
rect 44398 8741 44399 8742
rect 43642 8208 43710 8656
rect 43744 8208 43778 8656
rect 43642 8118 43732 8208
rect 43738 8158 43784 8208
rect 43738 8146 43760 8158
rect 43762 8146 43784 8158
rect 43790 8118 43812 8208
rect 44398 8142 44399 8143
rect 44397 8141 44398 8142
rect 44410 8130 44444 8754
rect 44456 8742 44457 8743
rect 45155 8742 45156 8743
rect 44455 8741 44456 8742
rect 45156 8741 45157 8742
rect 44455 8142 44456 8143
rect 45156 8142 45157 8143
rect 44456 8141 44457 8142
rect 45155 8141 45156 8142
rect 45168 8130 45202 8754
rect 45214 8742 45215 8743
rect 45913 8742 45914 8743
rect 45213 8741 45214 8742
rect 45914 8741 45915 8742
rect 45213 8142 45214 8143
rect 45914 8142 45915 8143
rect 45214 8141 45215 8142
rect 45913 8141 45914 8142
rect 45926 8130 45960 8754
rect 45972 8742 45973 8743
rect 46671 8742 46672 8743
rect 45971 8741 45972 8742
rect 46672 8741 46673 8742
rect 45971 8142 45972 8143
rect 46672 8142 46673 8143
rect 45972 8141 45973 8142
rect 46671 8141 46672 8142
rect 46684 8130 46718 8754
rect 46730 8742 46731 8743
rect 47429 8742 47430 8743
rect 46729 8741 46730 8742
rect 47430 8741 47431 8742
rect 46729 8142 46730 8143
rect 47430 8142 47431 8143
rect 46730 8141 46731 8142
rect 47429 8141 47430 8142
rect 47442 8130 47476 8754
rect 47488 8742 47489 8743
rect 48187 8742 48188 8743
rect 47487 8741 47488 8742
rect 48188 8741 48189 8742
rect 47487 8142 47488 8143
rect 48188 8142 48189 8143
rect 47488 8141 47489 8142
rect 48187 8141 48188 8142
rect 48200 8130 48234 8754
rect 48246 8742 48247 8743
rect 48945 8742 48946 8743
rect 48245 8741 48246 8742
rect 48946 8741 48947 8742
rect 48245 8142 48246 8143
rect 48946 8142 48947 8143
rect 48246 8141 48247 8142
rect 48945 8141 48946 8142
rect 48958 8130 48992 8754
rect 49004 8742 49005 8743
rect 49703 8742 49704 8743
rect 49003 8741 49004 8742
rect 49704 8741 49705 8742
rect 49003 8142 49004 8143
rect 49704 8142 49705 8143
rect 49004 8141 49005 8142
rect 49703 8141 49704 8142
rect 49716 8130 49750 8754
rect 49762 8742 49763 8743
rect 50461 8742 50462 8743
rect 49761 8741 49762 8742
rect 50462 8741 50463 8742
rect 49761 8142 49762 8143
rect 50462 8142 50463 8143
rect 49762 8141 49763 8142
rect 50461 8141 50462 8142
rect 50474 8130 50508 8754
rect 50520 8742 50521 8743
rect 51219 8742 51220 8743
rect 50519 8741 50520 8742
rect 51220 8741 51221 8742
rect 50519 8142 50520 8143
rect 51220 8142 51221 8143
rect 50520 8141 50521 8142
rect 51219 8141 51220 8142
rect 51232 8130 51266 8754
rect 51278 8742 51279 8743
rect 51277 8741 51278 8742
rect 51816 8726 51888 8764
rect 51854 8158 51888 8726
rect 51277 8142 51278 8143
rect 51278 8141 51279 8142
rect 51804 8130 51815 8141
rect 43642 8108 43710 8118
rect 43642 8106 43732 8108
rect 43642 8080 43778 8106
rect 43642 8068 43784 8080
rect 43642 7950 43732 8068
rect 43642 7448 43710 7950
rect 43738 7922 43784 8068
rect 43744 7500 43784 7922
rect 43762 7488 43784 7500
rect 43790 7460 43812 8108
rect 43828 8096 51815 8130
rect 44397 8084 44398 8085
rect 44398 8083 44399 8084
rect 44398 7484 44399 7485
rect 44397 7483 44398 7484
rect 44410 7472 44444 8096
rect 44456 8084 44457 8085
rect 45155 8084 45156 8085
rect 44455 8083 44456 8084
rect 45156 8083 45157 8084
rect 45168 7490 45202 8096
rect 45214 8084 45215 8085
rect 45913 8084 45914 8085
rect 45213 8083 45214 8084
rect 45914 8083 45915 8084
rect 44455 7484 44456 7485
rect 44456 7483 44457 7484
rect 44518 7472 45202 7490
rect 45213 7484 45214 7485
rect 45914 7484 45915 7485
rect 45214 7483 45215 7484
rect 45913 7483 45914 7484
rect 45926 7472 45960 8096
rect 45972 8084 45973 8085
rect 46671 8084 46672 8085
rect 45971 8083 45972 8084
rect 46672 8083 46673 8084
rect 45971 7484 45972 7485
rect 46672 7484 46673 7485
rect 45972 7483 45973 7484
rect 46671 7483 46672 7484
rect 46684 7472 46718 8096
rect 46730 8084 46731 8085
rect 47429 8084 47430 8085
rect 46729 8083 46730 8084
rect 47430 8083 47431 8084
rect 46729 7484 46730 7485
rect 47430 7484 47431 7485
rect 46730 7483 46731 7484
rect 47429 7483 47430 7484
rect 47442 7472 47476 8096
rect 47488 8084 47489 8085
rect 48187 8084 48188 8085
rect 47487 8083 47488 8084
rect 48188 8083 48189 8084
rect 47487 7484 47488 7485
rect 48188 7484 48189 7485
rect 47488 7483 47489 7484
rect 48187 7483 48188 7484
rect 47664 7472 47986 7474
rect 48200 7472 48234 8096
rect 48246 8084 48247 8085
rect 48945 8084 48946 8085
rect 48245 8083 48246 8084
rect 48946 8083 48947 8084
rect 48245 7484 48246 7485
rect 48946 7484 48947 7485
rect 48246 7483 48247 7484
rect 48945 7483 48946 7484
rect 48958 7472 48992 8096
rect 49004 8084 49005 8085
rect 49703 8084 49704 8085
rect 49003 8083 49004 8084
rect 49704 8083 49705 8084
rect 49003 7484 49004 7485
rect 49704 7484 49705 7485
rect 49004 7483 49005 7484
rect 49703 7483 49704 7484
rect 49716 7472 49750 8096
rect 49762 8084 49763 8085
rect 50461 8084 50462 8085
rect 49761 8083 49762 8084
rect 50462 8083 50463 8084
rect 49761 7484 49762 7485
rect 50462 7484 50463 7485
rect 49762 7483 49763 7484
rect 50461 7483 50462 7484
rect 50474 7472 50508 8096
rect 50520 8084 50521 8085
rect 51219 8084 51220 8085
rect 50519 8083 50520 8084
rect 51220 8083 51221 8084
rect 50519 7484 50520 7485
rect 51220 7484 51221 7485
rect 50520 7483 50521 7484
rect 51219 7483 51220 7484
rect 51232 7472 51266 8096
rect 51278 8084 51279 8085
rect 51277 8083 51278 8084
rect 51816 8068 51888 8106
rect 51854 7500 51888 8068
rect 51277 7484 51278 7485
rect 51278 7483 51279 7484
rect 51804 7472 51815 7483
rect 43642 7422 43778 7448
rect 43642 7410 43784 7422
rect 43642 6790 43710 7410
rect 43744 7346 43784 7410
rect 43790 7346 43812 7450
rect 43828 7438 51815 7472
rect 44397 7426 44398 7427
rect 44398 7425 44399 7426
rect 43744 6898 43778 7346
rect 43744 6842 43784 6898
rect 43762 6830 43784 6842
rect 43790 6802 43812 6898
rect 44398 6826 44399 6827
rect 44397 6825 44398 6826
rect 44410 6814 44444 7438
rect 44456 7426 44457 7427
rect 44455 7425 44456 7426
rect 44518 7416 45202 7438
rect 45214 7426 45215 7427
rect 45913 7426 45914 7427
rect 45213 7425 45214 7426
rect 45914 7425 45915 7426
rect 44624 6958 44946 7416
rect 44455 6826 44456 6827
rect 45156 6826 45157 6827
rect 44456 6825 44457 6826
rect 45155 6825 45156 6826
rect 45168 6814 45202 7416
rect 45213 6826 45214 6827
rect 45914 6826 45915 6827
rect 45214 6825 45215 6826
rect 45913 6825 45914 6826
rect 45926 6814 45960 7438
rect 45972 7426 45973 7427
rect 46671 7426 46672 7427
rect 45971 7425 45972 7426
rect 46672 7425 46673 7426
rect 45971 6826 45972 6827
rect 46672 6826 46673 6827
rect 45972 6825 45973 6826
rect 46671 6825 46672 6826
rect 46684 6814 46718 7438
rect 46730 7426 46731 7427
rect 47429 7426 47430 7427
rect 46729 7425 46730 7426
rect 47430 7425 47431 7426
rect 46729 6826 46730 6827
rect 47430 6826 47431 6827
rect 46730 6825 46731 6826
rect 47429 6825 47430 6826
rect 47442 6814 47476 7438
rect 47488 7426 47489 7427
rect 47487 7425 47488 7426
rect 47664 7230 47986 7438
rect 48187 7426 48188 7427
rect 48188 7425 48189 7426
rect 47516 7018 47986 7230
rect 47664 6966 47986 7018
rect 47487 6826 47488 6827
rect 48188 6826 48189 6827
rect 47488 6825 47489 6826
rect 48187 6825 48188 6826
rect 48200 6814 48234 7438
rect 48246 7426 48247 7427
rect 48945 7426 48946 7427
rect 48245 7425 48246 7426
rect 48946 7425 48947 7426
rect 48245 6826 48246 6827
rect 48946 6826 48947 6827
rect 48246 6825 48247 6826
rect 48945 6825 48946 6826
rect 48958 6814 48992 7438
rect 49004 7426 49005 7427
rect 49703 7426 49704 7427
rect 49003 7425 49004 7426
rect 49704 7425 49705 7426
rect 49003 6826 49004 6827
rect 49704 6826 49705 6827
rect 49004 6825 49005 6826
rect 49703 6825 49704 6826
rect 49716 6814 49750 7438
rect 49762 7426 49763 7427
rect 50461 7426 50462 7427
rect 49761 7425 49762 7426
rect 50462 7425 50463 7426
rect 49761 6826 49762 6827
rect 50462 6826 50463 6827
rect 49762 6825 49763 6826
rect 50461 6825 50462 6826
rect 50474 6814 50508 7438
rect 50520 7426 50521 7427
rect 51219 7426 51220 7427
rect 50519 7425 50520 7426
rect 51220 7425 51221 7426
rect 51232 6882 51266 7438
rect 51278 7426 51279 7427
rect 51277 7425 51278 7426
rect 51816 7410 51888 7448
rect 50519 6826 50520 6827
rect 50520 6825 50521 6826
rect 51198 6820 51222 6854
rect 51226 6820 51266 6882
rect 51854 6842 51888 7410
rect 51277 6826 51278 6827
rect 51278 6825 51279 6826
rect 51232 6814 51266 6820
rect 51804 6814 51815 6825
rect 43642 6764 43778 6790
rect 43642 6752 43784 6764
rect 43642 6132 43710 6752
rect 43744 6682 43784 6752
rect 43790 6682 43812 6792
rect 43828 6780 51815 6814
rect 44397 6768 44398 6769
rect 44398 6767 44399 6768
rect 43744 6234 43778 6682
rect 43744 6184 43784 6234
rect 43762 6172 43784 6184
rect 43790 6144 43812 6234
rect 44398 6168 44399 6169
rect 44397 6167 44398 6168
rect 44410 6156 44444 6780
rect 44456 6768 44457 6769
rect 45155 6768 45156 6769
rect 44455 6767 44456 6768
rect 45156 6767 45157 6768
rect 44455 6168 44456 6169
rect 45156 6168 45157 6169
rect 44456 6167 44457 6168
rect 45155 6167 45156 6168
rect 45168 6156 45202 6780
rect 45214 6768 45215 6769
rect 45913 6768 45914 6769
rect 45213 6767 45214 6768
rect 45914 6767 45915 6768
rect 45213 6168 45214 6169
rect 45914 6168 45915 6169
rect 45214 6167 45215 6168
rect 45913 6167 45914 6168
rect 45926 6156 45960 6780
rect 45972 6768 45973 6769
rect 46671 6768 46672 6769
rect 45971 6767 45972 6768
rect 46672 6767 46673 6768
rect 45971 6168 45972 6169
rect 46672 6168 46673 6169
rect 45972 6167 45973 6168
rect 46671 6167 46672 6168
rect 46684 6156 46718 6780
rect 46730 6768 46731 6769
rect 47429 6768 47430 6769
rect 46729 6767 46730 6768
rect 47430 6767 47431 6768
rect 46729 6168 46730 6169
rect 47430 6168 47431 6169
rect 46730 6167 46731 6168
rect 47429 6167 47430 6168
rect 47442 6156 47476 6780
rect 47488 6768 47489 6769
rect 48187 6768 48188 6769
rect 47487 6767 47488 6768
rect 48188 6767 48189 6768
rect 47487 6168 47488 6169
rect 48188 6168 48189 6169
rect 47488 6167 47489 6168
rect 48187 6167 48188 6168
rect 48200 6156 48234 6780
rect 48246 6768 48247 6769
rect 48945 6768 48946 6769
rect 48245 6767 48246 6768
rect 48946 6767 48947 6768
rect 48245 6168 48246 6169
rect 48946 6168 48947 6169
rect 48246 6167 48247 6168
rect 48945 6167 48946 6168
rect 48958 6156 48992 6780
rect 49004 6768 49005 6769
rect 49703 6768 49704 6769
rect 49003 6767 49004 6768
rect 49704 6767 49705 6768
rect 49003 6168 49004 6169
rect 49704 6168 49705 6169
rect 49004 6167 49005 6168
rect 49703 6167 49704 6168
rect 49716 6156 49750 6780
rect 49762 6768 49763 6769
rect 50461 6768 50462 6769
rect 49761 6767 49762 6768
rect 50462 6767 50463 6768
rect 49761 6168 49762 6169
rect 50462 6168 50463 6169
rect 49762 6167 49763 6168
rect 50461 6167 50462 6168
rect 50474 6156 50508 6780
rect 51232 6774 51266 6780
rect 50520 6768 50521 6769
rect 50519 6767 50520 6768
rect 51198 6718 51222 6774
rect 51226 6690 51266 6774
rect 51278 6768 51279 6769
rect 51277 6767 51278 6768
rect 51816 6752 51888 6790
rect 50519 6168 50520 6169
rect 51220 6168 51221 6169
rect 50520 6167 50521 6168
rect 51219 6167 51220 6168
rect 51232 6156 51266 6690
rect 51854 6184 51888 6752
rect 51912 6234 51914 6514
rect 51940 6206 51942 6486
rect 51277 6168 51278 6169
rect 51278 6167 51279 6168
rect 51804 6156 51815 6167
rect 43642 6106 43778 6132
rect 43642 6094 43784 6106
rect 43642 5446 43710 6094
rect 43744 6030 43784 6094
rect 43790 6030 43812 6134
rect 43828 6122 51815 6156
rect 44397 6110 44398 6111
rect 44398 6109 44399 6110
rect 43744 5582 43778 6030
rect 43744 5526 43784 5582
rect 43762 5514 43784 5526
rect 43790 5486 43812 5582
rect 44398 5510 44399 5511
rect 44397 5509 44398 5510
rect 44410 5498 44444 6122
rect 44456 6110 44457 6111
rect 45155 6110 45156 6111
rect 44455 6109 44456 6110
rect 45156 6109 45157 6110
rect 44455 5510 44456 5511
rect 45156 5510 45157 5511
rect 44456 5509 44457 5510
rect 45155 5509 45156 5510
rect 45168 5498 45202 6122
rect 45214 6110 45215 6111
rect 45913 6110 45914 6111
rect 45213 6109 45214 6110
rect 45914 6109 45915 6110
rect 45213 5510 45214 5511
rect 45914 5510 45915 5511
rect 45214 5509 45215 5510
rect 45913 5509 45914 5510
rect 45926 5498 45960 6122
rect 45972 6110 45973 6111
rect 46671 6110 46672 6111
rect 45971 6109 45972 6110
rect 46672 6109 46673 6110
rect 45971 5510 45972 5511
rect 46672 5510 46673 5511
rect 45972 5509 45973 5510
rect 46671 5509 46672 5510
rect 46684 5498 46718 6122
rect 46730 6110 46731 6111
rect 47429 6110 47430 6111
rect 46729 6109 46730 6110
rect 47430 6109 47431 6110
rect 47442 5764 47476 6122
rect 47488 6110 47489 6111
rect 48187 6110 48188 6111
rect 47487 6109 47488 6110
rect 48188 6109 48189 6110
rect 47498 5764 47946 5918
rect 47398 5706 47946 5764
rect 47398 5616 47518 5706
rect 46729 5510 46730 5511
rect 47430 5510 47431 5511
rect 46730 5509 46731 5510
rect 47429 5509 47430 5510
rect 47442 5498 47476 5616
rect 47487 5510 47488 5511
rect 48188 5510 48189 5511
rect 47488 5509 47489 5510
rect 48187 5509 48188 5510
rect 48200 5498 48234 6122
rect 48246 6110 48247 6111
rect 48945 6110 48946 6111
rect 48245 6109 48246 6110
rect 48946 6109 48947 6110
rect 48245 5510 48246 5511
rect 48946 5510 48947 5511
rect 48246 5509 48247 5510
rect 48945 5509 48946 5510
rect 48958 5498 48992 6122
rect 49004 6110 49005 6111
rect 49703 6110 49704 6111
rect 49003 6109 49004 6110
rect 49704 6109 49705 6110
rect 49003 5510 49004 5511
rect 49704 5510 49705 5511
rect 49004 5509 49005 5510
rect 49703 5509 49704 5510
rect 49716 5498 49750 6122
rect 49762 6110 49763 6111
rect 50461 6110 50462 6111
rect 49761 6109 49762 6110
rect 50462 6109 50463 6110
rect 49761 5510 49762 5511
rect 50462 5510 50463 5511
rect 49762 5509 49763 5510
rect 50461 5509 50462 5510
rect 50474 5498 50508 6122
rect 50520 6110 50521 6111
rect 51219 6110 51220 6111
rect 50519 6109 50520 6110
rect 51220 6109 51221 6110
rect 51232 5574 51266 6122
rect 51278 6110 51279 6111
rect 51277 6109 51278 6110
rect 51816 6094 51888 6132
rect 50519 5510 50520 5511
rect 50520 5509 50521 5510
rect 51198 5504 51224 5546
rect 51226 5504 51266 5574
rect 51854 5526 51888 6094
rect 51912 5582 51920 6030
rect 51940 5554 51948 6058
rect 51277 5510 51278 5511
rect 51278 5509 51279 5510
rect 51232 5498 51266 5504
rect 51804 5498 51815 5509
rect 43828 5464 51815 5498
rect 43642 5384 43686 5446
rect 44410 5384 44444 5464
rect 45168 5384 45202 5464
rect 45926 5384 45960 5464
rect 46684 5384 46718 5464
rect 47442 5384 47476 5464
rect 48200 5384 48234 5464
rect 48958 5384 48992 5464
rect 49716 5384 49750 5464
rect 50474 5384 50508 5464
rect 51232 5458 51266 5464
rect 51198 5410 51224 5458
rect 51226 5384 51266 5458
rect 51956 5384 51990 8868
rect 55644 8672 55812 8786
rect 55644 8616 55856 8672
rect 55736 8524 55856 8616
rect 55796 8496 55814 8520
rect 55792 8192 55814 8496
rect 55830 8360 55938 8486
rect 55830 8230 55852 8360
rect 56018 8058 58326 9496
rect 58596 8052 60904 9490
rect 61086 7784 61120 9444
rect 60552 7472 62202 7784
rect 56766 7288 57088 7428
rect 58276 7288 58598 7462
rect 59798 7288 60120 7464
rect 56766 6956 60120 7288
rect 60546 6964 62202 7472
rect 56766 6926 60006 6956
rect 56692 6920 60006 6926
rect 56692 6756 56860 6920
rect 57040 6350 60006 6920
rect 60552 6346 62202 6964
rect 62638 6348 64288 7786
rect 64742 6346 68092 9666
rect 82892 9564 84406 9578
rect 82626 9512 82650 9548
rect 82604 9502 82650 9512
rect 94996 9507 95012 9609
rect 95024 9535 95068 9581
rect 89776 9446 89846 9492
rect 95357 9461 95391 12247
rect 99414 12216 99436 12247
rect 99442 12216 99492 12247
rect 103065 12223 103111 12247
rect 103071 12219 103105 12223
rect 95514 12201 103012 12205
rect 95502 12179 103028 12201
rect 103037 12195 103139 12218
rect 95502 12173 103139 12179
rect 103024 12167 103139 12173
rect 103173 12167 103207 12247
rect 95536 12161 103105 12167
rect 95412 12105 95493 12152
rect 95536 12139 103121 12161
rect 95552 12133 103121 12139
rect 103139 12133 103241 12167
rect 95644 12127 95678 12133
rect 95446 11602 95453 11618
rect 95418 11574 95453 11590
rect 95459 11561 95493 12105
rect 95644 12099 95650 12122
rect 103024 12121 103121 12133
rect 95499 11602 96778 11618
rect 95499 11574 96750 11590
rect 103071 11577 103105 12121
rect 95443 11549 95540 11561
rect 95752 11549 96406 11570
rect 103012 11555 103023 11560
rect 101802 11549 103024 11555
rect 95443 11546 103024 11549
rect 95443 11543 103023 11546
rect 95443 11522 103028 11543
rect 95443 11521 103105 11522
rect 95502 11515 103139 11521
rect 95752 11509 96902 11515
rect 103024 11509 103139 11515
rect 103173 11509 103207 12133
rect 95536 11503 103105 11509
rect 95412 11487 95493 11494
rect 95412 11482 95527 11487
rect 95412 11459 95493 11482
rect 95536 11481 103121 11503
rect 95552 11475 103121 11481
rect 103139 11475 103241 11509
rect 95412 11454 95499 11459
rect 96248 11456 96902 11475
rect 103024 11463 103121 11475
rect 95412 11447 95493 11454
rect 95459 10903 95493 11447
rect 95842 11438 97244 11456
rect 95814 11410 97272 11428
rect 101344 10950 102752 10968
rect 101372 10922 102724 10940
rect 103071 10924 103105 11463
rect 103065 10907 103111 10924
rect 95443 10891 95540 10903
rect 103012 10891 103023 10902
rect 95443 10885 103023 10891
rect 95443 10864 103028 10885
rect 103037 10879 103139 10896
rect 95443 10863 103105 10864
rect 95502 10857 103139 10863
rect 103024 10851 103139 10857
rect 103173 10851 103207 11475
rect 115190 10896 115191 16570
rect 121664 16514 121672 17216
rect 121674 12328 122380 12364
rect 122477 12328 122511 17257
rect 130216 17216 130278 17262
rect 130344 17216 130428 17262
rect 130216 17188 130306 17212
rect 130316 17188 130372 17212
rect 130420 16514 130428 17216
rect 128286 12554 128292 12754
rect 128314 12526 128320 12782
rect 121674 12294 123076 12328
rect 95536 10845 103105 10851
rect 95412 10789 95493 10836
rect 95536 10823 103121 10845
rect 95552 10817 103121 10823
rect 103139 10817 103241 10851
rect 103024 10805 103121 10817
rect 95446 10280 95453 10298
rect 95418 10252 95453 10270
rect 95459 10245 95493 10789
rect 101888 10768 103065 10786
rect 101860 10740 103065 10758
rect 95499 10280 96756 10298
rect 95499 10252 96728 10270
rect 103071 10261 103105 10805
rect 103111 10768 103152 10786
rect 103111 10740 103124 10758
rect 95443 10233 95540 10245
rect 95732 10233 96386 10252
rect 103012 10233 103023 10244
rect 95443 10227 103023 10233
rect 95443 10206 103028 10227
rect 95443 10205 103105 10206
rect 95502 10199 103139 10205
rect 95732 10193 96922 10199
rect 103024 10193 103139 10199
rect 103173 10193 103207 10817
rect 95536 10187 103105 10193
rect 95412 10171 95493 10178
rect 95412 10162 95527 10171
rect 95536 10165 103121 10187
rect 95412 10143 95493 10162
rect 95552 10159 103121 10165
rect 103139 10159 103241 10193
rect 95412 10134 95499 10143
rect 96268 10138 96922 10159
rect 101286 10153 102750 10159
rect 103024 10147 103121 10159
rect 95412 10131 95493 10134
rect 95459 9587 95493 10131
rect 95864 10118 97266 10134
rect 95836 10090 97294 10106
rect 103071 9614 103105 10147
rect 103065 9591 103111 9614
rect 95443 9575 95540 9587
rect 103012 9575 103023 9586
rect 95443 9569 103023 9575
rect 95443 9547 103028 9569
rect 103037 9563 103139 9586
rect 95502 9541 103028 9547
rect 95536 9507 103062 9535
rect 95552 9503 103050 9507
rect 95459 9473 95493 9495
rect 103173 9461 103207 10159
rect 89776 9418 89790 9440
rect 94937 9427 103207 9461
rect 115190 9494 115218 10896
rect 85670 8862 85942 8866
rect 82654 8848 88986 8862
rect 85654 8846 85954 8848
rect 85654 8842 85952 8846
rect 82682 8814 88986 8834
rect 95357 8825 95391 9427
rect 101826 9402 102750 9408
rect 115190 9185 115191 9494
rect 116430 9472 116446 10874
rect 115151 9182 115191 9185
rect 115145 9170 115191 9182
rect 119966 8974 120904 11342
rect 121674 10126 122380 12294
rect 122477 12214 122511 12294
rect 122591 12214 122625 12294
rect 122881 12214 122892 12225
rect 122443 12180 122892 12214
rect 122477 11556 122511 12180
rect 122591 12150 122625 12180
rect 122637 12168 122638 12169
rect 122636 12167 122637 12168
rect 122893 12152 122974 12199
rect 122591 12120 122631 12150
rect 122650 12148 122659 12150
rect 122591 11556 122625 12120
rect 122940 11584 122974 12152
rect 122636 11568 122637 11569
rect 122637 11567 122638 11568
rect 122881 11556 122892 11567
rect 122443 11522 122892 11556
rect 122477 10898 122511 11522
rect 122591 10898 122625 11522
rect 122637 11510 122638 11511
rect 122636 11509 122637 11510
rect 122893 11494 122974 11541
rect 122940 10926 122974 11494
rect 122636 10910 122637 10911
rect 122637 10909 122638 10910
rect 122881 10898 122892 10909
rect 122443 10864 122892 10898
rect 122477 10240 122511 10864
rect 122591 10542 122625 10864
rect 122637 10852 122638 10853
rect 122636 10851 122637 10852
rect 122893 10836 122974 10883
rect 122940 10542 122974 10836
rect 122591 10320 122636 10542
rect 122940 10365 123021 10542
rect 122893 10352 123021 10365
rect 123042 10352 123076 12294
rect 123260 11348 124680 12340
rect 130260 11440 130284 11640
rect 130288 11412 130312 11668
rect 123718 11196 123848 11216
rect 124572 11150 124599 11182
rect 122591 10240 122625 10320
rect 122764 10318 123154 10352
rect 122636 10252 122637 10253
rect 122637 10251 122638 10252
rect 122764 10240 122798 10318
rect 122940 10252 122974 10318
rect 122881 10240 122892 10251
rect 122978 10250 123025 10297
rect 122443 10206 122897 10240
rect 122924 10218 123025 10250
rect 122924 10216 122931 10218
rect 122940 10216 123025 10218
rect 122477 10126 122511 10206
rect 122591 10126 122625 10206
rect 122764 10126 122798 10206
rect 122878 10168 122912 10173
rect 123008 10168 123040 10173
rect 122867 10157 122912 10168
rect 122995 10157 123040 10168
rect 122878 10126 122912 10157
rect 123006 10126 123040 10157
rect 123042 10126 123076 10318
rect 121674 10092 123076 10126
rect 121674 10056 122380 10092
rect 121668 9750 122380 9786
rect 122477 9750 122511 10092
rect 122764 9820 122798 10092
rect 122878 9981 122912 10092
rect 123006 9981 123040 10092
rect 122978 9922 123025 9969
rect 122940 9888 123025 9922
rect 123120 9820 123154 10318
rect 123260 10158 124680 11150
rect 130260 11040 130284 11240
rect 130288 11012 130312 11268
rect 123886 9898 123960 10158
rect 124572 10114 124599 10158
rect 124606 10148 124633 10158
rect 125223 9840 125257 9878
rect 122764 9786 123154 9820
rect 121668 9736 123070 9750
rect 121668 9716 123168 9736
rect 121668 8974 122380 9716
rect 122477 9636 122511 9716
rect 122591 9636 122625 9716
rect 122746 9636 123168 9716
rect 122443 9602 123168 9636
rect 122477 9021 122511 9602
rect 122591 9192 122625 9602
rect 122637 9590 122638 9591
rect 122636 9589 122637 9590
rect 122591 9182 122636 9192
rect 122746 9170 123168 9602
rect 122606 9123 123168 9170
rect 122653 9116 123168 9123
rect 122653 9089 123070 9116
rect 122934 9021 122968 9089
rect 123036 9021 123070 9089
rect 123252 9021 125272 9840
rect 122477 8987 125272 9021
rect 82682 8792 85654 8814
rect 85954 8792 88986 8814
rect 98446 8763 99066 8764
rect 95453 8729 100800 8763
rect 97474 8724 97586 8729
rect 98446 8693 99066 8729
rect 99212 8716 99586 8729
rect 82472 8644 83472 8648
rect 83908 8644 85558 8646
rect 86012 8644 89636 8648
rect 82034 8484 82618 8510
rect 82034 8476 82602 8484
rect 80468 8422 80474 8425
rect 80468 8236 80494 8422
rect 82602 8278 82624 8420
rect 83254 8406 83266 8408
rect 83282 8378 83294 8408
rect 80468 7925 80474 8236
rect 82602 8156 83234 8278
rect 83402 8260 83436 8516
rect 82614 7856 83234 8156
rect 83284 8226 83334 8260
rect 83380 8226 83754 8260
rect 83284 8154 83318 8226
rect 83284 7978 83328 8154
rect 83332 8006 83356 8126
rect 83402 8118 83436 8226
rect 83467 8146 83490 8158
rect 83402 8046 83454 8118
rect 83463 8112 83490 8146
rect 83467 8100 83490 8112
rect 83284 7904 83318 7978
rect 83402 7904 83436 8046
rect 83467 8018 83490 8030
rect 83463 7984 83490 8018
rect 83467 7972 83490 7984
rect 83284 7870 83334 7904
rect 83380 7870 83754 7904
rect 83402 7342 83436 7870
rect 83908 7834 84140 8550
rect 82095 7210 83472 7295
rect 83908 7208 85558 7295
rect 76960 6990 77134 7022
rect 76994 6956 77168 6988
rect 77270 6936 77294 6954
rect 77270 6900 77330 6936
rect 77288 6888 77348 6900
rect 77288 6852 77330 6888
rect 68150 6556 68172 6752
rect 77324 6072 77358 6804
rect 80718 6508 80740 6718
rect 79926 6168 79936 6222
rect 80042 6168 80050 6202
rect 82104 6168 82138 6810
rect 82349 6204 82428 7041
rect 86048 7005 86082 8516
rect 89566 7005 89600 8516
rect 82481 6971 90655 7005
rect 86048 6891 86082 6971
rect 86162 6891 86196 6971
rect 86820 6891 86854 6971
rect 87478 6891 87512 6971
rect 88136 6891 88170 6971
rect 88794 6891 88828 6971
rect 89452 6891 89486 6971
rect 89566 6891 89600 6971
rect 82453 6644 82466 6879
rect 86014 6857 89600 6891
rect 82487 6644 82500 6845
rect 82544 6261 82564 6267
rect 82540 6211 82564 6261
rect 82385 6168 82419 6204
rect 82453 6188 82564 6211
rect 82568 6202 82592 6239
rect 86048 6233 86082 6857
rect 86162 6233 86196 6857
rect 86208 6845 86209 6846
rect 86807 6845 86808 6846
rect 86207 6844 86208 6845
rect 86808 6844 86809 6845
rect 86207 6245 86208 6246
rect 86808 6245 86809 6246
rect 86208 6244 86209 6245
rect 86807 6244 86808 6245
rect 86820 6233 86854 6857
rect 86866 6845 86867 6846
rect 87465 6845 87466 6846
rect 86865 6844 86866 6845
rect 87466 6844 87467 6845
rect 86865 6245 86866 6246
rect 87466 6245 87467 6246
rect 86866 6244 86867 6245
rect 87465 6244 87466 6245
rect 87478 6233 87512 6857
rect 87524 6845 87525 6846
rect 88123 6845 88124 6846
rect 87523 6844 87524 6845
rect 88124 6844 88125 6845
rect 87523 6245 87524 6246
rect 88124 6245 88125 6246
rect 87524 6244 87525 6245
rect 88123 6244 88124 6245
rect 88136 6233 88170 6857
rect 88182 6845 88183 6846
rect 88781 6845 88782 6846
rect 88181 6844 88182 6845
rect 88782 6844 88783 6845
rect 88181 6245 88182 6246
rect 88782 6245 88783 6246
rect 88182 6244 88183 6245
rect 88781 6244 88782 6245
rect 88794 6233 88828 6857
rect 88840 6845 88841 6846
rect 89439 6845 89440 6846
rect 88839 6844 88840 6845
rect 89440 6844 89441 6845
rect 88839 6245 88840 6246
rect 89440 6245 89441 6246
rect 88840 6244 88841 6245
rect 89439 6244 89440 6245
rect 89452 6233 89486 6857
rect 89566 6233 89600 6857
rect 90581 6774 90588 6869
rect 90609 6774 90616 6841
rect 100800 6444 103026 6478
rect 82568 6199 83470 6202
rect 86014 6199 89600 6233
rect 90581 6221 90588 6326
rect 90609 6249 90616 6326
rect 99672 6229 103137 6240
rect 99672 6217 103126 6229
rect 82568 6193 82592 6199
rect 82487 6183 82521 6188
rect 82481 6168 82527 6183
rect 77876 6132 79454 6166
rect 76500 6026 76546 6032
rect 76612 6026 76654 6032
rect 76500 5998 76574 6004
rect 76584 5998 76654 6004
rect 76496 5830 76642 5982
rect 76550 5726 76604 5830
rect 77324 5630 77368 6072
rect 43642 5350 51990 5384
rect 77334 5350 77368 5630
rect 77876 5568 77910 6132
rect 78005 6064 78260 6111
rect 78620 6064 78667 6111
rect 78012 5996 78036 6064
rect 78040 6030 78667 6064
rect 78040 6024 78064 6030
rect 78084 5983 78142 6030
rect 78670 5996 78688 6098
rect 78754 6080 78801 6111
rect 78698 6064 78716 6070
rect 78742 6064 78801 6080
rect 79278 6064 79325 6111
rect 78698 6030 79325 6064
rect 78698 6028 78716 6030
rect 78742 6028 78800 6030
rect 78698 6024 78800 6028
rect 78742 6000 78800 6024
rect 78718 5996 78800 6000
rect 77979 5971 78035 5982
rect 77990 5717 78035 5971
rect 78096 5729 78141 5983
rect 78637 5971 78682 5982
rect 78648 5717 78682 5971
rect 78690 5802 78712 5978
rect 78718 5774 78740 5996
rect 78742 5983 78800 5996
rect 78754 5729 78788 5983
rect 79295 5971 79340 5982
rect 79306 5717 79340 5971
rect 77978 5670 78260 5717
rect 78636 5670 78695 5717
rect 78726 5676 78773 5717
rect 78714 5670 78773 5676
rect 79294 5670 79352 5717
rect 77978 5636 78115 5670
rect 78158 5636 78773 5670
rect 78816 5636 79352 5670
rect 79386 5636 79400 5670
rect 77978 5620 78036 5636
rect 78060 5630 78080 5636
rect 77978 5605 77993 5620
rect 78088 5602 78108 5636
rect 78636 5620 78694 5636
rect 78714 5630 78738 5636
rect 78742 5602 78766 5636
rect 79294 5620 79352 5636
rect 79337 5605 79352 5620
rect 77990 5568 78024 5602
rect 78648 5568 78682 5602
rect 79306 5568 79340 5602
rect 79420 5568 79454 6132
rect 79980 6112 79990 6168
rect 80004 6134 83532 6168
rect 80004 6112 80014 6134
rect 79980 5574 80014 6112
rect 80016 5719 80048 6112
rect 80674 6082 80721 6113
rect 80662 6072 80721 6082
rect 80724 6072 80771 6113
rect 81332 6082 81379 6113
rect 80662 6066 80771 6072
rect 81320 6066 81379 6082
rect 81382 6066 81429 6113
rect 81990 6082 82036 6113
rect 82104 6100 82138 6134
rect 81978 6066 82036 6082
rect 82096 6066 82138 6100
rect 80156 6032 80771 6066
rect 80814 6032 81429 6066
rect 81472 6032 82036 6066
rect 80662 6026 80736 6032
rect 80060 5984 80084 6013
rect 80662 5985 80720 6026
rect 81320 5985 81378 6032
rect 81978 5985 82036 6032
rect 82040 6032 82058 6066
rect 82040 6026 82052 6032
rect 82104 6007 82110 6039
rect 82114 6007 82138 6066
rect 82104 5996 82138 6007
rect 80088 5984 80112 5985
rect 80060 5973 80128 5984
rect 80060 5730 80084 5973
rect 80088 5723 80128 5973
rect 80674 5766 80714 5985
rect 80741 5980 80786 5984
rect 80724 5973 80786 5980
rect 80724 5794 80742 5973
rect 80674 5735 80708 5766
rect 80752 5723 80786 5973
rect 81332 5735 81366 5985
rect 81399 5973 81444 5984
rect 81410 5723 81444 5973
rect 81990 5735 82024 5985
rect 82040 5973 82138 5996
rect 82040 5970 82102 5973
rect 80082 5676 80141 5723
rect 80646 5676 80693 5723
rect 80740 5676 80799 5723
rect 81304 5676 81351 5723
rect 81398 5676 81457 5723
rect 81962 5676 82009 5723
rect 80082 5642 80693 5676
rect 80736 5642 81351 5676
rect 81394 5642 82009 5676
rect 80082 5626 80140 5642
rect 80740 5626 80798 5642
rect 81398 5626 81456 5642
rect 80082 5611 80097 5626
rect 80094 5574 80128 5608
rect 80752 5574 80786 5608
rect 80788 5574 80792 5626
rect 81410 5574 81444 5608
rect 82034 5574 82040 5774
rect 82062 5574 82096 5774
rect 82104 5574 82138 5973
rect 77420 5534 79464 5568
rect 79980 5540 82138 5574
rect 82385 6066 82419 6134
rect 82453 6066 82466 6112
rect 82487 6066 82521 6134
rect 82698 6066 82745 6113
rect 83356 6066 83403 6113
rect 82385 6032 82745 6066
rect 82788 6032 83403 6066
rect 77876 5430 77910 5534
rect 77770 5410 78432 5430
rect 77812 5390 78378 5410
rect 77876 5386 77910 5390
rect 77840 5362 78378 5386
rect 77876 5350 77910 5362
rect 79420 5350 79454 5534
rect 79980 5358 80014 5540
rect 80788 5358 80792 5540
rect 43652 5240 43686 5350
rect 43652 5154 43752 5240
rect 43652 4896 43686 5154
rect 44286 5048 44294 5078
rect 44314 5076 44322 5078
rect 44376 5076 44400 5078
rect 44404 5048 44428 5078
rect 43784 4878 44332 4912
rect 43784 4850 43818 4878
rect 44298 4850 44332 4878
rect 43750 4846 43852 4850
rect 44264 4846 44366 4850
rect 43784 4744 43818 4846
rect 43824 4844 44332 4846
rect 43932 4832 44184 4836
rect 43920 4812 44196 4832
rect 44298 4812 44332 4844
rect 43828 4810 43978 4812
rect 44138 4810 44332 4812
rect 43828 4806 44332 4810
rect 43828 4796 44288 4806
rect 43886 4744 43920 4770
rect 43954 4764 44162 4796
rect 44192 4778 44282 4784
rect 44196 4744 44230 4770
rect 44298 4744 44332 4806
rect 44382 4744 45020 4966
rect 77312 4766 77404 5350
rect 77840 4954 78304 5350
rect 77840 4764 78318 4954
rect 78322 4902 78378 4920
rect 78432 4902 78484 4920
rect 41360 4722 45020 4744
rect 41360 4721 43936 4722
rect 41360 4720 43947 4721
rect 43958 4720 45020 4722
rect 41360 4710 45020 4720
rect 43784 4658 43818 4710
rect 44298 4658 44332 4710
rect 44382 4674 45020 4710
rect 53462 4314 56054 4394
rect 78280 4322 78318 4764
rect 78340 4382 78378 4894
rect 78432 4874 78456 4892
rect 78502 4764 79490 5350
rect 53394 3756 56054 4314
rect 53462 3500 56054 3756
rect 79944 3338 80804 5358
rect 80980 3346 81972 5366
rect 80120 3168 80134 3338
rect 80148 3196 80162 3338
rect 79478 1830 79504 2754
rect 79512 1830 79538 2720
rect 80788 2000 80792 3338
rect 81410 3332 81444 3346
rect 81314 3238 81648 3332
rect 81314 3154 81878 3238
rect 80752 1997 80792 2000
rect 81410 1997 81444 3154
rect 82034 2184 82040 5540
rect 82062 2184 82096 5540
rect 82385 5370 82419 6032
rect 82453 5560 82466 6032
rect 82487 5603 82521 6032
rect 82568 5985 82569 5986
rect 82567 5984 82568 5985
rect 82715 5973 82760 5984
rect 83373 5973 83418 5984
rect 82487 5587 82500 5603
rect 82714 5587 82715 5588
rect 82713 5586 82714 5587
rect 82726 5575 82760 5973
rect 82771 5587 82772 5588
rect 83372 5587 83373 5588
rect 82772 5586 82773 5587
rect 83371 5586 83372 5587
rect 83384 5575 83418 5973
rect 83498 5575 83532 6134
rect 86048 5575 86082 6199
rect 86162 5575 86196 6199
rect 86208 6187 86209 6188
rect 86807 6187 86808 6188
rect 86207 6186 86208 6187
rect 86808 6186 86809 6187
rect 86207 5587 86208 5588
rect 86808 5587 86809 5588
rect 86208 5586 86209 5587
rect 86807 5586 86808 5587
rect 86820 5575 86854 6199
rect 86866 6187 86867 6188
rect 87465 6187 87466 6188
rect 86865 6186 86866 6187
rect 87466 6186 87467 6187
rect 86865 5587 86866 5588
rect 87466 5587 87467 5588
rect 86866 5586 86867 5587
rect 87465 5586 87466 5587
rect 87478 5575 87512 6199
rect 87524 6187 87525 6188
rect 88123 6187 88124 6188
rect 87523 6186 87524 6187
rect 88124 6186 88125 6187
rect 87523 5587 87524 5588
rect 88124 5587 88125 5588
rect 87524 5586 87525 5587
rect 88123 5586 88124 5587
rect 88136 5575 88170 6199
rect 88182 6187 88183 6188
rect 88781 6187 88782 6188
rect 88181 6186 88182 6187
rect 88782 6186 88783 6187
rect 88181 5587 88182 5588
rect 88782 5587 88783 5588
rect 88182 5586 88183 5587
rect 88781 5586 88782 5587
rect 88794 5575 88828 6199
rect 88840 6187 88841 6188
rect 89439 6187 89440 6188
rect 88839 6186 88840 6187
rect 89440 6186 89441 6187
rect 88839 5587 88840 5588
rect 89440 5587 89441 5588
rect 88840 5586 88841 5587
rect 89439 5586 89440 5587
rect 89452 5575 89486 6199
rect 89566 5575 89600 6199
rect 90581 6116 90588 6211
rect 99672 6206 103137 6217
rect 90609 6116 90616 6183
rect 99672 5820 99706 6206
rect 100416 6138 100454 6176
rect 101074 6138 101112 6176
rect 101732 6138 101770 6176
rect 102390 6138 102428 6176
rect 103076 6172 103086 6176
rect 99848 6104 100454 6138
rect 100506 6104 101112 6138
rect 101164 6104 101770 6138
rect 101822 6104 102428 6138
rect 102480 6104 103064 6138
rect 103076 6070 103098 6172
rect 103178 6144 103212 7812
rect 122268 7664 122380 7668
rect 123036 7610 123070 8987
rect 123252 8951 125272 8987
rect 123456 7398 123862 7402
rect 120134 7038 120140 7084
rect 120162 7010 120168 7084
rect 120184 7034 120336 7088
rect 120362 7034 120454 7050
rect 120184 7028 120454 7034
rect 120134 6930 120140 6972
rect 120162 6930 120168 7000
rect 120184 6980 120440 7028
rect 120184 6942 120336 6980
rect 124368 6664 125622 6672
rect 119362 6250 120536 6260
rect 120816 6250 121400 6272
rect 119362 6226 121400 6250
rect 120094 6216 121400 6226
rect 120816 6180 121400 6216
rect 103037 6066 103038 6067
rect 103076 6066 103086 6070
rect 103038 6065 103039 6066
rect 99775 6054 99820 6065
rect 100433 6054 100478 6065
rect 101091 6054 101136 6065
rect 101749 6056 101794 6065
rect 99786 5820 99820 6054
rect 99831 5832 99832 5833
rect 100432 5832 100433 5833
rect 99832 5831 99833 5832
rect 100431 5831 100432 5832
rect 100444 5820 100478 6054
rect 100489 5832 100490 5833
rect 101090 5832 101091 5833
rect 100490 5831 100491 5832
rect 101089 5831 101090 5832
rect 101102 5820 101136 6054
rect 101734 5844 101814 6056
rect 102407 6054 102452 6065
rect 101147 5832 101148 5833
rect 101148 5831 101149 5832
rect 101610 5820 102068 5844
rect 102406 5832 102407 5833
rect 102405 5831 102406 5832
rect 102418 5820 102452 6054
rect 103064 5854 103122 6066
rect 102463 5832 102464 5833
rect 103046 5832 103122 5854
rect 102464 5831 102465 5832
rect 103026 5826 103037 5831
rect 103018 5820 103038 5826
rect 99672 5786 103038 5820
rect 82440 5513 82521 5560
rect 82580 5541 83532 5575
rect 86014 5541 89600 5575
rect 90581 5563 90588 5668
rect 90609 5591 90616 5668
rect 82713 5529 82714 5530
rect 82714 5528 82715 5529
rect 82453 5478 82466 5513
rect 82487 5370 82521 5513
rect 82726 5370 82760 5541
rect 82772 5529 82773 5530
rect 83371 5529 83372 5530
rect 82771 5528 82772 5529
rect 83372 5528 83373 5529
rect 83318 5508 83378 5510
rect 83384 5370 83418 5541
rect 83498 5510 83532 5541
rect 83424 5508 83590 5510
rect 83498 5370 83532 5508
rect 82140 4259 85764 5370
rect 86048 4917 86082 5541
rect 86162 4917 86196 5541
rect 86208 5529 86209 5530
rect 86807 5529 86808 5530
rect 86207 5528 86208 5529
rect 86808 5528 86809 5529
rect 86207 4929 86208 4930
rect 86808 4929 86809 4930
rect 86208 4928 86209 4929
rect 86807 4928 86808 4929
rect 86820 4917 86854 5541
rect 86866 5529 86867 5530
rect 87465 5529 87466 5530
rect 86865 5528 86866 5529
rect 87466 5528 87467 5529
rect 86856 4923 86860 5006
rect 86865 4929 86866 4930
rect 87466 4929 87467 4930
rect 86866 4928 86867 4929
rect 87465 4928 87466 4929
rect 87478 4917 87512 5541
rect 87524 5529 87525 5530
rect 88123 5529 88124 5530
rect 87523 5528 87524 5529
rect 88124 5528 88125 5529
rect 87523 4929 87524 4930
rect 88124 4929 88125 4930
rect 87524 4928 87525 4929
rect 88123 4928 88124 4929
rect 88136 4917 88170 5541
rect 88182 5529 88183 5530
rect 88781 5529 88782 5530
rect 88181 5528 88182 5529
rect 88782 5528 88783 5529
rect 88181 4929 88182 4930
rect 88782 4929 88783 4930
rect 88182 4928 88183 4929
rect 88781 4928 88782 4929
rect 88794 4917 88828 5541
rect 88840 5529 88841 5530
rect 89439 5529 89440 5530
rect 88839 5528 88840 5529
rect 89440 5528 89441 5529
rect 88839 4929 88840 4930
rect 89440 4929 89441 4930
rect 88840 4928 88841 4929
rect 89439 4928 89440 4929
rect 89452 4917 89486 5541
rect 89566 4917 89600 5541
rect 90581 5454 90588 5553
rect 90609 5454 90616 5525
rect 95248 5240 96080 5254
rect 94982 5202 95006 5224
rect 94960 5178 95006 5202
rect 99672 5162 99706 5786
rect 99786 5162 99820 5786
rect 99832 5774 99833 5775
rect 100431 5774 100432 5775
rect 99831 5773 99832 5774
rect 100432 5773 100433 5774
rect 99831 5174 99832 5175
rect 100432 5174 100433 5175
rect 99832 5173 99833 5174
rect 100431 5173 100432 5174
rect 100444 5162 100478 5786
rect 100490 5774 100491 5775
rect 101089 5774 101090 5775
rect 100489 5773 100490 5774
rect 101090 5773 101091 5774
rect 100489 5174 100490 5175
rect 101090 5174 101091 5175
rect 100490 5173 100491 5174
rect 101089 5173 101090 5174
rect 101102 5162 101136 5786
rect 101148 5774 101149 5775
rect 101147 5773 101148 5774
rect 101610 5752 102068 5786
rect 102405 5774 102406 5775
rect 102406 5773 102407 5774
rect 101147 5174 101148 5175
rect 101748 5174 101749 5175
rect 101148 5173 101149 5174
rect 101747 5173 101748 5174
rect 101760 5162 101794 5752
rect 101805 5174 101806 5175
rect 102406 5174 102407 5175
rect 101806 5173 101807 5174
rect 102405 5173 102406 5174
rect 102418 5162 102452 5786
rect 103018 5780 103038 5786
rect 102464 5774 102465 5775
rect 103046 5774 103066 5832
rect 103107 5817 103122 5832
rect 103107 5774 103122 5789
rect 102463 5773 102464 5774
rect 103046 5752 103122 5774
rect 102463 5174 102464 5175
rect 103064 5174 103122 5752
rect 102464 5173 102465 5174
rect 103026 5162 103037 5173
rect 99672 5128 103037 5162
rect 103070 5146 103094 5174
rect 103107 5159 103122 5174
rect 96024 5090 96136 5092
rect 86014 4883 89600 4917
rect 86048 4280 86082 4883
rect 86162 4441 86196 4883
rect 86208 4871 86209 4872
rect 86807 4871 86808 4872
rect 86207 4870 86208 4871
rect 86808 4870 86809 4871
rect 86820 4441 86854 4883
rect 86856 4784 86860 4877
rect 86866 4871 86867 4872
rect 87465 4871 87466 4872
rect 86865 4870 86866 4871
rect 87466 4870 87467 4871
rect 87478 4492 87512 4883
rect 87524 4871 87525 4872
rect 88123 4871 88124 4872
rect 87523 4870 87524 4871
rect 88124 4870 88125 4871
rect 88136 4492 88170 4883
rect 88182 4871 88183 4872
rect 88781 4871 88782 4872
rect 88181 4870 88182 4871
rect 88782 4870 88783 4871
rect 88794 4492 88828 4883
rect 88840 4871 88841 4872
rect 89439 4871 89440 4872
rect 88839 4870 88840 4871
rect 89440 4870 89441 4871
rect 89452 4492 89486 4883
rect 87478 4441 87523 4492
rect 88136 4441 88181 4492
rect 88794 4441 88839 4492
rect 89452 4441 89497 4492
rect 86792 4382 86839 4429
rect 87426 4382 89471 4429
rect 86224 4348 86839 4382
rect 86882 4348 87497 4382
rect 87540 4348 88155 4382
rect 88198 4348 88813 4382
rect 88856 4348 89471 4382
rect 86144 4280 89504 4293
rect 89566 4280 89600 4883
rect 98810 4694 99144 4872
rect 97344 4618 98264 4652
rect 97344 4504 97378 4618
rect 98088 4550 98126 4588
rect 97520 4538 98126 4550
rect 97504 4516 98126 4538
rect 97504 4504 98104 4516
rect 98230 4504 98264 4618
rect 98512 4610 99432 4644
rect 98512 4504 98546 4610
rect 99256 4542 99294 4580
rect 98688 4538 99294 4542
rect 98672 4508 99294 4538
rect 98672 4504 99272 4508
rect 99398 4504 99432 4610
rect 99672 4504 99706 5128
rect 99786 4504 99820 5128
rect 99832 5116 99833 5117
rect 100431 5116 100432 5117
rect 99831 5115 99832 5116
rect 100432 5115 100433 5116
rect 99831 4516 99832 4517
rect 100432 4516 100433 4517
rect 99832 4515 99833 4516
rect 100431 4515 100432 4516
rect 100444 4504 100478 5128
rect 100490 5116 100491 5117
rect 101089 5116 101090 5117
rect 100489 5115 100490 5116
rect 101090 5115 101091 5116
rect 100489 4516 100490 4517
rect 101090 4516 101091 4517
rect 100490 4515 100491 4516
rect 101089 4515 101090 4516
rect 101102 4504 101136 5128
rect 101148 5116 101149 5117
rect 101747 5116 101748 5117
rect 101147 5115 101148 5116
rect 101748 5115 101749 5116
rect 101147 4516 101148 4517
rect 101748 4516 101749 4517
rect 101148 4515 101149 4516
rect 101747 4515 101748 4516
rect 101760 4504 101794 5128
rect 101806 5116 101807 5117
rect 102405 5116 102406 5117
rect 101805 5115 101806 5116
rect 102406 5115 102407 5116
rect 101805 4516 101806 4517
rect 102406 4516 102407 4517
rect 101806 4515 101807 4516
rect 102405 4515 102406 4516
rect 102418 4504 102452 5128
rect 102464 5116 102465 5117
rect 103107 5116 103122 5131
rect 102463 5115 102464 5116
rect 102463 4516 102464 4517
rect 103064 4516 103122 5116
rect 102464 4515 102465 4516
rect 103026 4504 103037 4515
rect 95050 4470 103037 4504
rect 103107 4501 103122 4516
rect 86048 4259 89600 4280
rect 90577 4259 90586 4398
rect 90615 4287 90624 4436
rect 96298 4390 96680 4470
rect 97344 4390 97378 4470
rect 97458 4432 97492 4466
rect 98116 4432 98150 4466
rect 97458 4390 97492 4424
rect 98116 4390 98150 4424
rect 98230 4390 98264 4470
rect 98512 4390 98546 4470
rect 98626 4398 98660 4458
rect 98626 4390 99262 4398
rect 99284 4390 99318 4458
rect 99398 4390 99432 4470
rect 99672 4390 99706 4470
rect 99786 4390 99820 4470
rect 100444 4390 100478 4470
rect 101102 4390 101136 4470
rect 101760 4390 101794 4470
rect 102418 4390 102452 4470
rect 103178 4452 103224 6144
rect 120598 5708 120632 6164
rect 124368 6006 124424 6008
rect 125566 6006 125622 6008
rect 124368 5950 124424 5952
rect 125566 5950 125622 5952
rect 120736 5772 120756 5814
rect 120736 5708 120776 5772
rect 120780 5708 120804 5744
rect 120816 5708 121402 5744
rect 103076 4390 103110 4424
rect 94960 4356 103144 4390
rect 96298 4294 96680 4356
rect 96264 4268 96680 4294
rect 82140 4225 90586 4259
rect 96216 4260 96680 4268
rect 82140 3417 85764 4225
rect 90577 4026 90586 4225
rect 90615 3988 90624 4197
rect 95520 4018 95538 4240
rect 95548 4018 95566 4212
rect 96216 4182 96298 4260
rect 97344 4074 97378 4356
rect 98230 4074 98264 4356
rect 98512 4074 98546 4356
rect 98626 4260 99262 4356
rect 99284 4260 99318 4356
rect 98626 4074 99342 4260
rect 99398 4074 99432 4356
rect 97308 4062 98300 4074
rect 95046 3924 95588 3952
rect 95006 3884 95554 3918
rect 94972 3822 94992 3856
rect 88886 3628 90238 3644
rect 95006 3602 95040 3884
rect 95368 3804 95379 3815
rect 95070 3760 95142 3798
rect 95192 3770 95379 3804
rect 95380 3760 95452 3798
rect 95108 3726 95142 3760
rect 95368 3716 95379 3727
rect 95418 3726 95452 3760
rect 95192 3682 95379 3716
rect 95520 3602 95554 3884
rect 95604 3870 95800 3972
rect 95602 3630 95800 3870
rect 95006 3568 95554 3602
rect 95604 3510 95800 3630
rect 95998 3510 96242 3972
rect 80746 1985 80792 1997
rect 82034 1957 82040 2046
rect 82062 2000 82096 2046
rect 82062 1997 82102 2000
rect 82062 1985 82108 1997
rect 82140 1934 83568 3417
rect 83594 1960 83652 1988
rect 84252 1960 84310 1988
rect 84910 1960 84968 1988
rect 85568 1960 85626 1988
rect 83606 1956 83640 1960
rect 84264 1956 84298 1960
rect 84922 1956 84956 1960
rect 85580 1956 85614 1960
rect 85694 1934 85728 3417
rect 87117 2713 87262 2812
rect 97344 2800 97378 4062
rect 98230 2800 98264 4062
rect 98476 4056 99468 4074
rect 98512 4018 98546 4056
rect 98626 4026 99342 4056
rect 98626 4018 98660 4026
rect 99284 4018 99318 4026
rect 99398 4018 99432 4056
rect 98420 4000 99524 4018
rect 98512 2792 98546 4000
rect 98626 2882 98660 4000
rect 99284 2882 99318 4000
rect 99398 2792 99432 4000
rect 99672 2788 99706 4356
rect 100476 2866 100484 3958
rect 101196 3218 101198 3958
rect 101196 2834 101222 2890
rect 101152 2810 101198 2834
rect 103190 2788 103224 4452
rect 120000 5674 121402 5708
rect 120000 4164 120034 5674
rect 120449 5594 120561 5606
rect 120598 5594 120632 5674
rect 120195 5591 120561 5594
rect 120055 5572 120136 5579
rect 120055 5548 120170 5572
rect 120195 5560 120546 5591
rect 120564 5560 120632 5594
rect 120449 5548 120546 5560
rect 120055 5544 120136 5548
rect 120055 5532 120142 5544
rect 120096 5520 120142 5532
rect 120496 5524 120530 5548
rect 120102 5501 120136 5520
rect 120490 5504 120536 5524
rect 120055 5500 120136 5501
rect 120055 5488 120183 5500
rect 120437 5488 120448 5499
rect 120055 5454 120448 5488
rect 120462 5476 120564 5496
rect 120086 5442 120183 5454
rect 120102 4964 120136 5442
rect 120449 5426 120530 5473
rect 120496 4949 120530 5426
rect 120449 4948 120530 4949
rect 120449 4936 120546 4948
rect 120598 4936 120632 5560
rect 120736 5206 120776 5674
rect 120780 5206 120804 5674
rect 120816 5304 121402 5674
rect 124368 5348 124424 5350
rect 125566 5348 125622 5350
rect 120816 5280 121844 5304
rect 124368 5292 124424 5294
rect 125566 5292 125622 5294
rect 121212 5266 121844 5280
rect 121246 5206 121264 5262
rect 121272 5206 121784 5244
rect 120736 5152 120756 5206
rect 121246 5100 121264 5152
rect 121274 5128 121292 5152
rect 120055 4914 120136 4921
rect 120055 4896 120170 4914
rect 120195 4902 120546 4936
rect 120564 4902 120632 4936
rect 120055 4886 120136 4896
rect 120055 4874 120142 4886
rect 120096 4868 120142 4874
rect 120188 4872 120364 4894
rect 120449 4890 120546 4902
rect 120496 4870 120530 4890
rect 120102 4843 120136 4868
rect 120055 4842 120136 4843
rect 120138 4842 120142 4868
rect 120166 4844 120392 4866
rect 120490 4846 120536 4870
rect 120166 4842 120170 4844
rect 120055 4830 120183 4842
rect 120437 4830 120448 4841
rect 120055 4796 120448 4830
rect 120462 4818 120564 4842
rect 120086 4784 120183 4796
rect 120102 4306 120136 4784
rect 120449 4768 120530 4815
rect 120496 4291 120530 4768
rect 120449 4290 120530 4291
rect 120449 4278 120546 4290
rect 120598 4278 120632 4902
rect 120195 4247 120546 4278
rect 120195 4244 120561 4247
rect 120564 4244 120632 4278
rect 120449 4232 120561 4244
rect 120496 4200 120530 4202
rect 120496 4184 120530 4198
rect 120598 4164 120632 4244
rect 120816 4164 121402 5082
rect 120000 4130 121402 4164
rect 124368 4132 124424 4134
rect 125566 4132 125622 4134
rect 120598 4120 120632 4130
rect 120816 4094 121402 4130
rect 123412 4080 124336 4106
rect 124368 4076 124424 4078
rect 125566 4076 125622 4078
rect 123446 4046 124336 4072
rect 119944 3648 120592 3658
rect 120808 3604 122828 3640
rect 120094 3602 122828 3604
rect 120054 3580 122828 3602
rect 119998 3570 122828 3580
rect 119998 3542 120032 3570
rect 120054 3542 120447 3568
rect 119964 3536 120447 3542
rect 119964 3534 120066 3536
rect 87371 2350 87516 2713
rect 94844 2712 95764 2736
rect 96034 2712 96084 2736
rect 96109 2713 96954 2731
rect 97344 2713 98264 2731
rect 98512 2730 98546 2731
rect 99398 2730 99432 2731
rect 98512 2713 99432 2730
rect 99672 2726 99706 2731
rect 103190 2726 103224 2736
rect 99672 2713 99768 2726
rect 96109 2712 96990 2713
rect 94810 2678 95798 2682
rect 96000 2678 96030 2682
rect 96127 2676 96990 2712
rect 97308 2668 98300 2713
rect 98476 2660 99468 2713
rect 99636 2692 99768 2713
rect 101180 2692 103224 2726
rect 99636 2656 99751 2692
rect 101234 2658 103258 2682
rect 89550 2586 89628 2609
rect 89545 2558 89628 2581
rect 87371 1934 90792 1970
rect 82140 1922 90792 1934
rect 93216 1932 93220 2536
rect 93244 2496 93290 2508
rect 93244 2484 93284 2496
rect 94784 2492 96066 2528
rect 96163 2492 96197 2581
rect 93244 1932 93276 2484
rect 94784 2458 97056 2492
rect 82140 1911 83594 1922
rect 83652 1911 84252 1922
rect 84310 1911 84910 1922
rect 84968 1911 90792 1922
rect 82140 1900 83605 1911
rect 83641 1900 84263 1911
rect 84299 1900 84921 1911
rect 84957 1900 90792 1911
rect 82140 1884 83568 1900
rect 85694 1890 85728 1900
rect 85276 1888 85764 1890
rect 82140 1882 83590 1884
rect 83656 1882 84248 1884
rect 85694 1882 85728 1888
rect 82140 1856 83568 1882
rect 82140 1854 83618 1856
rect 83628 1854 84276 1856
rect 82140 1820 83568 1854
rect 85276 1832 85820 1862
rect 85694 1820 85728 1832
rect 82140 1798 85728 1820
rect 82140 1786 86204 1798
rect 82140 1774 83752 1786
rect 84162 1780 86204 1786
rect 84162 1774 84280 1780
rect 82140 1766 84280 1774
rect 73566 1272 74602 1280
rect 74522 1192 74602 1200
rect 76912 600 76920 1742
rect 82408 0 82442 1766
rect 82878 1748 84280 1766
rect 83752 1742 84162 1746
rect 82850 1720 84308 1742
rect 82884 532 84286 546
rect 87371 -1654 90792 1900
rect 89062 -1764 89274 -1654
rect 92592 -5480 92626 0
rect 93216 -1612 93220 828
rect 93244 0 93276 828
rect 93376 772 93398 1988
rect 94566 1518 94600 1538
rect 94642 1518 94662 1914
rect 94566 1490 94704 1518
rect 94542 1262 94742 1490
rect 93244 -1668 93284 0
rect 93250 -5480 93284 -1668
rect 93908 -5480 93942 0
rect 94566 -5480 94600 1262
rect 94642 1222 94662 1244
rect 94784 1160 96066 2458
rect 96163 1160 96197 2458
rect 96277 2452 96311 2458
rect 96222 2356 96231 2390
rect 96265 2356 96269 2437
rect 96271 2406 96311 2452
rect 96271 2396 96323 2406
rect 96277 2390 96323 2396
rect 96880 2390 96927 2437
rect 96277 2356 96927 2390
rect 96277 2309 96323 2356
rect 96214 2026 96240 2298
rect 96277 2297 96311 2309
rect 96897 2297 96923 2308
rect 96935 2297 96969 2458
rect 96250 1321 96311 2297
rect 96908 1666 96969 2297
rect 96908 1512 96988 1666
rect 96894 1324 96988 1512
rect 96908 1321 96988 1324
rect 96277 1309 96311 1321
rect 96918 1309 96988 1321
rect 96222 1228 96231 1262
rect 96265 1228 96269 1309
rect 96277 1262 96323 1309
rect 96880 1262 96988 1309
rect 96277 1228 96988 1262
rect 96277 1222 96323 1228
rect 96271 1212 96323 1222
rect 96271 1166 96311 1212
rect 96918 1210 96988 1228
rect 96277 1160 96311 1166
rect 96935 1160 96969 1210
rect 97022 1160 97056 2458
rect 94784 1126 97056 1160
rect 97398 2452 99613 2486
rect 97398 1154 97432 2452
rect 97593 2400 97640 2431
rect 97581 2384 97640 2400
rect 98142 2384 98189 2431
rect 98251 2400 98298 2431
rect 98239 2384 98298 2400
rect 98800 2384 98847 2431
rect 98909 2400 98956 2431
rect 98897 2384 98956 2400
rect 99458 2384 99505 2431
rect 97574 2350 98189 2384
rect 98232 2350 98847 2384
rect 98890 2359 99505 2384
rect 98878 2350 99505 2359
rect 97478 2296 97500 2331
rect 97581 2303 97639 2350
rect 97506 2302 97528 2303
rect 97501 2291 97546 2302
rect 97512 2000 97546 2291
rect 97559 2000 97580 2296
rect 97478 1275 97500 2000
rect 97506 1315 97546 2000
rect 97587 1972 97627 2303
rect 98136 2302 98162 2331
rect 98239 2303 98297 2350
rect 98878 2344 98956 2350
rect 98897 2303 98956 2344
rect 98164 2302 98210 2303
rect 98136 2291 98210 2302
rect 98136 2250 98162 2291
rect 97506 1303 97528 1315
rect 97593 1303 97627 1972
rect 98108 1518 98162 2250
rect 98164 2194 98210 2291
rect 98164 1882 98204 2194
rect 98251 1882 98285 2303
rect 98847 2302 98868 2303
rect 98903 2302 98956 2303
rect 98817 2291 98900 2302
rect 98828 2020 98900 2291
rect 98828 1882 98868 2020
rect 98903 1882 98943 2302
rect 99475 2291 99520 2302
rect 99486 1882 99520 2291
rect 99561 2164 99582 2359
rect 98164 1518 98215 1882
rect 98170 1315 98215 1518
rect 98230 1310 98238 1526
rect 98108 1303 98162 1308
rect 98164 1303 98190 1308
rect 98251 1303 98296 1882
rect 98828 1315 98873 1882
rect 98847 1303 98868 1315
rect 98903 1303 98954 1882
rect 99486 1315 99531 1882
rect 97581 1256 97640 1303
rect 98108 1256 99505 1303
rect 97574 1222 98189 1256
rect 98232 1222 98847 1256
rect 98878 1247 99505 1256
rect 97581 1206 97639 1222
rect 98146 1194 98162 1222
rect 98239 1206 98297 1222
rect 98878 1216 98888 1247
rect 98890 1222 99505 1247
rect 98897 1206 98955 1222
rect 99567 1154 99572 1188
rect 99600 1154 99613 2452
rect 94784 1090 96066 1126
rect 95806 284 96066 320
rect 96163 284 96197 1126
rect 97398 1120 99613 1154
rect 99681 780 99715 2581
rect 99354 746 100800 780
rect 95806 250 98736 284
rect 95806 -548 96066 250
rect 96163 -548 96197 250
rect 96277 213 96324 229
rect 96265 182 96324 213
rect 96586 182 96633 229
rect 96935 198 96982 229
rect 96923 182 96982 198
rect 97244 182 97291 229
rect 97593 198 97640 229
rect 97581 182 97640 198
rect 97902 182 97949 229
rect 98251 198 98298 229
rect 98239 182 98298 198
rect 98560 182 98607 229
rect 96265 148 96633 182
rect 96676 148 97291 182
rect 97334 148 97949 182
rect 97992 148 98607 182
rect 96265 101 96323 148
rect 96923 101 96981 148
rect 97581 101 97639 148
rect 98239 101 98297 148
rect 96277 -399 96311 101
rect 96603 89 96648 100
rect 96614 -387 96648 89
rect 96935 -399 96969 101
rect 97261 89 97306 100
rect 97272 -387 97306 89
rect 97593 -399 97627 101
rect 97919 89 97964 100
rect 97930 -387 97964 89
rect 98251 -399 98285 101
rect 98577 89 98622 100
rect 98588 -387 98622 89
rect 96265 -446 96324 -399
rect 96586 -446 96633 -399
rect 96923 -446 96982 -399
rect 97244 -446 97291 -399
rect 97581 -446 97640 -399
rect 97902 -446 97949 -399
rect 98239 -446 98298 -399
rect 98560 -446 98607 -399
rect 96265 -480 96633 -446
rect 96676 -480 97291 -446
rect 97334 -480 97949 -446
rect 97992 -480 98607 -446
rect 96265 -496 96323 -480
rect 96923 -496 96981 -480
rect 97581 -496 97639 -480
rect 98239 -496 98297 -480
rect 96265 -511 96280 -496
rect 98702 -548 98736 250
rect 95806 -582 98736 -548
rect 99354 -552 99388 746
rect 99483 678 99613 725
rect 99530 644 99613 678
rect 99555 597 99613 644
rect 99457 585 99513 596
rect 99468 564 99513 585
rect 99567 564 99612 597
rect 99468 -391 99502 564
rect 99567 -403 99601 564
rect 99555 -450 99613 -403
rect 99530 -484 99613 -450
rect 99555 -500 99613 -484
rect 99598 -515 99613 -500
rect 99681 -552 99715 746
rect 101240 466 101286 482
rect 99354 -558 100800 -552
rect 95806 -618 96066 -582
rect 96163 -5593 96197 -582
rect 99354 -586 100968 -558
rect 96450 -4358 96840 -4324
rect 96450 -4856 96484 -4358
rect 96664 -4426 96711 -4379
rect 96626 -4460 96711 -4426
rect 96553 -4519 96598 -4508
rect 96681 -4519 96726 -4508
rect 96564 -4695 96598 -4519
rect 96692 -4695 96726 -4519
rect 96664 -4754 96711 -4707
rect 96626 -4788 96711 -4754
rect 96806 -4856 96840 -4358
rect 96450 -4890 96840 -4856
rect 96432 -5560 96854 -4940
rect 99681 -5593 99715 -586
rect 100102 -622 100968 -586
rect 101404 -620 103054 818
rect 103398 810 103418 1914
rect 103322 -1048 103356 0
rect 103508 -622 104822 2718
rect 119998 1480 120032 3534
rect 120153 3500 120436 3524
rect 120490 3506 120524 3524
rect 120443 3496 120555 3502
rect 120181 3487 120555 3496
rect 120592 3490 120626 3570
rect 120053 3428 120134 3475
rect 120181 3472 120540 3487
rect 120193 3456 120540 3472
rect 120558 3456 120626 3490
rect 120443 3444 120540 3456
rect 120100 2923 120134 3428
rect 120490 2938 120524 3444
rect 120053 2922 120134 2923
rect 120053 2910 120181 2922
rect 120431 2910 120442 2921
rect 120053 2876 120442 2910
rect 120084 2870 120400 2876
rect 120084 2864 120181 2870
rect 120100 2860 120134 2864
rect 120186 2842 120372 2860
rect 120443 2848 120524 2895
rect 120490 2845 120524 2848
rect 120443 2844 120524 2845
rect 120443 2832 120540 2844
rect 120592 2832 120626 3456
rect 120053 2770 120134 2817
rect 120193 2798 120540 2832
rect 120558 2798 120626 2832
rect 120443 2786 120540 2798
rect 120100 2265 120134 2770
rect 120490 2280 120524 2786
rect 120053 2264 120134 2265
rect 120053 2252 120181 2264
rect 120431 2252 120442 2263
rect 120053 2218 120442 2252
rect 120084 2206 120181 2218
rect 120100 2202 120140 2206
rect 120132 2190 120140 2202
rect 120160 2180 120168 2206
rect 120443 2190 120524 2237
rect 120490 2187 120524 2190
rect 120443 2186 120524 2187
rect 120443 2174 120540 2186
rect 120592 2174 120626 2798
rect 120808 3464 122828 3570
rect 120808 3450 122998 3464
rect 120808 3436 122828 3450
rect 120808 3422 122970 3436
rect 120808 2780 122828 3422
rect 120053 2112 120134 2159
rect 120193 2140 120540 2174
rect 120558 2140 120626 2174
rect 120443 2128 120540 2140
rect 120100 1607 120134 2112
rect 120490 1622 120524 2128
rect 120053 1606 120134 1607
rect 120053 1594 120181 1606
rect 120431 1594 120442 1605
rect 120053 1560 120442 1594
rect 120069 1554 120420 1560
rect 120069 1550 120181 1554
rect 120069 1548 120392 1550
rect 120170 1526 120392 1548
rect 120066 1480 120168 1488
rect 120193 1482 120564 1514
rect 120592 1480 120626 2140
rect 120800 2174 122820 2604
rect 120800 2140 124169 2174
rect 120800 1612 122820 2140
rect 119356 1446 120626 1480
rect 119998 148 120032 1446
rect 120796 16 124400 1444
rect 120934 -10 120968 16
rect 121030 -6 121358 16
rect 103454 -792 103476 -788
rect 103426 -820 103448 -816
rect 103426 -1046 103450 -820
rect 103426 -1048 103448 -1046
rect 103454 -1048 103478 -792
rect 103132 -1060 103478 -1048
rect 103322 -5480 103356 -1060
rect 103454 -1074 103478 -1060
rect 103454 -1078 103476 -1074
<< metal1 >>
rect 115246 37884 116090 37976
rect 115246 36592 115344 37884
rect 115990 36592 116090 37884
rect 115246 7558 116090 36592
rect 116630 19234 118352 19318
rect 116630 18934 117242 19234
rect 117738 18934 118352 19234
rect 116630 18826 118352 18934
rect 115246 7544 117490 7558
rect 115246 6510 117510 7544
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
rect 0 -2400 200 -2200
rect 0 -2800 200 -2600
rect 0 -3200 200 -3000
rect 0 -3600 200 -3400
rect 0 -4000 200 -3800
rect 0 -4400 200 -4200
rect 0 -4800 200 -4600
rect 0 -5200 200 -5000
rect 0 -5600 200 -5400
rect 0 -6000 200 -5800
rect 116710 -6192 117510 6510
rect 124560 -6762 125568 -2142
rect 124560 -7340 124626 -6762
rect 125510 -7340 125568 -6762
rect 124560 -7412 125568 -7340
<< via1 >>
rect 115344 36592 115990 37884
rect 117242 18934 117738 19234
rect 124626 -7340 125510 -6762
<< metal2 >>
rect 38638 51484 131148 52740
rect 38638 46984 74732 51484
rect 85778 46984 131148 51484
rect 38638 40548 131148 46984
rect 38568 37884 131148 40548
rect 38568 37356 115344 37884
rect 34294 36152 35444 36428
rect 34294 33872 34506 36152
rect 35272 33872 35444 36152
rect 31892 23726 33640 23732
rect 9654 23718 33640 23726
rect 9654 23350 33664 23718
rect 9654 21480 10088 23350
rect 11798 21480 33664 23350
rect 9654 20970 33664 21480
rect 31892 1200 33640 20970
rect 34294 14406 35444 33872
rect 38568 32790 77824 37356
rect 106022 36592 115344 37356
rect 115990 37356 131148 37884
rect 115990 36592 118004 37356
rect 106022 36356 118004 36592
rect 117070 19234 117886 19328
rect 117070 18934 117242 19234
rect 117738 18934 117886 19234
rect 117070 18836 117886 18934
rect 34294 14002 38616 14406
rect 34294 12490 37552 14002
rect 38318 12490 38616 14002
rect 34294 12212 38616 12490
rect 31892 1054 36900 1200
rect 31892 278 36224 1054
rect 36752 278 36900 1054
rect 31892 142 36900 278
rect 41102 -5498 74748 2998
rect 124096 -5026 124576 -4942
rect 124096 -5452 124144 -5026
rect 124488 -5452 124576 -5026
rect 40590 -6576 115178 -5498
rect 124096 -5518 124576 -5452
rect 40590 -6758 125590 -6576
rect 126230 -6758 130010 18604
rect 40590 -6762 130010 -6758
rect 40590 -7340 124626 -6762
rect 125510 -7340 130010 -6762
rect 40590 -12342 130010 -7340
rect 40590 -14092 77484 -12342
rect 40704 -16842 77484 -14092
rect 88530 -16842 130010 -12342
rect 40704 -18276 130010 -16842
rect 40704 -18560 129728 -18276
<< via2 >>
rect 74732 46984 85778 51484
rect 34506 33872 35272 36152
rect 10088 21480 11798 23350
rect 118568 33404 119192 34818
rect 118564 24274 119418 25920
rect 132062 20278 132868 35914
rect 117242 18934 117738 19234
rect 37552 12490 38318 14002
rect 36224 278 36752 1054
rect 124144 -5452 124488 -5026
rect 77484 -16842 88530 -12342
<< metal3 >>
rect 73654 51484 87112 52368
rect 73654 46984 74732 51484
rect 85778 46984 87112 51484
rect 73654 46042 87112 46984
rect 73958 43414 76222 43718
rect 73958 41284 74396 43414
rect 75884 41284 76222 43414
rect 34378 36152 35464 36364
rect 34378 33872 34506 36152
rect 35272 33872 35464 36152
rect 34378 33596 35464 33872
rect 34328 31840 35374 32224
rect 34328 29770 34564 31840
rect 35204 29770 35374 31840
rect 9564 27608 33764 28046
rect 9564 25666 9960 27608
rect 11782 25666 33764 27608
rect 9564 25212 33764 25666
rect 9854 23350 11996 23570
rect 9854 21480 10088 23350
rect 11798 21480 11996 23350
rect 9854 21184 11996 21480
rect 31854 -366 33700 25212
rect 34328 24368 35374 29770
rect 73958 26428 76222 41284
rect 131792 35914 133096 36374
rect 118380 34818 119406 35048
rect 118380 33404 118568 34818
rect 119192 33404 119406 34818
rect 118380 33242 119406 33404
rect 34328 23580 38810 24368
rect 70006 23786 76222 26428
rect 118440 25920 119530 26070
rect 118440 24274 118564 25920
rect 119418 24274 119530 25920
rect 118440 24092 119530 24274
rect 70006 22762 76138 23786
rect 70006 21552 74518 22762
rect 75942 21552 76138 22762
rect 70006 21386 76138 21552
rect 131792 20278 132062 35914
rect 132868 20278 133096 35914
rect 131792 19972 133096 20278
rect 117070 19234 117886 19328
rect 117070 18934 117242 19234
rect 117738 18934 117886 19234
rect 117070 18836 117886 18934
rect 37382 14002 38660 14384
rect 37382 12490 37552 14002
rect 38318 12490 38660 14002
rect 37382 12190 38660 12490
rect 113712 6498 115052 6502
rect 74602 1200 75588 6492
rect 113712 5590 118242 6498
rect 36100 1054 75588 1200
rect 36100 278 36224 1054
rect 36752 278 75588 1054
rect 36100 154 75588 278
rect 74602 118 75588 154
rect 31854 -398 94850 -366
rect 113712 -398 115052 5590
rect 31854 -1610 115052 -398
rect 31854 -1612 94850 -1610
rect 113712 -1626 115052 -1610
rect 121048 -1858 121444 -1614
rect 124086 -4720 124652 -4566
rect 124086 -5026 124148 -4720
rect 124086 -5452 124144 -5026
rect 124086 -5702 124148 -5452
rect 124542 -5702 124652 -4720
rect 124086 -5854 124652 -5702
rect 75650 -12342 89972 -11570
rect 75650 -16842 77484 -12342
rect 88530 -16842 89972 -12342
rect 75650 -17872 89972 -16842
<< via3 >>
rect 74732 46984 85778 51484
rect 74396 41284 75884 43414
rect 34506 33872 35272 36152
rect 34564 29770 35204 31840
rect 9960 25666 11782 27608
rect 10088 21480 11798 23350
rect 37940 27438 38382 29510
rect 78850 33204 79772 34172
rect 118568 33404 119192 34818
rect 78878 30960 79800 31928
rect 78920 24196 79842 25164
rect 118564 24274 119418 25920
rect 74518 21552 75942 22762
rect 78906 22036 79828 23004
rect 78934 19876 79856 20844
rect 132062 20278 132868 35914
rect 117242 18934 117738 19234
rect 37774 6508 38902 7930
rect 78640 2238 79568 3180
rect 124148 -5026 124542 -4720
rect 124148 -5452 124488 -5026
rect 124488 -5452 124542 -5026
rect 124148 -5702 124542 -5452
rect 77484 -16842 88530 -12342
<< metal4 >>
rect 73654 51484 87112 52368
rect 73654 46984 74732 51484
rect 85778 46984 87112 51484
rect 73654 46042 87112 46984
rect 31626 44780 33968 45110
rect 31626 42372 31940 44780
rect 33600 42372 33968 44780
rect 9792 27608 11934 27828
rect 9792 25666 9960 27608
rect 11782 25666 11934 27608
rect 9792 25442 11934 25666
rect 9854 23350 11996 23570
rect 9854 21480 10088 23350
rect 11798 21480 11996 23350
rect 9854 21184 11996 21480
rect 9474 18854 31096 19376
rect 9474 17130 9896 18854
rect 11568 17130 31096 18854
rect 9474 16546 31096 17130
rect 29446 3306 31096 16546
rect 31626 8892 33968 42372
rect 74126 43414 76222 43718
rect 74126 41284 74396 43414
rect 75884 41284 76222 43414
rect 74126 40880 76222 41284
rect 35804 40318 38372 40424
rect 35804 38110 36186 40318
rect 37862 38110 38372 40318
rect 34378 36152 35464 36364
rect 34378 33872 34506 36152
rect 35272 33872 35464 36152
rect 34378 33596 35464 33872
rect 34350 31840 35416 32202
rect 34350 29770 34564 31840
rect 35204 29770 35416 31840
rect 34350 29556 35416 29770
rect 35804 29984 38372 38110
rect 127328 35914 133002 36562
rect 118380 34818 119406 35048
rect 78638 34172 80048 34440
rect 78638 33204 78850 34172
rect 79772 33204 80048 34172
rect 118380 33404 118568 34818
rect 119192 33404 119406 34818
rect 118380 33242 119406 33404
rect 78638 32942 80048 33204
rect 78660 31928 80070 32170
rect 78660 30960 78878 31928
rect 79800 30960 80070 31928
rect 78660 30672 80070 30960
rect 35804 29510 38498 29984
rect 35804 27438 37940 29510
rect 38382 27438 38498 29510
rect 35804 26930 38498 27438
rect 113388 25920 119628 26604
rect 78682 25164 80092 25450
rect 78682 24196 78920 25164
rect 79842 24196 80092 25164
rect 78682 23952 80092 24196
rect 113388 24274 118564 25920
rect 119418 24274 119628 25920
rect 113388 23456 119628 24274
rect 78690 23004 80100 23252
rect 74290 22762 76138 22942
rect 74290 21552 74518 22762
rect 75942 21552 76138 22762
rect 78690 22036 78906 23004
rect 79828 22036 80100 23004
rect 78690 21754 80100 22036
rect 74290 19474 76138 21552
rect 78696 20844 80106 21134
rect 78696 19876 78934 20844
rect 79856 19876 80106 20844
rect 78696 19636 80106 19876
rect 127328 20278 132062 35914
rect 132868 20278 133002 35914
rect 117070 19234 117886 19328
rect 117070 18934 117242 19234
rect 117738 18934 117886 19234
rect 117070 18836 117886 18934
rect 127328 11774 133002 20278
rect 31626 7930 39404 8892
rect 31626 6508 37774 7930
rect 38902 6508 39404 7930
rect 119950 7034 133002 11774
rect 119950 6730 132996 7034
rect 31626 5588 39404 6508
rect 29446 3180 79670 3306
rect 29446 2238 78640 3180
rect 79568 2238 79670 3180
rect 29446 2148 79670 2238
rect 124116 -3612 124996 -3456
rect 124116 -4720 124202 -3612
rect 124116 -5702 124148 -4720
rect 124116 -6046 124202 -5702
rect 124846 -6046 124996 -3612
rect 124116 -6172 124996 -6046
rect 75650 -12342 89972 -11570
rect 75650 -16842 77484 -12342
rect 88530 -16842 89972 -12342
rect 75650 -17872 89972 -16842
<< via4 >>
rect 74732 46984 85778 51484
rect 31940 42372 33600 44780
rect 9960 25666 11782 27608
rect 10088 21480 11798 23350
rect 9896 17130 11568 18854
rect 74396 41284 75884 43414
rect 36186 38110 37862 40318
rect 34506 33872 35272 36152
rect 34564 29770 35204 31840
rect 78850 33204 79772 34172
rect 118568 33404 119192 34818
rect 78878 30960 79800 31928
rect 78920 24196 79842 25164
rect 78906 22036 79828 23004
rect 78934 19876 79856 20844
rect 117242 18934 117738 19234
rect 124202 -4720 124846 -3612
rect 124202 -5702 124542 -4720
rect 124542 -5702 124846 -4720
rect 124202 -6046 124846 -5702
rect 77484 -16842 88530 -12342
<< metal5 >>
rect 35738 51484 131268 52674
rect 35738 46984 74732 51484
rect 85778 46984 131268 51484
rect 35738 45616 131268 46984
rect 9536 44984 12182 44994
rect 9536 44976 13158 44984
rect 31480 44976 33926 44984
rect 9536 44780 34012 44976
rect 9536 42372 31940 44780
rect 33600 42372 34012 44780
rect 9536 42222 34012 42372
rect 9540 42182 34012 42222
rect 74060 43414 119596 43718
rect 74060 41284 74396 43414
rect 75884 41284 119596 43414
rect 74060 40914 119596 41284
rect 9568 40558 13158 40572
rect 31480 40558 38308 40572
rect 9568 40318 38308 40558
rect 9568 38110 36186 40318
rect 37862 38110 38308 40318
rect 9568 37814 38308 38110
rect 9600 37788 12246 37814
rect 9564 36364 12210 36380
rect 9564 36338 13158 36364
rect 31480 36338 35422 36364
rect 9564 36152 35422 36338
rect 9564 33872 34506 36152
rect 35272 33872 35422 36152
rect 115914 34818 119596 40914
rect 9564 33608 35422 33872
rect 78518 34418 87750 34528
rect 78518 34172 87776 34418
rect 78518 33204 78850 34172
rect 79772 33204 87776 34172
rect 78518 32832 87776 33204
rect 9564 32224 12210 32228
rect 9564 32216 13158 32224
rect 31480 32216 35396 32224
rect 9564 31840 35396 32216
rect 9564 29770 34564 31840
rect 35204 29770 35396 31840
rect 78540 32176 85238 32256
rect 78540 31928 85262 32176
rect 78540 30960 78878 31928
rect 79800 30960 85262 31928
rect 78540 30612 85262 30960
rect 9564 29456 35396 29770
rect 9564 27608 12210 27984
rect 9564 25666 9960 27608
rect 11782 25666 12210 27608
rect 9564 25212 12210 25666
rect 13446 25642 16160 25798
rect 13446 25164 80184 25642
rect 13446 24196 78920 25164
rect 79842 24196 80184 25164
rect 13446 23814 80184 24196
rect 9654 23350 12300 23742
rect 9654 21480 10088 23350
rect 11798 21480 12300 23350
rect 9654 20970 12300 21480
rect 9474 18854 12120 19318
rect 9474 17130 9896 18854
rect 11568 17130 12120 18854
rect 9474 16546 12120 17130
rect 13446 14938 16160 23814
rect 80900 23336 82746 23338
rect 78584 23004 82788 23336
rect 78584 22036 78906 23004
rect 79828 22036 82788 23004
rect 78584 21670 82788 22036
rect 17816 21178 19798 21266
rect 17784 20844 80214 21178
rect 17784 19876 78934 20844
rect 79856 19876 80214 20844
rect 17784 19532 80214 19876
rect 9474 12124 16162 14938
rect 17816 10500 19798 19532
rect 9382 7700 19850 10500
rect 9382 6010 12028 6050
rect 80900 6010 82746 21670
rect 9382 3820 82746 6010
rect 9382 3284 82740 3820
rect 9382 3278 82632 3284
rect 83112 1632 85262 30612
rect 9292 -1124 85262 1632
rect 9292 -1146 84814 -1124
rect 86016 -2672 87776 32832
rect 115914 33404 118568 34818
rect 119192 33404 119596 34818
rect 115914 32400 119596 33404
rect 116636 19234 118340 19322
rect 116636 18934 117242 19234
rect 117738 18934 118340 19234
rect 9112 -5478 87778 -2672
rect 116636 -6888 118340 18934
rect 124100 -3442 125862 -3428
rect 133226 -3442 135962 -3422
rect 124100 -3612 135962 -3442
rect 124100 -6046 124202 -3612
rect 124846 -6046 135962 -3612
rect 124100 -6194 135962 -6046
rect 124100 -6212 135950 -6194
rect 124946 -6222 135950 -6212
rect 9022 -9722 120478 -6888
rect 116636 -9730 118340 -9722
rect 34564 -12342 130094 -11238
rect 34564 -16842 77484 -12342
rect 88530 -16842 130094 -12342
rect 34564 -18296 130094 -16842
use buffer  buffer_0
timestamp 1695698273
transform 1 0 70830 0 1 -1726
box -6068 -1844 19288 11182
use diffamp  diffamp_0
timestamp 1695698273
transform 1 0 -27400 0 1 32314
box 0 -31714 61184 4684
use integrator  integrator_0
timestamp 1695698273
transform 1 0 19202 0 1 11168
box 0 -10568 125722 37774
use mux2_1  mux2_1_0
timestamp 1695698273
transform 1 0 85918 0 1 -7822
box -476 -1200 20872 33492
use diffamp  x1
timestamp 1695698273
transform 1 0 10044 0 1 31138
box 0 -31714 61184 4684
use integrator  x2
timestamp 1695698273
transform 1 0 57968 0 1 4200
box 0 -10568 125722 37774
use mux2_1  x3
timestamp 1695698273
transform 1 0 112232 0 1 6854
box -476 -1200 20872 33492
use buffer  x7
timestamp 1695698273
transform 0 -1 127892 -1 0 12754
box -6068 -1844 19288 11182
<< labels >>
rlabel metal5 34564 -18296 130094 -11238 1 GROUND
port 2 nsew
rlabel metal5 35738 45616 131268 52674 1 VDD
port 1 nsew
rlabel metal5 9536 42222 12182 44994 1 AIn0
port 3 nsew
rlabel metal5 9600 37788 12246 40560 1 AIn1
port 4 nsew
rlabel metal5 9564 33608 12210 36380 1 AIn2
port 5 nsew
rlabel metal5 9564 29456 12210 32228 1 AIn3
port 6 nsew
rlabel metal5 9564 25212 12210 27984 1 AIn4
port 7 nsew
rlabel metal5 9654 20970 12300 23742 1 AIn5
port 8 nsew
rlabel metal5 9474 16546 12120 19318 1 REG0
port 9 nsew
rlabel metal5 9474 12124 12120 14896 1 REG1
port 10 nsew
rlabel metal5 9382 7700 12028 10472 1 REG2
port 11 nsew
rlabel metal5 9382 3278 12028 6050 1 REG3
port 12 nsew
rlabel metal5 9292 -1146 11938 1626 1 REG4
port 13 nsew
rlabel metal5 9112 -5478 11758 -2706 1 REG5
port 14 nsew
rlabel metal5 9022 -9722 11668 -6950 1 REG6
port 15 nsew
rlabel metal5 133316 -6194 135962 -3422 1 AOut
port 16 nsew
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 GROUND
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 AIn0
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 AOut
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 AIn1
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 AIn2
flabel metal1 0 -2400 200 -2200 0 FreeSans 256 0 0 0 AIn3
flabel metal1 0 -2800 200 -2600 0 FreeSans 256 0 0 0 AIn4
flabel metal1 0 -3200 200 -3000 0 FreeSans 256 0 0 0 AIn5
flabel metal1 0 -3600 200 -3400 0 FreeSans 256 0 0 0 REG0
flabel metal1 0 -4000 200 -3800 0 FreeSans 256 0 0 0 REG1
flabel metal1 0 -4400 200 -4200 0 FreeSans 256 0 0 0 REG2
flabel metal1 0 -4800 200 -4600 0 FreeSans 256 0 0 0 REG3
flabel metal1 0 -5200 200 -5000 0 FreeSans 256 0 0 0 REG4
flabel metal1 0 -5600 200 -5400 0 FreeSans 256 0 0 0 REG5
flabel metal1 0 -6000 200 -5800 0 FreeSans 256 0 0 0 REG6
<< end >>
