magic
tech sky130A
magscale 1 2
timestamp 1695461801
<< error_p >>
rect 52128 43866 52130 43916
rect 52156 43866 52158 43944
rect 51576 43626 52214 43866
rect 57342 43822 57344 43900
rect 57370 43822 57372 43872
rect 57286 43582 57924 43822
rect 52110 43320 52130 43440
rect 52138 43314 52158 43468
rect 57342 43270 57362 43424
rect 57370 43276 57390 43396
rect 74349 43234 74383 46377
rect 77095 43234 77129 46278
rect 77867 43234 77901 46377
rect 79420 43234 79454 46382
rect 82938 43234 82972 43838
rect 185426 4780 185432 4800
rect 185618 4782 185858 5334
rect 185618 4780 185908 4782
rect 185426 4752 185460 4772
rect 185618 4754 185858 4780
rect 185618 4752 185936 4754
rect 185618 4696 185858 4752
rect 120999 -3470 121033 -1704
rect 121075 -3460 121076 -3378
rect 121113 -3436 121114 -3340
rect 121113 -3470 121174 -3436
rect 120960 -3504 121236 -3470
rect 120999 -3572 121033 -3504
rect 121006 -3615 121033 -3572
rect 121101 -3606 121107 -3525
rect 120965 -3857 120994 -3649
rect 120999 -3891 121033 -3615
rect 121113 -3665 121147 -3504
rect 121088 -3841 121147 -3665
rect 121006 -3934 121033 -3891
rect 121094 -3924 121098 -3898
rect 121101 -3934 121107 -3853
rect 120999 -3968 121033 -3934
rect 121113 -3968 121147 -3841
rect 120980 -3988 121080 -3968
rect 120999 -3996 121033 -3988
rect 120974 -4002 121080 -3996
rect 121113 -4002 121174 -3968
rect 121202 -4002 121236 -3504
rect 120960 -4036 121236 -4002
rect 121322 -3504 121712 -3470
rect 121322 -4002 121356 -3504
rect 121536 -3572 121583 -3525
rect 121498 -3606 121583 -3572
rect 121425 -3665 121470 -3654
rect 121553 -3665 121598 -3654
rect 121436 -3841 121470 -3665
rect 121564 -3841 121598 -3665
rect 121536 -3900 121583 -3853
rect 121498 -3934 121583 -3900
rect 121678 -4002 121712 -3504
rect 121322 -4036 121712 -4002
rect 121860 -4014 121870 -3664
rect 121888 -4014 121898 -3636
rect 120994 -4048 121033 -4036
rect 120999 -4086 121033 -4048
rect 120963 -4706 121250 -4086
rect 121304 -4706 121726 -4086
rect 121860 -4488 121870 -4200
rect 121888 -4516 121898 -4200
rect 121135 -4767 121162 -4706
rect 121163 -4739 121190 -4706
rect 25484 -7786 25556 -7778
rect 34680 -7786 34752 -7778
rect 25484 -7788 25552 -7786
rect 34680 -7788 34748 -7786
rect 19680 -8276 19684 -7956
rect 19718 -8276 19722 -7956
rect 34762 -8006 34782 -7827
rect 34762 -8027 34792 -8006
rect 34728 -8366 34786 -8364
rect 34702 -8400 34752 -8398
<< error_s >>
rect 77095 40320 77129 43234
rect 74349 40013 74383 40320
rect 74463 40109 74497 40143
rect 75121 40109 75155 40143
rect 75779 40109 75813 40143
rect 76437 40109 76471 40143
rect 77095 40109 77129 40143
rect 77753 40109 77807 40143
rect 74413 40075 74417 40109
rect 74429 40075 77807 40109
rect 5526 36898 5528 36948
rect 5554 36898 5556 36976
rect 4974 36658 5612 36898
rect 10740 36854 10742 36932
rect 10768 36854 10770 36904
rect 10684 36614 11322 36854
rect 5508 36352 5528 36472
rect 5536 36346 5556 36500
rect 10740 36302 10760 36456
rect 10768 36308 10788 36428
rect -1996 30763 -1962 35702
rect 1440 35684 2922 35796
rect 0 35650 6166 35684
rect 1440 35026 2922 35650
rect 0 34992 6166 35026
rect 1440 34368 2922 34992
rect 4974 34368 5612 34466
rect 5662 34380 6210 34408
rect 5662 34374 6178 34380
rect 5662 34368 5696 34374
rect 0 34340 6170 34368
rect 6176 34353 6178 34374
rect 6199 34369 6210 34380
rect 0 34334 6166 34340
rect 1440 34220 2922 34334
rect 4974 34004 5612 34334
rect 5662 34092 5696 34334
rect 6024 34294 6035 34305
rect 5726 34250 5798 34288
rect 5848 34278 6035 34294
rect 6036 34278 6108 34288
rect 5836 34254 6108 34278
rect 6036 34250 6108 34254
rect 5764 34216 5798 34250
rect 5808 34226 6064 34250
rect 6024 34206 6035 34217
rect 6074 34216 6108 34250
rect 5848 34172 6035 34206
rect 6176 34092 6210 34353
rect 5662 34058 6210 34092
rect 4974 33732 5612 33990
rect 4822 33710 5612 33732
rect 0 33676 5612 33710
rect 4822 33658 5612 33676
rect 4974 33528 5612 33658
rect 5662 33898 6210 33932
rect 5662 33710 5696 33898
rect 5726 33774 5798 33812
rect 5802 33802 5834 33822
rect 6024 33818 6035 33829
rect 5802 33774 5806 33794
rect 5848 33784 6035 33818
rect 6036 33774 6108 33812
rect 5764 33724 5798 33774
rect 6024 33730 6035 33741
rect 5848 33722 6035 33730
rect 6074 33724 6108 33774
rect 5848 33710 6024 33722
rect 6176 33711 6210 33898
rect 6216 33816 6250 34306
rect 6318 33816 6352 35702
rect 6216 33738 6352 33816
rect 5662 33676 6166 33710
rect 6176 33695 6200 33711
rect 6176 33688 6210 33695
rect 5662 33616 5696 33676
rect 6176 33672 6284 33688
rect 6176 33660 6210 33672
rect 6176 33644 6256 33660
rect 6176 33616 6210 33644
rect 5662 33582 6210 33616
rect 6216 33340 6250 33644
rect 6318 33340 6352 33738
rect 6216 33254 6352 33340
rect 6216 33144 6250 33254
rect -1921 33133 6277 33144
rect -1910 33121 6266 33133
rect -1921 33110 6277 33121
rect -1894 33064 -1860 33110
rect -880 33064 -422 33084
rect 6216 33080 6250 33110
rect -880 33052 -382 33064
rect -1810 33006 6166 33052
rect -1810 32996 6177 33006
rect -880 32992 -382 32996
rect -1894 32400 -1860 32990
rect -840 32972 -382 32992
rect -1230 32948 -126 32968
rect -1258 32920 -98 32940
rect 2030 32788 2478 32816
rect 2030 32604 2496 32788
rect 2048 32576 2496 32604
rect 4794 32405 5448 32418
rect 1144 32394 3276 32405
rect 3894 32394 6177 32405
rect 6216 32400 6250 32990
rect -1810 32384 6177 32394
rect -1810 32338 6166 32384
rect 4830 32320 5484 32338
rect -1894 32310 -1860 32314
rect 6216 32310 6250 32314
rect -1941 32246 6297 32280
rect 6318 32168 6352 33254
rect 9944 33772 9978 35658
rect 10086 34330 10634 34364
rect 10046 33772 10080 34262
rect 10086 34048 10120 34330
rect 10600 34324 10634 34330
rect 10126 34296 10634 34324
rect 10130 34290 10154 34296
rect 10566 34290 10634 34296
rect 10448 34250 10459 34261
rect 10150 34206 10222 34244
rect 10272 34234 10459 34250
rect 10460 34234 10532 34244
rect 10260 34210 10532 34234
rect 10460 34206 10532 34210
rect 10188 34172 10222 34206
rect 10232 34182 10488 34206
rect 10448 34162 10459 34173
rect 10498 34172 10532 34206
rect 10272 34128 10459 34162
rect 10600 34048 10634 34290
rect 10086 34014 10634 34048
rect 10684 33960 11322 34422
rect 9944 33694 10080 33772
rect 10086 33854 10634 33888
rect 9944 33296 9978 33694
rect 10086 33644 10120 33854
rect 10448 33774 10459 33785
rect 10150 33730 10222 33768
rect 10272 33740 10459 33774
rect 10462 33768 10494 33778
rect 10460 33730 10532 33768
rect 10188 33706 10222 33730
rect 10498 33706 10532 33730
rect 10188 33696 10260 33706
rect 10261 33686 10459 33697
rect 10498 33696 10570 33706
rect 10272 33678 10459 33686
rect 10272 33666 10448 33678
rect 10600 33666 10634 33854
rect 10012 33628 10120 33644
rect 10130 33632 10634 33666
rect 10086 33616 10120 33628
rect 10040 33600 10120 33616
rect 10046 33296 10080 33600
rect 10086 33572 10120 33600
rect 10600 33572 10634 33632
rect 10086 33538 10634 33572
rect 10684 33688 11322 33946
rect 10684 33666 11474 33688
rect 10684 33632 18106 33666
rect 10684 33614 11474 33632
rect 10684 33484 11322 33614
rect 9944 33210 10080 33296
rect 9944 32222 9978 33210
rect 10046 33100 10080 33210
rect 16658 33100 16714 33122
rect 10019 33089 18217 33100
rect 10030 33077 18206 33089
rect 10019 33066 18217 33077
rect 10046 33036 10080 33066
rect 16718 33020 17176 33040
rect 16682 33008 17176 33020
rect 10130 32962 18106 33008
rect 10130 32952 18117 32962
rect 16682 32948 17176 32952
rect 10046 32356 10080 32946
rect 16682 32928 17136 32948
rect 16658 32904 17526 32924
rect 15646 32890 15702 32896
rect 16658 32876 17554 32896
rect 16658 32848 16714 32876
rect 13818 32744 14266 32772
rect 13800 32560 14266 32744
rect 13800 32532 14248 32560
rect 10848 32361 11502 32374
rect 10119 32350 18117 32361
rect 18156 32356 18190 32946
rect 10130 32340 18117 32350
rect 10130 32294 18106 32340
rect 10812 32276 11466 32294
rect 10046 32266 10080 32270
rect 18156 32266 18190 32270
rect 9999 32222 18237 32236
rect 18258 32222 18292 35658
rect 9944 32202 18292 32222
rect 9944 32168 9978 32202
rect 18258 32168 18292 32202
rect 2036 31932 2484 32144
rect 3868 32134 20160 32168
rect 1498 31368 2136 31830
rect 2186 31742 2734 31776
rect 2186 31714 2220 31742
rect 2700 31714 2734 31742
rect 3868 31714 3902 32134
rect 4712 32066 4750 32104
rect 5470 32066 5508 32104
rect 6216 32066 6250 32134
rect 6260 32082 6266 32124
rect 4044 32032 4750 32066
rect 4802 32032 5508 32066
rect 5560 32032 6250 32066
rect 6177 31994 6178 31995
rect 6216 31994 6250 32032
rect 6302 32022 6308 32082
rect 6318 32032 6352 32134
rect 6314 32022 6352 32032
rect 6274 31998 6352 32022
rect 6256 31996 6352 31998
rect 6256 31994 6290 31996
rect 6302 31994 6308 31996
rect 6178 31993 6179 31994
rect 3971 31982 4016 31993
rect 4729 31982 4774 31993
rect 5487 31982 5532 31993
rect 3982 31714 4016 31982
rect 4027 31726 4028 31727
rect 4728 31726 4729 31727
rect 4028 31725 4029 31726
rect 4727 31725 4728 31726
rect 4740 31714 4774 31982
rect 4785 31726 4786 31727
rect 5486 31726 5487 31727
rect 4786 31725 4787 31726
rect 5485 31725 5486 31726
rect 5498 31714 5532 31982
rect 6216 31968 6296 31994
rect 6216 31742 6290 31968
rect 5543 31726 5544 31727
rect 6222 31726 6290 31742
rect 5544 31725 5545 31726
rect 6166 31714 6177 31725
rect 2186 31680 2254 31714
rect 2334 31696 2586 31700
rect 2332 31680 2588 31696
rect 2186 31676 2220 31680
rect 2332 31676 2364 31680
rect 2186 31674 2364 31676
rect 2558 31674 2588 31680
rect 2700 31680 2768 31714
rect 3834 31680 6177 31714
rect 2186 31460 2220 31674
rect 2360 31662 2560 31668
rect 2360 31656 2364 31662
rect 2250 31648 2364 31656
rect 2236 31646 2364 31648
rect 2372 31656 2560 31662
rect 2372 31646 2670 31656
rect 2250 31624 2360 31646
rect 2372 31628 2559 31646
rect 2560 31624 2670 31646
rect 2250 31622 2670 31624
rect 2250 31618 2360 31622
rect 2560 31618 2670 31622
rect 2288 31596 2360 31618
rect 2288 31594 2588 31596
rect 2288 31584 2360 31594
rect 2361 31574 2559 31585
rect 2598 31584 2670 31618
rect 2372 31540 2559 31574
rect 2700 31460 2734 31680
rect 2186 31426 2734 31460
rect 3868 31056 3902 31680
rect 3982 31056 4016 31680
rect 4028 31668 4029 31669
rect 4727 31668 4728 31669
rect 4027 31667 4028 31668
rect 4728 31667 4729 31668
rect 4027 31068 4028 31069
rect 4728 31068 4729 31069
rect 4028 31067 4029 31068
rect 4727 31067 4728 31068
rect 4740 31056 4774 31680
rect 4786 31668 4787 31669
rect 5485 31668 5486 31669
rect 4785 31667 4786 31668
rect 5486 31667 5487 31668
rect 4810 31078 4814 31090
rect 4785 31068 4786 31069
rect 4786 31067 4787 31068
rect 4822 31056 4826 31078
rect 5486 31068 5487 31069
rect 5485 31067 5486 31068
rect 5498 31056 5532 31680
rect 5544 31668 5545 31669
rect 6178 31668 6250 31690
rect 6256 31668 6290 31726
rect 5543 31667 5544 31668
rect 6178 31652 6290 31668
rect 6216 31084 6290 31652
rect 5543 31068 5544 31069
rect 6222 31068 6290 31084
rect 5544 31067 5545 31068
rect 6166 31056 6177 31067
rect 3834 31022 6177 31056
rect 2102 30828 2234 30946
rect 2034 30763 2482 30828
rect 3868 30763 3902 31022
rect 3982 30763 4016 31022
rect 4028 31010 4029 31011
rect 4727 31010 4728 31011
rect 4027 31009 4028 31010
rect 4728 31009 4729 31010
rect 4632 30980 4692 30994
rect 4740 30763 4774 31022
rect 4786 31010 4787 31011
rect 5485 31010 5486 31011
rect 4785 31009 4786 31010
rect 5486 31009 5487 31010
rect 4816 30980 4878 30994
rect 5382 30980 5492 30994
rect 5498 30763 5532 31022
rect 5544 31010 5545 31011
rect 6178 31010 6250 31032
rect 6256 31010 6290 31068
rect 5543 31009 5544 31010
rect 6178 30994 6290 31010
rect 5538 30980 5648 30994
rect 6216 30763 6290 30994
rect 6314 30763 6352 31996
rect -2027 29556 6411 30763
rect -1991 26860 -1957 29556
rect 3832 29303 6411 29556
rect -1808 29284 -1508 29303
rect -156 29284 1344 29303
rect 2912 29286 6411 29303
rect 3484 29186 3496 29252
rect 3726 29174 3742 29252
rect -1564 29158 -100 29174
rect 1534 29106 2100 29140
rect 1534 28784 1568 29106
rect 2066 29042 2100 29106
rect 2150 29042 2770 29158
rect 1718 29026 1916 29037
rect 1589 28964 1717 29011
rect 1729 28992 1916 29026
rect 2002 29011 2770 29042
rect 1917 28964 2770 29011
rect 1636 28926 1717 28964
rect 1964 28926 2770 28964
rect 1718 28898 1916 28909
rect 1974 28900 2770 28926
rect 1729 28864 1916 28898
rect 2002 28830 2770 28900
rect 2066 28784 2100 28830
rect 1534 28750 2100 28784
rect 2150 28736 2770 28830
rect 2010 28184 2458 28396
rect 2102 28174 2234 28184
rect 3832 28073 6411 29286
rect -1916 28062 6411 28073
rect -1905 28050 6411 28062
rect -1916 28039 6411 28050
rect -1889 27993 -1855 28039
rect -980 27981 -524 28000
rect 3832 27981 6411 28039
rect -1796 27925 6411 27981
rect -1889 27329 -1855 27919
rect -942 27910 -486 27925
rect 2010 27720 2458 27730
rect 2002 27518 2458 27720
rect 2002 27508 2450 27518
rect 1144 27323 3276 27334
rect 3832 27323 6411 27925
rect 7014 27434 7048 31982
rect 9288 27434 9322 31982
rect 9944 30719 9978 32134
rect 13350 32130 13636 32134
rect 10046 32100 10056 32104
rect 10070 32100 10080 32104
rect 10008 32032 10034 32066
rect 10046 31998 10080 32100
rect 10776 32066 10814 32104
rect 11534 32066 11572 32104
rect 12292 32066 12330 32104
rect 13050 32066 13088 32104
rect 13384 32066 13602 32116
rect 13808 32100 13846 32104
rect 13808 32066 14260 32100
rect 14566 32066 14604 32104
rect 14730 32066 14952 32104
rect 15324 32066 15362 32104
rect 16082 32066 16120 32104
rect 16840 32066 16878 32104
rect 17598 32066 17636 32104
rect 18156 32066 18190 32134
rect 18258 32066 18292 32134
rect 10092 32032 10814 32066
rect 10866 32032 11572 32066
rect 11624 32032 12330 32066
rect 12382 32032 13088 32066
rect 13140 32032 14604 32066
rect 14656 32032 15362 32066
rect 15414 32032 16120 32066
rect 16172 32032 16878 32066
rect 16930 32032 17636 32066
rect 17688 32032 18292 32066
rect 10046 31994 10056 31998
rect 10070 31994 10080 31998
rect 10118 31994 10119 31995
rect 10034 31682 10092 31994
rect 10117 31993 10118 31994
rect 10793 31982 10838 31993
rect 11551 31982 11596 31993
rect 12309 31982 12354 31993
rect 13067 31982 13112 31993
rect 10792 31682 10793 31683
rect 10791 31681 10792 31682
rect 10804 31670 10838 31982
rect 10849 31682 10850 31683
rect 11550 31682 11551 31683
rect 10850 31681 10851 31682
rect 11549 31681 11550 31682
rect 11562 31670 11596 31982
rect 11607 31682 11608 31683
rect 12308 31682 12309 31683
rect 11608 31681 11609 31682
rect 12307 31681 12308 31682
rect 12320 31670 12354 31982
rect 12365 31682 12366 31683
rect 13066 31682 13067 31683
rect 12366 31681 12367 31682
rect 13065 31681 13066 31682
rect 13078 31670 13112 31982
rect 13812 31888 14260 32032
rect 18117 31994 18118 31995
rect 18118 31993 18119 31994
rect 14583 31982 14628 31993
rect 15341 31982 15386 31993
rect 16099 31982 16144 31993
rect 16857 31982 16902 31993
rect 17615 31982 17660 31993
rect 13710 31732 13736 31768
rect 13738 31732 13764 31768
rect 13836 31732 13870 31888
rect 14594 31786 14628 31982
rect 13562 31698 14110 31732
rect 13123 31682 13124 31683
rect 13124 31681 13125 31682
rect 13562 31681 13596 31698
rect 13384 31670 13602 31681
rect 13710 31676 13736 31698
rect 13738 31676 13764 31698
rect 13824 31682 13825 31683
rect 13823 31681 13824 31682
rect 13836 31670 13870 31698
rect 13881 31682 13882 31683
rect 13882 31681 13883 31682
rect 14076 31670 14110 31698
rect 14160 31681 14798 31786
rect 15340 31682 15341 31683
rect 15339 31681 15340 31682
rect 14160 31670 14952 31681
rect 15352 31670 15386 31982
rect 15397 31682 15398 31683
rect 16098 31682 16099 31683
rect 15398 31681 15399 31682
rect 16097 31681 16098 31682
rect 16110 31670 16144 31982
rect 16155 31682 16156 31683
rect 16856 31682 16857 31683
rect 16156 31681 16157 31682
rect 16855 31681 16856 31682
rect 16868 31670 16902 31982
rect 16913 31682 16914 31683
rect 17614 31682 17615 31683
rect 16914 31681 16915 31682
rect 17613 31681 17614 31682
rect 17626 31670 17660 31982
rect 18156 31698 18190 32032
rect 17671 31682 17672 31683
rect 17672 31681 17673 31682
rect 18106 31670 18117 31681
rect 10130 31636 18117 31670
rect 10791 31624 10792 31625
rect 10034 31024 10092 31624
rect 10792 31623 10793 31624
rect 10804 31168 10838 31636
rect 10850 31624 10851 31625
rect 11549 31624 11550 31625
rect 10849 31623 10850 31624
rect 11550 31623 11551 31624
rect 10758 31034 10878 31168
rect 10758 31020 11474 31034
rect 11550 31024 11551 31025
rect 11549 31023 11550 31024
rect 10804 31012 11474 31020
rect 11562 31012 11596 31636
rect 11608 31624 11609 31625
rect 12307 31624 12308 31625
rect 11607 31623 11608 31624
rect 12308 31623 12309 31624
rect 11607 31024 11608 31025
rect 12308 31024 12309 31025
rect 11608 31023 11609 31024
rect 12307 31023 12308 31024
rect 12320 31012 12354 31636
rect 12366 31624 12367 31625
rect 13065 31624 13066 31625
rect 12365 31623 12366 31624
rect 13066 31623 13067 31624
rect 12365 31024 12366 31025
rect 13066 31024 13067 31025
rect 12366 31023 12367 31024
rect 13065 31023 13066 31024
rect 13078 31012 13112 31636
rect 13124 31624 13125 31625
rect 13123 31623 13124 31624
rect 13562 31416 13596 31636
rect 13736 31630 13738 31636
rect 13710 31624 13736 31630
rect 13738 31624 13764 31630
rect 13823 31624 13824 31625
rect 13736 31618 13738 31624
rect 13824 31623 13825 31624
rect 13836 31618 13870 31636
rect 13932 31632 13964 31636
rect 13932 31630 13980 31632
rect 13882 31624 13883 31625
rect 13924 31624 13935 31629
rect 13881 31623 13882 31624
rect 13924 31618 13936 31624
rect 13732 31612 13940 31618
rect 13626 31574 13698 31612
rect 13732 31602 14008 31612
rect 13748 31584 13935 31602
rect 13736 31578 13796 31580
rect 13664 31540 13698 31574
rect 13736 31550 13796 31552
rect 13836 31530 13870 31584
rect 13936 31580 14008 31602
rect 13920 31578 14008 31580
rect 13936 31574 14008 31578
rect 13920 31550 13964 31552
rect 13924 31530 13935 31541
rect 13974 31540 14008 31574
rect 13748 31496 13935 31530
rect 13836 31416 13870 31496
rect 14076 31416 14110 31636
rect 13562 31382 14110 31416
rect 13836 31226 13870 31382
rect 14160 31324 14798 31636
rect 15339 31624 15340 31625
rect 15340 31623 15341 31624
rect 13818 31220 13932 31226
rect 13123 31024 13124 31025
rect 13824 31024 13825 31025
rect 13124 31023 13125 31024
rect 13823 31023 13824 31024
rect 13836 31012 13870 31220
rect 13881 31024 13882 31025
rect 14582 31024 14583 31025
rect 13882 31023 13883 31024
rect 14581 31023 14582 31024
rect 14594 31012 14628 31324
rect 14639 31024 14640 31025
rect 15340 31024 15341 31025
rect 14640 31023 14641 31024
rect 15339 31023 15340 31024
rect 15352 31012 15386 31636
rect 15398 31624 15399 31625
rect 16097 31624 16098 31625
rect 15397 31623 15398 31624
rect 16098 31623 16099 31624
rect 15397 31024 15398 31025
rect 16098 31024 16099 31025
rect 15398 31023 15399 31024
rect 16097 31023 16098 31024
rect 16110 31012 16144 31636
rect 16156 31624 16157 31625
rect 16855 31624 16856 31625
rect 16155 31623 16156 31624
rect 16856 31623 16857 31624
rect 16155 31024 16156 31025
rect 16856 31024 16857 31025
rect 16156 31023 16157 31024
rect 16855 31023 16856 31024
rect 16868 31012 16902 31636
rect 16914 31624 16915 31625
rect 17613 31624 17614 31625
rect 16913 31623 16914 31624
rect 17614 31623 17615 31624
rect 16913 31024 16914 31025
rect 17614 31024 17615 31025
rect 16914 31023 16915 31024
rect 17613 31023 17614 31024
rect 17626 31012 17660 31636
rect 17672 31624 17673 31625
rect 17671 31623 17672 31624
rect 18118 31608 18190 31646
rect 18156 31040 18190 31608
rect 17671 31024 17672 31025
rect 17672 31023 17673 31024
rect 18106 31012 18117 31023
rect 10130 30978 18117 31012
rect 10791 30966 10792 30967
rect 10034 30719 10092 30966
rect 10792 30965 10793 30966
rect 10804 30960 11474 30978
rect 11549 30966 11550 30967
rect 11550 30965 11551 30966
rect 10706 30936 10754 30950
rect 10804 30719 10838 30960
rect 10878 30936 10950 30950
rect 11454 30936 11556 30950
rect 11562 30719 11596 30978
rect 11608 30966 11609 30967
rect 12307 30966 12308 30967
rect 11607 30965 11608 30966
rect 12308 30965 12309 30966
rect 11602 30936 11718 30950
rect 12320 30719 12354 30978
rect 12366 30966 12367 30967
rect 13065 30966 13066 30967
rect 12365 30965 12366 30966
rect 13066 30965 13067 30966
rect 13078 30719 13112 30978
rect 13124 30966 13125 30967
rect 13823 30966 13824 30967
rect 13123 30965 13124 30966
rect 13824 30965 13825 30966
rect 13836 30784 13870 30978
rect 13882 30966 13883 30967
rect 14581 30966 14582 30967
rect 13881 30965 13882 30966
rect 14582 30965 14583 30966
rect 14062 30784 14194 30902
rect 13814 30719 14262 30784
rect 14594 30719 14628 30978
rect 14640 30966 14641 30967
rect 15339 30966 15340 30967
rect 14639 30965 14640 30966
rect 15340 30965 15341 30966
rect 15352 30719 15386 30978
rect 15398 30966 15399 30967
rect 16097 30966 16098 30967
rect 15397 30965 15398 30966
rect 16098 30965 16099 30966
rect 16110 30719 16144 30978
rect 16156 30966 16157 30967
rect 16855 30966 16856 30967
rect 16155 30965 16156 30966
rect 16856 30965 16857 30966
rect 16868 30719 16902 30978
rect 16914 30966 16915 30967
rect 17613 30966 17614 30967
rect 16913 30965 16914 30966
rect 17614 30965 17615 30966
rect 17626 30719 17660 30978
rect 17672 30966 17673 30967
rect 17671 30965 17672 30966
rect 18118 30950 18190 30988
rect 18156 30719 18190 30950
rect 18258 30719 18292 32032
rect -1796 27267 6411 27323
rect -1889 27239 -1855 27243
rect 3832 27212 6411 27267
rect 9885 27212 18323 30719
rect 19900 27434 19934 31982
rect 21358 31386 27278 35606
rect 21358 31366 27318 31386
rect 21318 29282 21319 29283
rect 21317 29281 21318 29282
rect 21358 29242 27278 31366
rect 27280 30947 27281 31366
rect 27318 30947 27338 31366
rect 27280 30946 27338 30947
rect 27566 29294 27630 35658
rect 27747 33045 27781 39409
rect 27911 39363 27978 39376
rect 28426 39363 28503 39376
rect 28569 39363 28636 39376
rect 29084 39363 29161 39376
rect 29227 39363 29298 39376
rect 29746 39363 29819 39376
rect 29885 39363 29968 39376
rect 30416 39363 30477 39376
rect 30543 39363 30620 39376
rect 31068 39363 31135 39376
rect 29177 36851 29211 39310
rect 30493 36851 30527 39310
rect 27849 36817 31197 36851
rect 27861 36783 27895 36817
rect 28519 36796 28553 36817
rect 29177 36796 29211 36817
rect 29835 36796 29869 36817
rect 30493 36796 30527 36817
rect 31151 36796 31185 36817
rect 28491 36783 28553 36796
rect 29149 36783 29211 36796
rect 29807 36783 29869 36796
rect 30465 36783 30527 36796
rect 27861 36681 27901 36783
rect 28491 36755 28559 36783
rect 29149 36755 29217 36783
rect 29807 36755 29875 36783
rect 30465 36755 30533 36783
rect 31123 36755 31185 36796
rect 27911 36749 27929 36755
rect 28485 36749 28559 36755
rect 28569 36749 28587 36755
rect 29143 36749 29217 36755
rect 29227 36749 29245 36755
rect 29801 36749 29875 36755
rect 29885 36749 29903 36755
rect 30459 36749 30533 36755
rect 30543 36749 30561 36755
rect 31117 36749 31185 36755
rect 27907 36715 28559 36749
rect 28565 36715 29217 36749
rect 29223 36715 29875 36749
rect 29881 36715 30533 36749
rect 30539 36715 31185 36749
rect 27911 36709 27929 36715
rect 28485 36709 28503 36715
rect 28513 36681 28559 36715
rect 28569 36709 28587 36715
rect 29143 36709 29161 36715
rect 29171 36681 29217 36715
rect 29227 36709 29245 36715
rect 29801 36709 29819 36715
rect 29829 36681 29875 36715
rect 29885 36709 29903 36715
rect 30459 36709 30477 36715
rect 30487 36681 30533 36715
rect 30543 36709 30561 36715
rect 31117 36709 31135 36715
rect 31145 36681 31185 36715
rect 27861 33141 27895 36681
rect 28420 35610 28426 36134
rect 28519 33141 28553 36681
rect 29177 35796 29211 36681
rect 29835 35796 29869 36681
rect 28840 35504 30322 35796
rect 28756 35056 30322 35504
rect 28840 34862 30322 35056
rect 30493 34862 30527 36681
rect 31108 35610 31124 36078
rect 28840 34490 30894 34862
rect 28840 34220 30322 34490
rect 29177 33141 29211 34220
rect 29835 33141 29869 34220
rect 30493 33141 30527 34490
rect 31151 33141 31185 36681
rect 27811 33107 27815 33141
rect 27849 33107 31197 33141
rect 27861 33086 27895 33107
rect 28519 33086 28553 33107
rect 29177 33086 29211 33107
rect 29835 33086 29869 33107
rect 30493 33086 30527 33107
rect 27715 32204 27781 33045
rect 27849 33039 30750 33086
rect 31091 33039 31138 33086
rect 27861 33005 28506 33039
rect 28519 33005 29164 33039
rect 29177 33005 29822 33039
rect 29835 33005 30480 33039
rect 30493 33005 31138 33039
rect 27861 32958 27907 33005
rect 27936 32999 27946 33005
rect 28426 32999 28471 33005
rect 28519 32999 28604 33005
rect 29084 32999 29129 33005
rect 27817 32946 27835 32958
rect 27861 32946 27906 32958
rect 27918 32956 27936 32999
rect 27946 32956 27964 32999
rect 28519 32958 28565 32999
rect 29136 32971 29157 33005
rect 29177 32958 29223 33005
rect 29244 32999 29266 33005
rect 29746 32999 29787 33005
rect 29835 32999 29936 33005
rect 30416 32999 30445 33005
rect 28476 32946 28507 32957
rect 28519 32946 28564 32958
rect 29134 32946 29165 32957
rect 29177 32946 29222 32958
rect 29238 32956 29244 32999
rect 29266 32956 29272 32999
rect 29835 32958 29881 32999
rect 30456 32971 30473 33005
rect 30493 32958 30539 33005
rect 30564 32999 30588 33005
rect 31068 32999 31103 33005
rect 29792 32946 29823 32957
rect 29835 32946 29880 32958
rect 30450 32946 30481 32957
rect 30493 32946 30538 32958
rect 30560 32956 30564 32999
rect 30588 32956 30592 32999
rect 31108 32946 31139 32957
rect 31151 32946 31185 33107
rect 27817 32204 27906 32946
rect 28487 32204 28564 32946
rect 29145 32204 29222 32946
rect 29803 32204 29880 32946
rect 30461 32204 30538 32946
rect 19204 27350 20160 27384
rect 6239 27209 6273 27212
rect -1927 27175 6311 27209
rect 6239 27020 6273 27175
rect 6239 26934 6328 27020
rect 6239 26860 6273 26934
rect -2027 25788 6388 26860
rect 9921 26532 9955 27212
rect 10008 27165 10628 27212
rect 10678 27165 10712 27212
rect 10812 27202 11466 27212
rect 11210 27165 11244 27202
rect 18151 27195 18185 27199
rect 9985 27131 18219 27165
rect 10008 27122 10628 27131
rect 9985 27036 10628 27122
rect 10008 26852 10628 27036
rect 10678 26904 10712 27131
rect 10718 27130 10860 27131
rect 10873 27130 11142 27131
rect 10733 27084 10814 27130
rect 10873 27112 11060 27130
rect 11061 27084 11142 27130
rect 10780 27046 10814 27084
rect 11108 27046 11142 27084
rect 11049 27018 11060 27029
rect 10873 26984 11060 27018
rect 11210 26904 11244 27131
rect 10678 26870 11244 26904
rect 10416 26698 10518 26714
rect 11056 26698 11462 26700
rect 9985 26589 10012 26646
rect 10023 26627 10050 26684
rect 10444 26670 10518 26686
rect 11056 26670 11434 26672
rect 9985 26560 10012 26575
rect 10116 26565 18092 26599
rect 9921 26502 10017 26532
rect 10023 26522 10050 26537
rect 10063 26502 10414 26532
rect 10444 26522 10718 26532
rect 9921 26486 9955 26502
rect 10063 26486 10244 26502
rect 10444 26486 10644 26522
rect 10860 26486 11434 26532
rect 16452 26516 17804 26532
rect 18253 26486 18287 27212
rect 9885 25824 18287 26486
rect 9866 25788 18287 25824
rect -2027 25754 18287 25788
rect -18495 21973 -18461 24531
rect -2027 24485 6388 25754
rect -20160 21939 -15721 21973
rect -18495 21859 -18461 21939
rect -18393 21893 -18359 21939
rect -15755 21881 -15721 21939
rect -18440 21859 -18359 21866
rect -18300 21859 -15721 21881
rect -18529 21847 -15721 21859
rect -18529 21835 -15916 21847
rect -18529 21825 -15905 21835
rect -18495 21201 -18461 21825
rect -18440 21819 -18312 21825
rect -18409 21813 -18312 21819
rect -18393 21251 -18359 21813
rect -15904 21797 -15823 21844
rect -15857 21235 -15823 21797
rect -15904 21223 -15807 21235
rect -15755 21223 -15721 21847
rect -1996 21789 -1962 24485
rect 3944 24170 4350 24485
rect 4594 24170 6388 24485
rect -1921 24159 6388 24170
rect -1910 24147 6388 24159
rect -1921 24136 6388 24147
rect -1894 24090 -1860 24136
rect -880 24090 -422 24110
rect -880 24078 -382 24090
rect 3944 24078 4350 24136
rect 4594 24078 6388 24136
rect -1810 24022 6388 24078
rect -880 24018 -382 24022
rect -1894 23426 -1860 24016
rect -840 23998 -382 24018
rect -1230 23974 -126 23994
rect -1258 23946 -98 23966
rect 3786 23960 3842 23966
rect 4470 23960 4526 23966
rect 2030 23814 2478 23842
rect 2030 23630 2496 23814
rect 2048 23602 2496 23630
rect 4480 23434 4526 23458
rect 4594 23431 6388 24022
rect 1144 23420 6388 23431
rect -1810 23364 6388 23420
rect -1894 23336 -1860 23340
rect 4594 23306 6388 23364
rect -1941 23272 6388 23306
rect 2036 22958 2484 23170
rect 1498 22394 2136 22856
rect 2186 22768 2734 22802
rect 2186 22740 2220 22768
rect 2700 22740 2734 22768
rect 2186 22706 2254 22740
rect 2334 22722 2586 22726
rect 2332 22706 2588 22722
rect 2186 22702 2220 22706
rect 2332 22702 2364 22706
rect 2186 22700 2364 22702
rect 2558 22700 2588 22706
rect 2700 22706 2768 22740
rect 2186 22486 2220 22700
rect 2360 22688 2560 22694
rect 2360 22682 2364 22688
rect 2250 22674 2364 22682
rect 2236 22672 2364 22674
rect 2372 22682 2560 22688
rect 2372 22672 2670 22682
rect 2250 22650 2360 22672
rect 2372 22654 2559 22672
rect 2560 22650 2670 22672
rect 2250 22648 2670 22650
rect 2250 22644 2360 22648
rect 2560 22644 2670 22648
rect 2288 22622 2360 22644
rect 2288 22620 2588 22622
rect 2288 22610 2360 22620
rect 2361 22600 2559 22611
rect 2598 22610 2670 22644
rect 2372 22566 2559 22600
rect 2700 22486 2734 22706
rect 2186 22452 2734 22486
rect 4594 22020 6388 23272
rect 4474 22006 6388 22020
rect 2102 21854 2234 21972
rect 2034 21789 2482 21854
rect 4594 21789 6388 22006
rect -18300 21201 -15721 21223
rect -18495 21189 -15721 21201
rect -18495 21167 -15916 21189
rect -15904 21177 -15776 21186
rect -18495 21109 -18461 21167
rect -15857 21139 -15823 21143
rect -15755 21109 -15721 21189
rect -18495 21075 -10225 21109
rect -15755 20160 -15721 21075
rect -2027 20582 6388 21789
rect 9866 24511 18287 25754
rect 21326 27032 27278 29242
rect 9866 24441 18286 24511
rect 9866 24134 14102 24441
rect 9866 23922 14220 24134
rect 9866 23796 14102 23922
rect 9866 23785 18175 23796
rect 9866 23773 18164 23785
rect 9866 23762 18175 23773
rect 9866 23704 14102 23762
rect 16676 23716 17134 23736
rect 18114 23716 18148 23762
rect 16636 23704 17134 23716
rect 9866 23658 18064 23704
rect 9866 23648 18075 23658
rect 9866 23468 14102 23648
rect 16636 23644 17134 23648
rect 16636 23624 17094 23644
rect 16380 23600 17484 23620
rect 16352 23572 17512 23592
rect 9866 23256 14224 23468
rect 9866 23228 14206 23256
rect 9866 23046 14102 23228
rect 18064 23046 18075 23057
rect 18114 23052 18148 23642
rect 9866 23036 18075 23046
rect 9866 22990 18064 23036
rect 9866 22932 14102 22990
rect 18114 22962 18148 22966
rect 9866 22898 18182 22932
rect 9866 22796 14102 22898
rect 9866 22584 14218 22796
rect 9866 21598 14102 22584
rect 14118 22020 14756 22482
rect 18114 21736 18148 22304
rect 17472 21674 18172 21708
rect 9866 21480 14152 21598
rect 18114 21510 18148 21646
rect 18216 21510 18250 24441
rect 21286 22610 21287 22611
rect 21285 22609 21286 22610
rect 21326 22570 27246 27032
rect 27286 26992 27287 26993
rect 27285 26991 27286 26992
rect 27534 26980 27630 29294
rect 27679 32030 30696 32204
rect 27679 31836 30894 32030
rect 27679 31322 30696 31836
rect 31119 31768 31185 32946
rect 31233 33045 31251 33107
rect 31265 33045 31299 39409
rect 32130 35650 32166 35666
rect 32818 33050 32852 39414
rect 32982 39368 33064 39376
rect 33512 39368 33574 39376
rect 33640 39368 33716 39376
rect 34164 39368 34232 39376
rect 34298 39368 34374 39376
rect 34822 39368 34890 39376
rect 34956 39368 35038 39376
rect 35486 39368 35548 39376
rect 35614 39368 35690 39376
rect 36138 39368 36206 39376
rect 32920 36822 36268 36856
rect 32932 36788 32966 36822
rect 33590 36792 33624 36822
rect 34248 36792 34282 36822
rect 34906 36792 34940 36822
rect 35564 36792 35598 36822
rect 36222 36792 36256 36822
rect 33562 36788 33624 36792
rect 32932 36686 32972 36788
rect 33562 36760 33630 36788
rect 34220 36760 35228 36792
rect 35536 36788 35598 36792
rect 35536 36760 35604 36788
rect 36194 36760 36256 36792
rect 32982 36754 33000 36760
rect 33556 36754 33630 36760
rect 33640 36754 33658 36760
rect 34214 36754 35228 36760
rect 35530 36754 35604 36760
rect 35614 36754 35632 36760
rect 36188 36754 36256 36760
rect 32978 36720 33630 36754
rect 33636 36720 34288 36754
rect 32982 36714 33000 36720
rect 33556 36714 33574 36720
rect 33584 36686 33630 36720
rect 33640 36714 33658 36720
rect 34214 36714 34232 36720
rect 34242 36686 34288 36720
rect 34298 36720 34946 36754
rect 34298 36714 34316 36720
rect 34872 36714 34890 36720
rect 34900 36686 34946 36720
rect 34956 36720 35604 36754
rect 35610 36720 36256 36754
rect 34956 36714 34974 36720
rect 35530 36714 35548 36720
rect 35558 36686 35604 36720
rect 35614 36714 35632 36720
rect 36188 36714 36206 36720
rect 36216 36686 36256 36720
rect 32932 33146 32966 36686
rect 33590 33146 33624 36686
rect 34248 33146 34282 36686
rect 34906 33146 34940 36686
rect 35564 33146 35598 36686
rect 36222 33146 36256 36686
rect 32882 33112 32886 33146
rect 32920 33112 36268 33146
rect 32932 33082 32966 33112
rect 33590 33082 33624 33112
rect 34248 33082 34282 33112
rect 34906 33082 34940 33112
rect 35564 33082 35598 33112
rect 31233 32204 31299 33045
rect 31048 31322 31068 31768
rect 31076 31322 31185 31768
rect 27679 31241 31185 31322
rect 27679 31173 30696 31241
rect 31107 31225 31185 31241
rect 31113 31173 31185 31225
rect 27679 31139 31219 31173
rect 27679 30487 30696 31139
rect 31113 30794 31185 31139
rect 31119 30521 31185 30794
rect 31119 30487 31205 30521
rect 27679 30453 31205 30487
rect 27679 30385 30696 30453
rect 31119 30432 31185 30453
rect 31091 30385 31185 30432
rect 27679 30351 31185 30385
rect 27679 28621 30696 30351
rect 31048 28938 31068 29606
rect 31076 28938 31096 29606
rect 31119 28680 31185 30351
rect 31119 28668 31153 28680
rect 31107 28621 31165 28668
rect 27679 28587 31165 28621
rect 27679 28519 30696 28587
rect 31107 28571 31153 28587
rect 27679 28485 31165 28519
rect 27679 27212 30696 28485
rect 27534 22622 27598 26980
rect 27715 26373 27749 27212
rect 27829 26469 27863 27212
rect 28487 26469 28521 27212
rect 29145 26469 29179 27212
rect 29803 26469 29837 27212
rect 30066 26469 30278 26486
rect 30461 26469 30495 27212
rect 31119 26469 31153 28485
rect 31232 28449 31335 32204
rect 32786 32168 32852 33050
rect 32928 33044 33568 33082
rect 33586 33044 34226 33082
rect 34244 33044 34884 33082
rect 34902 33044 35542 33082
rect 35560 33044 36200 33082
rect 32932 33010 33568 33044
rect 33590 33040 34226 33044
rect 33590 33010 34228 33040
rect 32932 32972 32978 33010
rect 33004 33004 33032 33010
rect 33512 33004 33542 33010
rect 33590 33004 33684 33010
rect 34164 33004 34200 33010
rect 33590 32972 33636 33004
rect 34206 32976 34228 33010
rect 34248 33010 34884 33044
rect 34906 33010 35542 33044
rect 35564 33010 36200 33044
rect 34248 32972 34294 33010
rect 34314 33004 34342 33010
rect 34822 33004 34858 33010
rect 34906 33004 35006 33010
rect 35486 33004 35516 33010
rect 34906 32972 34952 33004
rect 35528 32976 35544 33004
rect 35564 32972 35610 33010
rect 35636 33004 35658 33010
rect 36138 33004 36174 33010
rect 32888 32960 32906 32972
rect 32932 32960 32977 32972
rect 33547 32960 33578 32971
rect 33590 32960 33635 32972
rect 34205 32960 34236 32971
rect 34248 32960 34293 32972
rect 34863 32960 34894 32971
rect 34906 32960 34951 32972
rect 35521 32960 35552 32971
rect 35564 32960 35609 32972
rect 32888 32168 32977 32960
rect 33558 32168 33635 32960
rect 34216 32168 34293 32960
rect 34874 32168 34951 32960
rect 35532 32168 35609 32960
rect 35630 32956 35636 33004
rect 35658 32956 35664 33004
rect 36179 32960 36210 32971
rect 36222 32960 36256 33112
rect 36190 32168 36256 32960
rect 36304 33050 36322 33112
rect 36336 33050 36370 39414
rect 74317 38203 74383 40013
rect 74459 40023 74463 40041
rect 74459 40007 74509 40023
rect 74520 40013 74538 40028
rect 74548 40013 74566 40026
rect 75061 40007 75108 40054
rect 75117 40023 75121 40041
rect 75117 40007 75167 40023
rect 75719 40013 75766 40054
rect 75710 40007 75766 40013
rect 75775 40023 75779 40041
rect 75775 40007 75825 40023
rect 75840 40013 75846 40016
rect 75868 40013 75874 40026
rect 76377 40007 76424 40054
rect 76433 40023 76437 40041
rect 76433 40007 76483 40023
rect 77035 40013 77082 40054
rect 77030 40007 77082 40013
rect 77091 40023 77095 40041
rect 77091 40007 77141 40023
rect 77693 40007 77740 40054
rect 74463 39973 75108 40007
rect 75121 39973 75766 40007
rect 75779 39973 76424 40007
rect 76437 39973 77082 40007
rect 77095 39973 77740 40007
rect 74463 39926 74509 39973
rect 74419 39914 74437 39926
rect 74463 39914 74497 39926
rect 74419 38302 74497 39914
rect 74520 38626 74538 39967
rect 74548 38598 74566 39967
rect 75121 39926 75167 39973
rect 75710 39967 75731 39973
rect 75738 39939 75759 39973
rect 75779 39926 75825 39973
rect 75078 39914 75109 39925
rect 75121 39914 75155 39926
rect 75736 39914 75767 39925
rect 75779 39914 75813 39926
rect 74317 36394 74351 38203
rect 74419 38141 74465 38302
rect 75018 38249 75028 39648
rect 75046 38277 75056 39620
rect 75089 38302 75155 39914
rect 75747 38302 75813 39914
rect 75840 38614 75846 39967
rect 75868 38586 75874 39967
rect 76437 39926 76483 39973
rect 77030 39967 77047 39973
rect 77058 39939 77075 39973
rect 77095 39926 77141 39973
rect 76394 39914 76425 39925
rect 76437 39914 76471 39926
rect 77052 39914 77083 39925
rect 77095 39914 77129 39926
rect 75089 38290 75123 38302
rect 75747 38290 75781 38302
rect 75077 38277 75136 38290
rect 75046 38268 75136 38277
rect 75143 38268 75174 38277
rect 75077 38249 75136 38268
rect 75018 38243 75136 38249
rect 74525 38209 75136 38243
rect 75171 38243 75202 38249
rect 75735 38243 75794 38290
rect 76328 38249 76348 39654
rect 76356 38277 76376 39626
rect 76405 38302 76471 39914
rect 77063 38302 77129 39914
rect 77162 38592 77166 39967
rect 77190 38564 77194 39967
rect 77710 39914 77741 39925
rect 77753 39914 77787 40075
rect 76405 38290 76439 38302
rect 77063 38290 77097 38302
rect 76393 38277 76452 38290
rect 76356 38274 76452 38277
rect 76459 38274 76484 38277
rect 76393 38249 76452 38274
rect 76328 38246 76452 38249
rect 76487 38246 76512 38249
rect 76393 38243 76452 38246
rect 77051 38243 77110 38290
rect 77650 38249 77670 39624
rect 77678 38249 77698 39596
rect 77721 38302 77787 39914
rect 77835 40013 77853 40075
rect 77867 40013 77901 40320
rect 79420 40018 79454 40320
rect 79534 40114 79568 40148
rect 80192 40114 80226 40148
rect 80850 40114 80884 40148
rect 81508 40114 81542 40148
rect 82166 40114 82200 40148
rect 82824 40114 82878 40148
rect 79484 40080 79488 40114
rect 79500 40080 82878 40114
rect 77721 38290 77755 38302
rect 77709 38243 77767 38290
rect 75171 38240 75794 38243
rect 75183 38209 75794 38240
rect 75841 38209 76452 38243
rect 76499 38209 77110 38243
rect 77157 38209 77767 38243
rect 75077 38193 75123 38209
rect 75735 38193 75781 38209
rect 76393 38193 76439 38209
rect 77051 38193 77097 38209
rect 77709 38193 77755 38209
rect 77835 38203 77901 40013
rect 79388 38226 79454 40018
rect 79530 40028 79534 40046
rect 79530 40012 79580 40028
rect 80132 40012 80170 40050
rect 80188 40028 80192 40046
rect 80188 40012 80238 40028
rect 80790 40018 80828 40050
rect 80780 40012 80828 40018
rect 80846 40028 80850 40046
rect 80846 40012 80896 40028
rect 81448 40012 81486 40050
rect 81504 40028 81508 40046
rect 81504 40012 81554 40028
rect 82106 40012 82144 40050
rect 82162 40028 82166 40046
rect 82162 40012 82212 40028
rect 82764 40012 82802 40050
rect 79534 39978 80170 40012
rect 80192 40008 80828 40012
rect 80192 39978 80830 40008
rect 79534 39940 79580 39978
rect 80192 39940 80238 39978
rect 80780 39972 80802 39978
rect 80808 39944 80830 39978
rect 80850 39978 81486 40012
rect 81508 39978 82144 40012
rect 82166 39978 82802 40012
rect 80850 39940 80896 39978
rect 81508 39940 81554 39978
rect 82102 39972 82118 39978
rect 82130 39944 82146 39972
rect 82166 39940 82212 39978
rect 79490 39928 79508 39940
rect 79534 39928 79568 39940
rect 80149 39928 80180 39939
rect 80192 39928 80226 39940
rect 80807 39928 80838 39939
rect 80850 39928 80884 39940
rect 81465 39928 81496 39939
rect 81508 39928 81542 39940
rect 82123 39928 82154 39939
rect 82166 39928 82200 39940
rect 79490 38316 79568 39928
rect 77063 38141 77097 38193
rect 74419 38107 77767 38141
rect 77063 36394 77097 38107
rect 77835 36394 77869 38203
rect 74317 36356 77869 36394
rect 52150 35496 52156 35508
rect 52342 35496 52350 35508
rect 52122 35468 52156 35480
rect 52342 35468 52378 35480
rect 51612 35044 52178 35078
rect 51612 34949 51646 35044
rect 51983 34964 51994 34975
rect 51807 34961 51994 34964
rect 51807 34949 51983 34961
rect 52144 34949 52178 35044
rect 51578 34915 52178 34949
rect 51612 34722 51646 34915
rect 51667 34903 51795 34915
rect 51995 34903 52092 34915
rect 51667 34902 51748 34903
rect 51995 34902 52076 34903
rect 51714 34864 51748 34902
rect 52042 34864 52076 34902
rect 51704 34838 51756 34850
rect 51983 34836 51994 34847
rect 51676 34810 51784 34822
rect 51807 34802 51994 34836
rect 52128 34822 52130 34909
rect 52144 34722 52178 34915
rect 51612 34688 52178 34722
rect 52228 34887 52848 35092
rect 56986 34890 57116 34911
rect 52228 34670 52875 34887
rect 56800 34865 57116 34890
rect 57302 34865 57708 34911
rect 56828 34837 57116 34862
rect 57302 34837 57652 34862
rect 52841 34616 52875 34670
rect 51612 34568 52178 34602
rect 51612 34280 51646 34568
rect 51983 34488 51994 34499
rect 51667 34426 51748 34473
rect 51807 34454 51994 34488
rect 51995 34426 52076 34473
rect 51714 34388 51748 34426
rect 52042 34388 52076 34426
rect 52144 34374 52178 34568
rect 51983 34360 51994 34371
rect 52110 34360 52130 34374
rect 51807 34326 51994 34360
rect 52034 34346 52130 34360
rect 52138 34360 52178 34374
rect 52228 34464 52875 34616
rect 52228 34378 52930 34464
rect 52228 34360 52875 34378
rect 52138 34340 52875 34360
rect 52144 34332 52178 34340
rect 52228 34332 52875 34340
rect 52006 34319 52875 34332
rect 52006 34318 52848 34319
rect 52110 34312 52848 34318
rect 51769 34288 52021 34291
rect 52144 34280 52178 34312
rect 51612 34257 52178 34280
rect 51612 34246 51646 34257
rect 52144 34246 52178 34257
rect 51612 34245 52178 34246
rect 51646 34231 52144 34245
rect 51612 34212 52178 34231
rect 52228 34194 52848 34312
rect 56610 34296 57230 34718
rect 57280 34670 57846 34704
rect 57280 34348 57314 34670
rect 57651 34590 57662 34601
rect 57335 34528 57416 34575
rect 57475 34556 57662 34590
rect 57663 34528 57744 34575
rect 57382 34490 57416 34528
rect 57710 34490 57744 34528
rect 57651 34462 57662 34473
rect 57475 34428 57662 34462
rect 57812 34348 57846 34670
rect 57280 34314 57846 34348
rect 56668 34242 56686 34281
rect 56986 34253 57016 34288
rect 57042 34253 57044 34288
rect 56702 34242 56720 34247
rect 56610 34196 57230 34242
rect 57342 34228 57784 34262
rect 57280 34201 57846 34228
rect 56610 34194 57290 34196
rect 56610 34180 57348 34194
rect 56610 34168 57230 34180
rect 56610 34166 57262 34168
rect 56610 34133 57320 34166
rect 56610 34099 60480 34133
rect 56610 34063 57230 34099
rect 57280 33966 57320 34099
rect 57328 33972 57348 34092
rect 57382 34065 57416 34068
rect 57710 34065 57744 34068
rect 57280 33934 57314 33966
rect 57812 33934 57846 34099
rect 36304 32168 36370 33050
rect 37230 32204 37470 32540
rect 36754 32168 37216 32204
rect 31364 32134 37216 32168
rect 32094 32126 32252 32134
rect 31394 31998 31412 32100
rect 32786 32066 32852 32134
rect 32888 32130 32977 32134
rect 33558 32130 33635 32134
rect 32888 32066 32966 32130
rect 33558 32082 33624 32130
rect 34216 32104 34293 32134
rect 34874 32104 34951 32134
rect 35532 32130 35609 32134
rect 33546 32066 33624 32082
rect 33628 32066 33666 32104
rect 34216 32082 34424 32104
rect 34204 32066 34424 32082
rect 34438 32066 35182 32104
rect 35532 32082 35598 32130
rect 35520 32066 35598 32082
rect 35902 32066 35940 32104
rect 36190 32097 36256 32134
rect 36190 32082 36268 32097
rect 36178 32066 36268 32082
rect 31428 32032 31446 32066
rect 32202 32032 32886 32066
rect 32888 32032 33666 32066
rect 33718 32032 34424 32066
rect 34476 32032 35182 32066
rect 35234 32032 35940 32066
rect 35992 32032 36268 32066
rect 32048 31204 32166 31306
rect 32048 31184 32214 31204
rect 32094 31056 32214 31184
rect 32786 31196 32852 32032
rect 32888 31994 32966 32032
rect 33546 31994 33624 32032
rect 32900 31982 32966 31994
rect 32898 31360 32966 31982
rect 32976 31632 33004 31768
rect 32898 31202 32972 31360
rect 32982 31298 33000 31304
rect 33558 31298 33624 31994
rect 33656 31993 33658 31998
rect 34204 31994 34293 32032
rect 34862 31994 34951 32032
rect 35520 31994 35598 32032
rect 36178 31994 36268 32032
rect 33645 31982 33690 31993
rect 33656 31336 33690 31982
rect 34216 31768 34293 31994
rect 34403 31982 34459 31993
rect 34216 31336 34322 31768
rect 34342 31336 34378 31768
rect 34414 31336 34459 31982
rect 34874 31336 34951 31994
rect 35161 31982 35217 31993
rect 35172 31336 35217 31982
rect 33656 31298 33694 31336
rect 34216 31298 35228 31336
rect 35532 31298 35598 31994
rect 35919 31982 35964 31993
rect 35930 31336 35964 31982
rect 35930 31298 35968 31336
rect 36190 31298 36256 31994
rect 32978 31264 33624 31298
rect 33636 31264 34293 31298
rect 34310 31264 34951 31298
rect 34968 31264 35598 31298
rect 35610 31264 36256 31298
rect 32982 31258 33000 31264
rect 32898 31200 32966 31202
rect 33558 31200 33624 31264
rect 33656 31200 33690 31264
rect 34216 31258 34293 31264
rect 32898 31196 32977 31200
rect 33558 31196 33635 31200
rect 33656 31196 33701 31200
rect 34216 31196 34322 31258
rect 34342 31196 34378 31258
rect 34414 31196 34459 31264
rect 34874 31196 34951 31264
rect 35172 31196 35217 31264
rect 35532 31200 35598 31264
rect 35930 31200 35964 31264
rect 36190 31200 36256 31264
rect 35532 31196 35609 31200
rect 35930 31196 35975 31200
rect 36190 31196 36267 31200
rect 36304 31196 36370 32134
rect 36406 32120 36636 32128
rect 36580 32026 36636 32034
rect 36754 31902 37216 32134
rect 37230 31902 37692 32204
rect 44606 32168 44640 33696
rect 52920 32168 52954 33696
rect 74317 33341 74351 36356
rect 77063 36338 77097 36356
rect 74386 36300 77804 36338
rect 74431 33437 74465 33471
rect 75089 33437 75123 33471
rect 75747 33437 75781 33471
rect 76405 33437 76439 33471
rect 77063 33437 77097 36300
rect 77721 33437 77755 33471
rect 74399 33403 77789 33437
rect 56504 32168 56538 33322
rect 40320 32134 58060 32168
rect 44606 32066 44640 32134
rect 44708 32066 44742 32134
rect 44998 32066 45036 32104
rect 45756 32066 45794 32104
rect 46514 32066 46552 32104
rect 47272 32066 47310 32104
rect 48030 32066 48068 32104
rect 48788 32066 48826 32104
rect 49546 32066 49584 32104
rect 50304 32066 50342 32104
rect 51062 32066 51100 32104
rect 51820 32066 51858 32104
rect 52578 32066 52616 32104
rect 52818 32066 52852 32134
rect 52920 32066 52954 32134
rect 44606 32032 45036 32066
rect 45088 32032 45794 32066
rect 45846 32032 46552 32066
rect 46604 32032 47310 32066
rect 47362 32032 48068 32066
rect 48120 32032 48826 32066
rect 48878 32032 49584 32066
rect 49636 32032 50342 32066
rect 50394 32032 51100 32066
rect 51152 32032 51858 32066
rect 51910 32032 52616 32066
rect 52668 32032 52954 32066
rect 55596 32032 55626 32066
rect 36808 31818 37158 31852
rect 36618 31778 36642 31804
rect 36646 31750 36670 31776
rect 36580 31704 36606 31730
rect 32786 31162 36370 31196
rect 32786 30492 32852 31162
rect 32898 30492 32977 31162
rect 33558 30492 33635 31162
rect 33656 30492 33701 31162
rect 34216 30794 34322 31162
rect 34342 30794 34378 31162
rect 34216 30492 34293 30794
rect 34414 30492 34459 31162
rect 34874 30492 34951 31162
rect 35172 30492 35217 31162
rect 35532 30492 35609 31162
rect 35930 30492 35975 31162
rect 36190 30526 36267 31162
rect 36190 30492 36276 30526
rect 36304 30492 36370 31162
rect 36618 31126 36630 31480
rect 36646 31126 36658 31480
rect 36808 31338 36842 31818
rect 37000 31750 37038 31788
rect 36966 31716 37038 31750
rect 36911 31666 36956 31677
rect 36999 31666 37044 31677
rect 36922 31490 36956 31666
rect 37010 31490 37044 31666
rect 37000 31440 37038 31478
rect 36966 31406 37038 31440
rect 37124 31338 37158 31818
rect 36808 31304 37158 31338
rect 37284 31818 37634 31852
rect 37284 31338 37318 31818
rect 37446 31784 37484 31788
rect 37446 31766 37510 31784
rect 37434 31716 37510 31766
rect 37434 31700 37492 31716
rect 37412 31678 37432 31682
rect 37412 31677 37438 31678
rect 37387 31666 37438 31677
rect 37398 31490 37438 31666
rect 37412 31478 37438 31490
rect 37440 31478 37480 31700
rect 37486 31677 37514 31682
rect 37486 31490 37520 31677
rect 37412 31474 37432 31478
rect 37440 31474 37484 31478
rect 37486 31474 37514 31490
rect 37440 31456 37510 31474
rect 37434 31406 37510 31456
rect 37434 31390 37492 31406
rect 37600 31338 37634 31818
rect 37284 31304 37634 31338
rect 36646 31070 36686 31126
rect 32786 30458 36370 30492
rect 31500 29072 31526 29078
rect 31528 29072 31554 29106
rect 31908 29014 32370 29652
rect 31966 28930 32316 28964
rect 31966 28450 32000 28930
rect 32086 28896 32178 28900
rect 32086 28862 32192 28896
rect 32124 28828 32192 28862
rect 32128 28790 32174 28828
rect 32069 28778 32125 28789
rect 32080 28602 32125 28778
rect 32140 28778 32174 28790
rect 32186 28778 32213 28789
rect 32140 28602 32213 28778
rect 32140 28590 32174 28602
rect 32086 28586 32178 28590
rect 32086 28552 32192 28586
rect 32124 28518 32192 28552
rect 32128 28502 32174 28518
rect 32282 28450 32316 28930
rect 31232 28424 31303 28449
rect 31966 28424 32316 28450
rect 32786 28542 32852 30458
rect 32898 30428 32977 30458
rect 33558 30428 33635 30458
rect 33656 30428 33701 30458
rect 34216 30428 34293 30458
rect 34414 30428 34459 30458
rect 34874 30428 34951 30458
rect 35172 30428 35217 30458
rect 35532 30428 35609 30458
rect 35930 30428 35975 30458
rect 36190 30428 36267 30458
rect 32898 30356 36267 30428
rect 32898 30100 32977 30356
rect 33558 30100 33635 30356
rect 33656 30100 33701 30356
rect 32898 29962 32966 30100
rect 33558 29962 33624 30100
rect 33656 29962 33690 30100
rect 34216 30038 34293 30356
rect 32898 29606 32977 29962
rect 32898 29016 33004 29606
rect 32898 28946 32977 29016
rect 32978 28978 32994 28994
rect 32994 28974 33000 28978
rect 32898 28938 32978 28946
rect 32994 28938 33006 28974
rect 32898 28922 32994 28938
rect 32898 28694 32977 28922
rect 33558 28694 33635 29962
rect 32898 28542 32934 28694
rect 32944 28542 32945 28694
rect 33558 28682 33603 28694
rect 33656 28682 33701 29962
rect 34216 29930 34304 30038
rect 33912 29606 34304 29930
rect 33912 29422 34322 29606
rect 34216 28938 34322 29422
rect 34342 28938 34378 29606
rect 34216 28694 34293 28938
rect 34216 28682 34261 28694
rect 34414 28682 34459 30356
rect 34874 28694 34951 30356
rect 34874 28682 34919 28694
rect 35172 28682 35217 30356
rect 35532 30288 35609 30356
rect 35930 30288 35975 30356
rect 35532 30030 35598 30288
rect 35532 29964 35620 30030
rect 35384 29456 35706 29964
rect 35930 29962 35964 30288
rect 35990 30272 35998 30288
rect 36190 30262 36267 30356
rect 36190 29962 36256 30262
rect 35532 29376 35620 29456
rect 35532 28694 35609 29376
rect 35532 28682 35577 28694
rect 35930 28682 35975 29962
rect 36190 28694 36267 29962
rect 36190 28682 36235 28694
rect 32956 28644 33603 28682
rect 33614 28644 34261 28682
rect 34272 28644 34919 28682
rect 34930 28644 35577 28682
rect 35588 28644 36235 28682
rect 32994 28610 33603 28644
rect 33652 28621 34261 28644
rect 33645 28610 34261 28621
rect 34310 28610 34919 28644
rect 34968 28610 35577 28644
rect 35626 28610 36235 28644
rect 33558 28542 33603 28610
rect 33656 28542 33701 28610
rect 34216 28542 34261 28610
rect 34414 28542 34459 28610
rect 34874 28542 34919 28610
rect 35172 28542 35217 28610
rect 35532 28542 35577 28610
rect 35930 28542 35975 28610
rect 36190 28542 36235 28610
rect 36304 28542 36370 30458
rect 36754 29248 37216 29886
rect 37230 29248 37692 29886
rect 36808 29164 37158 29198
rect 36580 29050 36606 29076
rect 36580 28994 36662 29020
rect 36808 28684 36842 29164
rect 36948 29136 36954 29138
rect 37018 29136 37028 29138
rect 36928 29096 37038 29134
rect 36966 29066 37038 29096
rect 36948 29064 37038 29066
rect 36966 29062 37038 29064
rect 36911 29012 36967 29023
rect 36999 29012 37055 29023
rect 36922 28836 36967 29012
rect 37010 28836 37055 29012
rect 36928 28786 37038 28824
rect 36966 28752 37038 28786
rect 37124 28684 37158 29164
rect 36808 28650 37158 28684
rect 37284 29164 37634 29198
rect 37284 28684 37318 29164
rect 37424 29136 37430 29138
rect 37404 29130 37484 29134
rect 37404 29096 37510 29130
rect 37434 29066 37510 29096
rect 37424 29064 37510 29066
rect 37434 29062 37510 29064
rect 37434 29046 37492 29062
rect 37392 29023 37438 29024
rect 37387 29020 37438 29023
rect 37384 28962 37438 29020
rect 37440 29020 37480 29046
rect 37492 29020 37531 29023
rect 37440 28962 37531 29020
rect 37398 28836 37434 28962
rect 37444 28824 37480 28962
rect 37486 28836 37531 28962
rect 37404 28820 37484 28824
rect 37404 28786 37510 28820
rect 37434 28752 37510 28786
rect 37434 28736 37492 28752
rect 37600 28684 37634 29164
rect 37284 28650 37634 28684
rect 32786 28508 36370 28542
rect 32786 28424 32820 28508
rect 32898 28424 32934 28508
rect 32944 28424 32945 28508
rect 33558 28424 33603 28508
rect 33656 28424 33701 28508
rect 34216 28424 34261 28508
rect 34414 28424 34459 28508
rect 34874 28424 34919 28508
rect 35172 28424 35217 28508
rect 35532 28424 35577 28508
rect 35930 28424 35975 28508
rect 36190 28424 36235 28508
rect 36304 28424 36338 28508
rect 43510 28424 43544 31982
rect 44606 30274 44640 32032
rect 44708 31732 44742 32032
rect 44780 31994 44781 31995
rect 52779 31994 52780 31995
rect 44779 31993 44780 31994
rect 52780 31993 52781 31994
rect 45015 31982 45060 31993
rect 45773 31982 45818 31993
rect 46531 31982 46576 31993
rect 47289 31982 47334 31993
rect 48047 31982 48092 31993
rect 48805 31982 48850 31993
rect 49563 31982 49608 31993
rect 50321 31982 50366 31993
rect 51079 31982 51124 31993
rect 51837 31982 51882 31993
rect 52595 31982 52640 31993
rect 45014 31716 45015 31717
rect 45013 31715 45014 31716
rect 45026 31704 45060 31982
rect 45071 31716 45072 31717
rect 45772 31716 45773 31717
rect 45072 31715 45073 31716
rect 45771 31715 45772 31716
rect 45784 31704 45818 31982
rect 45829 31716 45830 31717
rect 46530 31716 46531 31717
rect 45830 31715 45831 31716
rect 46529 31715 46530 31716
rect 46542 31704 46576 31982
rect 46587 31716 46588 31717
rect 47288 31716 47289 31717
rect 46588 31715 46589 31716
rect 47287 31715 47288 31716
rect 47300 31704 47334 31982
rect 47345 31716 47346 31717
rect 48046 31716 48047 31717
rect 47346 31715 47347 31716
rect 48045 31715 48046 31716
rect 48058 31704 48092 31982
rect 48742 31796 48810 31804
rect 48770 31768 48810 31776
rect 48103 31716 48104 31717
rect 48804 31716 48805 31717
rect 48104 31715 48105 31716
rect 48803 31715 48804 31716
rect 48816 31704 48850 31982
rect 48856 31796 48922 31804
rect 48856 31768 48894 31776
rect 48861 31716 48862 31717
rect 49562 31716 49563 31717
rect 48862 31715 48863 31716
rect 49561 31715 49562 31716
rect 49574 31704 49608 31982
rect 50256 31796 50326 31816
rect 50284 31768 50326 31788
rect 49619 31716 49620 31717
rect 50320 31716 50321 31717
rect 49620 31715 49621 31716
rect 50319 31715 50320 31716
rect 50332 31704 50366 31982
rect 50372 31796 50436 31816
rect 50372 31768 50408 31788
rect 50377 31716 50378 31717
rect 51078 31716 51079 31717
rect 50378 31715 50379 31716
rect 51077 31715 51078 31716
rect 51090 31704 51124 31982
rect 51135 31716 51136 31717
rect 51836 31716 51837 31717
rect 51136 31715 51137 31716
rect 51835 31715 51836 31716
rect 51848 31704 51882 31982
rect 51893 31716 51894 31717
rect 52594 31716 52595 31717
rect 51894 31715 51895 31716
rect 52593 31715 52594 31716
rect 52606 31704 52640 31982
rect 52818 31732 52852 32032
rect 52651 31716 52652 31717
rect 52652 31715 52653 31716
rect 52768 31704 52779 31715
rect 44670 31642 44742 31680
rect 44792 31670 52779 31704
rect 45013 31658 45014 31659
rect 45014 31657 45015 31658
rect 44708 31074 44742 31642
rect 45014 31058 45015 31059
rect 45013 31057 45014 31058
rect 45026 31046 45060 31670
rect 45072 31658 45073 31659
rect 45771 31658 45772 31659
rect 45071 31657 45072 31658
rect 45772 31657 45773 31658
rect 45784 31090 45818 31670
rect 45830 31658 45831 31659
rect 46529 31658 46530 31659
rect 45829 31657 45830 31658
rect 46530 31657 46531 31658
rect 45740 31084 45860 31090
rect 45071 31058 45072 31059
rect 45772 31058 45773 31059
rect 45072 31057 45073 31058
rect 45771 31057 45772 31058
rect 45784 31046 45818 31084
rect 45829 31058 45830 31059
rect 46530 31058 46531 31059
rect 45830 31057 45831 31058
rect 46529 31057 46530 31058
rect 46542 31046 46576 31670
rect 46588 31658 46589 31659
rect 47287 31658 47288 31659
rect 46587 31657 46588 31658
rect 47288 31657 47289 31658
rect 46587 31058 46588 31059
rect 47288 31058 47289 31059
rect 46588 31057 46589 31058
rect 47287 31057 47288 31058
rect 47300 31046 47334 31670
rect 47346 31658 47347 31659
rect 48045 31658 48046 31659
rect 47345 31657 47346 31658
rect 48046 31657 48047 31658
rect 47345 31058 47346 31059
rect 48046 31058 48047 31059
rect 47346 31057 47347 31058
rect 48045 31057 48046 31058
rect 48058 31046 48092 31670
rect 48104 31658 48105 31659
rect 48803 31658 48804 31659
rect 48103 31657 48104 31658
rect 48804 31657 48805 31658
rect 48103 31058 48104 31059
rect 48804 31058 48805 31059
rect 48104 31057 48105 31058
rect 48803 31057 48804 31058
rect 48816 31046 48850 31670
rect 48862 31658 48863 31659
rect 49561 31658 49562 31659
rect 48861 31657 48862 31658
rect 49562 31657 49563 31658
rect 48861 31058 48862 31059
rect 49562 31058 49563 31059
rect 48862 31057 48863 31058
rect 49561 31057 49562 31058
rect 49574 31046 49608 31670
rect 49620 31658 49621 31659
rect 50319 31658 50320 31659
rect 49619 31657 49620 31658
rect 50320 31657 50321 31658
rect 49619 31058 49620 31059
rect 50320 31058 50321 31059
rect 49620 31057 49621 31058
rect 50319 31057 50320 31058
rect 50332 31046 50366 31670
rect 50378 31658 50379 31659
rect 51077 31658 51078 31659
rect 50377 31657 50378 31658
rect 51078 31657 51079 31658
rect 50377 31058 50378 31059
rect 51078 31058 51079 31059
rect 50378 31057 50379 31058
rect 51077 31057 51078 31058
rect 51090 31046 51124 31670
rect 51136 31658 51137 31659
rect 51835 31658 51836 31659
rect 51135 31657 51136 31658
rect 51836 31657 51837 31658
rect 51135 31058 51136 31059
rect 51836 31058 51837 31059
rect 51136 31057 51137 31058
rect 51835 31057 51836 31058
rect 51848 31046 51882 31670
rect 51894 31658 51895 31659
rect 52593 31658 52594 31659
rect 51893 31657 51894 31658
rect 52594 31657 52595 31658
rect 51893 31058 51894 31059
rect 52594 31058 52595 31059
rect 51894 31057 51895 31058
rect 52593 31057 52594 31058
rect 52606 31046 52640 31670
rect 52652 31658 52653 31659
rect 52651 31657 52652 31658
rect 52780 31642 52852 31680
rect 52818 31074 52852 31642
rect 52651 31058 52652 31059
rect 52652 31057 52653 31058
rect 52768 31046 52779 31057
rect 44670 30984 44742 31022
rect 44792 31012 52779 31046
rect 45013 31000 45014 31001
rect 45014 30999 45015 31000
rect 44708 30416 44742 30984
rect 45014 30400 45015 30401
rect 45013 30399 45014 30400
rect 45026 30388 45060 31012
rect 45072 31000 45073 31001
rect 45771 31000 45772 31001
rect 45071 30999 45072 31000
rect 45772 30999 45773 31000
rect 45071 30400 45072 30401
rect 45772 30400 45773 30401
rect 45072 30399 45073 30400
rect 45771 30399 45772 30400
rect 45784 30388 45818 31012
rect 45830 31000 45831 31001
rect 46529 31000 46530 31001
rect 45829 30999 45830 31000
rect 46530 30999 46531 31000
rect 45829 30400 45830 30401
rect 46530 30400 46531 30401
rect 45830 30399 45831 30400
rect 46529 30399 46530 30400
rect 46542 30388 46576 31012
rect 46588 31000 46589 31001
rect 47287 31000 47288 31001
rect 46587 30999 46588 31000
rect 47288 30999 47289 31000
rect 46587 30400 46588 30401
rect 47288 30400 47289 30401
rect 46588 30399 46589 30400
rect 47287 30399 47288 30400
rect 47300 30388 47334 31012
rect 47346 31000 47347 31001
rect 48045 31000 48046 31001
rect 47345 30999 47346 31000
rect 48046 30999 48047 31000
rect 47345 30400 47346 30401
rect 48046 30400 48047 30401
rect 47346 30399 47347 30400
rect 48045 30399 48046 30400
rect 48058 30388 48092 31012
rect 48104 31000 48105 31001
rect 48803 31000 48804 31001
rect 48103 30999 48104 31000
rect 48804 30999 48805 31000
rect 48708 30420 48718 30486
rect 48736 30448 48746 30486
rect 48103 30400 48104 30401
rect 48804 30400 48805 30401
rect 48104 30399 48105 30400
rect 48803 30399 48804 30400
rect 48816 30388 48850 31012
rect 48862 31000 48863 31001
rect 49561 31000 49562 31001
rect 48861 30999 48862 31000
rect 49562 30999 49563 31000
rect 48861 30400 48862 30401
rect 49562 30400 49563 30401
rect 48862 30399 48863 30400
rect 49561 30399 49562 30400
rect 49574 30388 49608 31012
rect 49620 31000 49621 31001
rect 50319 31000 50320 31001
rect 49619 30999 49620 31000
rect 50320 30999 50321 31000
rect 49619 30400 49620 30401
rect 49620 30399 49621 30400
rect 50284 30398 50326 30422
rect 50256 30388 50326 30394
rect 50332 30388 50366 31012
rect 50378 31000 50379 31001
rect 51077 31000 51078 31001
rect 50377 30999 50378 31000
rect 51078 30999 51079 31000
rect 50372 30398 50408 30422
rect 51078 30400 51079 30401
rect 51077 30399 51078 30400
rect 50372 30388 50436 30394
rect 51090 30388 51124 31012
rect 51136 31000 51137 31001
rect 51835 31000 51836 31001
rect 51135 30999 51136 31000
rect 51836 30999 51837 31000
rect 51135 30400 51136 30401
rect 51836 30400 51837 30401
rect 51136 30399 51137 30400
rect 51835 30399 51836 30400
rect 51848 30388 51882 31012
rect 51894 31000 51895 31001
rect 52593 31000 52594 31001
rect 51893 30999 51894 31000
rect 52594 30999 52595 31000
rect 51893 30400 51894 30401
rect 52594 30400 52595 30401
rect 51894 30399 51895 30400
rect 52593 30399 52594 30400
rect 52606 30388 52640 31012
rect 52652 31000 52653 31001
rect 52651 30999 52652 31000
rect 52780 30984 52852 31022
rect 52818 30416 52852 30984
rect 52651 30400 52652 30401
rect 52652 30399 52653 30400
rect 52768 30388 52779 30399
rect 44792 30354 52779 30388
rect 45026 30274 45060 30354
rect 45784 30274 45818 30354
rect 46542 30274 46576 30354
rect 47300 30274 47334 30354
rect 48058 30274 48092 30354
rect 48816 30274 48850 30354
rect 49574 30274 49608 30354
rect 50332 30274 50366 30354
rect 51090 30274 51124 30354
rect 51848 30274 51882 30354
rect 52606 30274 52640 30354
rect 52920 30274 52954 32032
rect 55630 31998 55660 32100
rect 56504 32066 56538 32134
rect 56582 32086 56600 32100
rect 56554 32066 56600 32072
rect 56606 32066 56640 32134
rect 57126 32100 57164 32104
rect 57884 32100 57922 32104
rect 56646 32086 57166 32100
rect 57176 32086 57924 32100
rect 57126 32072 57164 32086
rect 57884 32072 57922 32086
rect 56646 32066 57164 32072
rect 56504 32032 57164 32066
rect 57204 32058 57922 32072
rect 57216 32032 57922 32058
rect 55656 30532 55672 31050
rect 55694 30570 55710 31012
rect 44606 30240 52954 30274
rect 48058 28757 48092 30240
rect 48692 29906 48718 29936
rect 48720 29934 48746 29936
rect 48782 29934 48806 29936
rect 48810 29906 48834 29936
rect 56504 29900 56538 32032
rect 56606 32016 56640 32032
rect 56678 31994 57142 32000
rect 57200 31994 57900 32000
rect 58026 31988 58060 32134
rect 56568 31926 56640 31964
rect 56690 31954 58060 31988
rect 57141 31942 57142 31943
rect 57142 31941 57143 31942
rect 56606 31358 56640 31926
rect 57142 31342 57143 31343
rect 57141 31341 57142 31342
rect 57154 31330 57188 31954
rect 57200 31942 57201 31943
rect 57899 31942 57900 31943
rect 57199 31941 57200 31942
rect 57900 31941 57901 31942
rect 57199 31342 57200 31343
rect 57900 31342 57901 31343
rect 57200 31341 57201 31342
rect 57899 31341 57900 31342
rect 57912 31330 57946 31954
rect 58026 31330 58060 31954
rect 56568 31268 56640 31306
rect 56690 31296 58060 31330
rect 57141 31284 57142 31285
rect 57142 31283 57143 31284
rect 56606 30700 56640 31268
rect 57142 30684 57143 30685
rect 57141 30683 57142 30684
rect 57154 30672 57188 31296
rect 57200 31284 57201 31285
rect 57899 31284 57900 31285
rect 57199 31283 57200 31284
rect 57900 31283 57901 31284
rect 57199 30684 57200 30685
rect 57900 30684 57901 30685
rect 57200 30683 57201 30684
rect 57899 30683 57900 30684
rect 57912 30672 57946 31296
rect 58026 30672 58060 31296
rect 56568 30610 56640 30648
rect 56690 30638 58060 30672
rect 57141 30626 57142 30627
rect 57142 30625 57143 30626
rect 56606 30042 56640 30610
rect 57142 30026 57143 30027
rect 57141 30025 57142 30026
rect 57154 30014 57188 30638
rect 57200 30626 57201 30627
rect 57899 30626 57900 30627
rect 57199 30625 57200 30626
rect 57900 30625 57901 30626
rect 57199 30026 57200 30027
rect 57900 30026 57901 30027
rect 57200 30025 57201 30026
rect 57899 30025 57900 30026
rect 57912 30014 57946 30638
rect 58026 30014 58060 30638
rect 56690 29996 58060 30014
rect 74303 31839 74351 33341
rect 74431 33351 74465 33403
rect 75089 33382 75123 33403
rect 75747 33382 75781 33403
rect 76405 33382 76439 33403
rect 77063 33382 77097 33403
rect 77721 33382 77755 33403
rect 75047 33351 75123 33382
rect 75705 33351 75781 33382
rect 76363 33351 76439 33382
rect 77021 33351 77097 33382
rect 74431 33254 74477 33351
rect 75047 33335 75135 33351
rect 75705 33335 75793 33351
rect 76363 33335 76451 33351
rect 77021 33335 77109 33351
rect 77679 33335 77755 33382
rect 77835 33341 77869 36356
rect 79388 36384 79422 38226
rect 79490 38164 79536 38316
rect 80088 38272 80114 39392
rect 80116 38272 80142 39364
rect 80160 38316 80226 39928
rect 80818 38316 80884 39928
rect 80160 38304 80194 38316
rect 80818 38304 80852 38316
rect 80148 38266 80198 38304
rect 80252 38272 80270 38288
rect 80806 38266 80856 38304
rect 81408 38272 81424 39374
rect 81436 38272 81452 39346
rect 81476 38316 81542 39928
rect 82134 38316 82200 39928
rect 82232 38570 82238 39972
rect 82260 38542 82266 39972
rect 82781 39928 82812 39939
rect 82824 39928 82858 40080
rect 81476 38304 81510 38316
rect 82134 38304 82168 38316
rect 81464 38266 81514 38304
rect 82122 38266 82172 38304
rect 82716 38272 82740 39376
rect 82744 38272 82768 39348
rect 82792 38316 82858 39928
rect 82906 40018 82924 40080
rect 82938 40018 82972 40320
rect 82792 38304 82826 38316
rect 82780 38266 82830 38304
rect 79596 38232 80198 38266
rect 80254 38232 80856 38266
rect 80912 38232 81514 38266
rect 81570 38232 82172 38266
rect 82228 38232 82830 38266
rect 80148 38216 80194 38232
rect 80806 38216 80852 38232
rect 81464 38216 81510 38232
rect 82122 38216 82168 38232
rect 82780 38216 82826 38232
rect 82906 38226 82972 40018
rect 83526 38954 83646 38974
rect 83832 38956 84072 39508
rect 83832 38954 84122 38956
rect 83520 38926 83674 38946
rect 83832 38928 84072 38954
rect 83832 38926 84150 38928
rect 83832 38870 84072 38926
rect 80160 38164 80194 38216
rect 79490 38130 82838 38164
rect 80160 36384 80194 38130
rect 82128 36384 82150 36574
rect 82906 36384 82940 38226
rect 90894 36898 90896 36948
rect 90922 36898 90924 36976
rect 90342 36658 90980 36898
rect 96108 36854 96110 36932
rect 96136 36854 96138 36904
rect 96052 36614 96690 36854
rect 79388 36356 82940 36384
rect 79082 35914 79084 35962
rect 79054 35886 79084 35906
rect 79388 33346 79422 36356
rect 80160 36328 80194 36356
rect 82128 36328 82150 36356
rect 79460 36300 82878 36328
rect 79502 33442 79536 33476
rect 80160 33442 80194 36300
rect 82128 35906 82150 36300
rect 80852 33644 80858 34718
rect 80852 33476 80884 33644
rect 80818 33442 80884 33476
rect 80908 33442 80912 33672
rect 81476 33442 81510 33476
rect 82070 33442 82096 33636
rect 82128 33608 82152 34718
rect 82098 33476 82152 33608
rect 82098 33442 82168 33476
rect 82792 33442 82826 33476
rect 79470 33408 82860 33442
rect 74479 33301 75135 33335
rect 75137 33301 75793 33335
rect 75795 33301 76451 33335
rect 76453 33301 77109 33335
rect 77111 33301 77755 33335
rect 75055 33295 75059 33301
rect 75083 33267 75087 33301
rect 75089 33254 75135 33301
rect 75747 33254 75793 33301
rect 76371 33295 76375 33301
rect 76399 33267 76403 33301
rect 76405 33254 76451 33301
rect 77063 33254 77109 33301
rect 77687 33295 77691 33301
rect 77715 33267 77719 33301
rect 74431 33242 74465 33254
rect 75064 33242 75077 33253
rect 75089 33242 75123 33254
rect 75722 33242 75735 33253
rect 75747 33242 75781 33254
rect 76380 33242 76393 33253
rect 76405 33242 76439 33254
rect 77038 33242 77051 33253
rect 77063 33242 77097 33254
rect 77696 33242 77709 33253
rect 77721 33242 77755 33301
rect 74417 31938 74465 33242
rect 75075 31938 75123 33242
rect 75733 31938 75781 33242
rect 56674 29980 58184 29996
rect 57154 29962 57188 29980
rect 57912 29962 57946 29980
rect 58026 29962 58060 29980
rect 56640 29946 58150 29962
rect 57154 29900 57188 29946
rect 57912 29900 57946 29946
rect 58026 29900 58060 29946
rect 48298 29824 48620 29896
rect 56504 29866 60480 29900
rect 48100 29362 48738 29824
rect 48788 29736 49336 29770
rect 48788 29454 48822 29736
rect 48963 29656 49161 29667
rect 48852 29612 48962 29650
rect 48974 29622 49161 29656
rect 49162 29612 49272 29650
rect 48890 29578 48962 29612
rect 48963 29568 49161 29579
rect 49200 29578 49272 29612
rect 48974 29534 49161 29568
rect 49302 29454 49336 29736
rect 48788 29420 49336 29454
rect 50298 29414 50316 29614
rect 50326 29386 50344 29642
rect 44575 28424 53013 28757
rect 31232 28390 31321 28424
rect 31370 28401 57958 28424
rect 58026 28401 58060 29866
rect 31370 28390 58060 28401
rect 31232 27282 31303 28390
rect 31382 27422 31416 28390
rect 32140 28360 32174 28390
rect 32786 28360 32820 28390
rect 32898 28360 32934 28390
rect 32944 28360 32945 28390
rect 33558 28360 33603 28390
rect 33656 28360 33701 28390
rect 34216 28360 34261 28390
rect 34414 28360 34459 28390
rect 34874 28360 34919 28390
rect 35172 28360 35217 28390
rect 35532 28360 35577 28390
rect 35930 28360 35975 28390
rect 36190 28360 36235 28390
rect 36304 28360 36338 28390
rect 36688 28360 36722 28390
rect 37446 28360 37480 28390
rect 38204 28360 38238 28390
rect 38962 28360 38996 28390
rect 39720 28360 39754 28390
rect 40478 28360 40512 28390
rect 41236 28360 41270 28390
rect 41994 28360 42028 28390
rect 42752 28360 42786 28390
rect 42796 28360 42820 28386
rect 43510 28360 43544 28390
rect 44268 28360 44302 28390
rect 44575 28360 53013 28390
rect 53364 28360 53398 28390
rect 54122 28360 54156 28390
rect 54880 28360 54914 28390
rect 55638 28360 55672 28390
rect 56396 28360 56430 28390
rect 58026 28383 58060 28390
rect 31962 28322 32700 28360
rect 32786 28322 36384 28360
rect 36660 28322 36722 28360
rect 37418 28322 37480 28360
rect 38176 28322 38238 28360
rect 38934 28322 38996 28360
rect 39692 28322 39754 28360
rect 40450 28322 40512 28360
rect 41208 28322 41270 28360
rect 41966 28322 42028 28360
rect 42724 28322 53013 28360
rect 53336 28322 53398 28360
rect 54094 28322 54156 28360
rect 54852 28322 54914 28360
rect 55610 28322 55672 28360
rect 56368 28356 56430 28360
rect 56368 28328 56436 28356
rect 56362 28322 56436 28328
rect 56445 28322 58096 28383
rect 31428 28288 32174 28322
rect 32202 28288 32934 28322
rect 32140 27422 32174 28288
rect 31382 27384 31456 27422
rect 32112 27384 32174 27422
rect 32786 27384 32820 28288
rect 32898 27422 32934 28288
rect 32870 27384 32934 27422
rect 31382 27282 31416 27384
rect 31444 27350 32174 27384
rect 32186 27350 32934 27384
rect 32140 27282 32174 27350
rect 32786 27282 32820 27350
rect 32898 27282 32934 27350
rect 32944 27384 32945 28322
rect 32960 28288 33701 28322
rect 33718 28288 34459 28322
rect 34476 28288 35217 28322
rect 35234 28288 35975 28322
rect 35992 28288 36722 28322
rect 36734 28288 37480 28322
rect 37492 28288 38238 28322
rect 38250 28288 38996 28322
rect 39008 28288 39754 28322
rect 39766 28288 40512 28322
rect 40524 28288 41270 28322
rect 41282 28288 42028 28322
rect 42040 28288 42786 28322
rect 33558 27446 33603 28288
rect 33656 27446 33701 28288
rect 33558 27384 33592 27446
rect 33656 27422 33690 27446
rect 34216 27422 34261 28288
rect 34414 27422 34459 28288
rect 34874 27422 34919 28288
rect 35172 27422 35217 28288
rect 33628 27384 33690 27422
rect 34212 27384 35217 27422
rect 35532 27634 35577 28288
rect 35930 27634 35975 28288
rect 35532 27384 35566 27634
rect 35930 27422 35964 27634
rect 35990 27618 35998 27634
rect 35902 27384 35964 27422
rect 36190 27608 36235 28288
rect 36190 27384 36224 27608
rect 36304 27384 36338 28288
rect 36688 28284 36722 28288
rect 37446 28284 37480 28288
rect 38204 28284 38238 28288
rect 38962 28284 38996 28288
rect 39720 28284 39754 28288
rect 36476 28254 40154 28284
rect 36688 27422 36722 28254
rect 37446 27422 37480 28254
rect 38204 27422 38238 28254
rect 38962 27422 38996 28254
rect 39720 27422 39754 28254
rect 40478 27422 40512 28288
rect 41236 27422 41270 28288
rect 41994 27422 42028 28288
rect 42752 27422 42786 28288
rect 42796 28288 43544 28322
rect 43572 28288 44302 28322
rect 44330 28288 53398 28322
rect 53410 28288 54156 28322
rect 54168 28288 54914 28322
rect 54926 28288 55672 28322
rect 55684 28288 56436 28322
rect 56442 28288 58096 28322
rect 42796 27422 42820 28288
rect 43510 27422 43544 28288
rect 44268 27422 44302 28288
rect 44575 27422 53013 28288
rect 53364 27422 53398 28288
rect 54122 27422 54156 28288
rect 54880 27422 54914 28288
rect 55638 27422 55672 28288
rect 56362 28282 56380 28288
rect 56390 28254 56436 28288
rect 56396 27422 56430 28254
rect 36452 27384 40212 27422
rect 40450 27418 40512 27422
rect 40450 27390 40518 27418
rect 40444 27384 40518 27390
rect 40528 27384 40546 27390
rect 41208 27384 41270 27422
rect 41966 27418 42028 27422
rect 41966 27390 42034 27418
rect 41960 27384 42034 27390
rect 42044 27384 42062 27390
rect 42724 27384 53013 27422
rect 53336 27384 53398 27422
rect 54094 27384 54156 27422
rect 54852 27384 54914 27422
rect 55610 27384 55672 27422
rect 56368 27384 56430 27422
rect 56445 27384 58096 28288
rect 32944 27350 33690 27384
rect 33702 27350 34459 27384
rect 34476 27350 35217 27384
rect 35234 27350 35964 27384
rect 35976 27350 36722 27384
rect 36750 27350 37486 27384
rect 32944 27282 32945 27350
rect 33558 27282 33592 27350
rect 33656 27282 33690 27350
rect 34216 27282 34261 27350
rect 34414 27282 34459 27350
rect 34874 27282 34919 27350
rect 35172 27282 35217 27350
rect 35532 27282 35566 27350
rect 35930 27282 35964 27350
rect 36190 27282 36224 27350
rect 36304 27282 36338 27350
rect 36688 27282 36722 27350
rect 37412 27344 37430 27350
rect 37440 27316 37486 27350
rect 37496 27350 38238 27384
rect 38266 27350 39002 27384
rect 37496 27344 37514 27350
rect 37446 27282 37480 27316
rect 38204 27282 38238 27350
rect 38928 27344 38946 27350
rect 38956 27316 39002 27350
rect 39012 27350 39754 27384
rect 39782 27350 40518 27384
rect 40524 27350 41270 27384
rect 41282 27350 42034 27384
rect 42040 27350 42786 27384
rect 39012 27344 39030 27350
rect 38962 27282 38996 27316
rect 39720 27282 39754 27350
rect 40444 27344 40462 27350
rect 40472 27316 40518 27350
rect 40528 27344 40546 27350
rect 40478 27282 40512 27316
rect 41236 27282 41270 27350
rect 41960 27344 41978 27350
rect 41988 27316 42034 27350
rect 42044 27344 42062 27350
rect 41994 27282 42028 27316
rect 42752 27282 42786 27350
rect 42796 27350 43550 27384
rect 42796 27282 42820 27350
rect 43476 27344 43494 27350
rect 43504 27316 43550 27350
rect 43560 27350 44302 27384
rect 44330 27350 53398 27384
rect 53410 27350 54156 27384
rect 54168 27350 54914 27384
rect 54926 27350 55672 27384
rect 55684 27350 56430 27384
rect 56442 27350 58096 27384
rect 43560 27344 43578 27350
rect 43510 27282 43544 27316
rect 44268 27282 44302 27350
rect 44575 27282 53013 27350
rect 53364 27282 53398 27350
rect 54122 27282 54156 27350
rect 54880 27282 54914 27350
rect 55638 27282 55672 27350
rect 56396 27282 56430 27350
rect 56445 27282 58096 27350
rect 31232 27248 31321 27282
rect 31364 27248 58096 27282
rect 31232 27004 31303 27248
rect 31164 26762 31202 26948
rect 31220 26762 31303 27004
rect 27817 26435 31187 26469
rect 9866 21415 14220 21480
rect 16668 21415 18286 21510
rect 9866 20702 18286 21415
rect 19470 20752 19526 20764
rect 20714 20752 20770 20764
rect 19470 20702 19526 20708
rect 9866 20668 20160 20702
rect 20714 20696 20770 20708
rect 21312 20668 27246 22570
rect 9866 20654 18286 20668
rect 9866 20652 18452 20654
rect -14496 20316 -14490 20458
rect -14502 20294 -14490 20316
rect -1808 20310 -1508 20329
rect -156 20310 1344 20329
rect 2912 20323 4620 20329
rect 4630 20323 4664 20582
rect 4744 20323 4778 20582
rect 4982 20368 5038 20385
rect 6239 20351 6273 20582
rect 4789 20335 4790 20336
rect 4790 20334 4791 20335
rect 4908 20323 5038 20329
rect 6180 20323 6191 20334
rect 2912 20312 6191 20323
rect -14506 20268 -14490 20294
rect 4596 20289 6191 20312
rect -14506 20238 -14480 20268
rect -1564 20184 -100 20200
rect -14506 20134 -14480 20162
rect -14506 20106 -14484 20134
rect -14502 20098 -14484 20106
rect -17612 19974 -16148 19990
rect -18840 19845 -18784 19862
rect -18438 19845 -17556 19862
rect -16204 19845 -15904 19862
rect -18840 19789 -18784 19806
rect -14496 19640 -14484 20098
rect -18508 19442 -15685 19592
rect -18508 19408 -10310 19442
rect -18508 18569 -15685 19408
rect -14510 19402 -14440 19404
rect -14454 19346 -14440 19348
rect -14372 18794 -14000 18822
rect -14410 18756 -13962 18784
rect -20160 18535 -15685 18569
rect -18508 18385 -15685 18535
rect -20084 17662 -20082 17804
rect -20094 17640 -20082 17662
rect -20098 17614 -20082 17640
rect -20098 17584 -20072 17614
rect -19380 17514 -19348 17584
rect -20098 17480 -20072 17508
rect -19346 17480 -19314 17618
rect -20098 17452 -20076 17480
rect -20094 17444 -20076 17452
rect -20084 16986 -20076 17444
rect -18472 16902 -18438 18385
rect -17996 18154 -16594 18168
rect -1991 17303 -1957 20160
rect 1534 20132 2100 20166
rect 1534 19810 1568 20132
rect 2066 20068 2100 20132
rect 2150 20068 2770 20184
rect 1718 20052 1916 20063
rect 1589 19990 1717 20037
rect 1729 20018 1916 20052
rect 2002 20037 2770 20068
rect 1917 19990 2770 20037
rect 1636 19952 1717 19990
rect 1964 19952 2770 19990
rect 1718 19924 1916 19935
rect 1974 19926 2770 19952
rect 1729 19890 1916 19924
rect 2002 19856 2770 19926
rect 2066 19810 2100 19856
rect 1534 19776 2100 19810
rect 2150 19762 2770 19856
rect 4630 19665 4664 20289
rect 4744 19665 4778 20289
rect 4790 20277 4791 20278
rect 4789 20276 4790 20277
rect 6192 20261 6273 20308
rect 4982 19752 5038 19754
rect 4982 19696 5038 19698
rect 6239 19693 6273 20261
rect 4789 19677 4790 19678
rect 4790 19676 4791 19677
rect 6180 19665 6191 19676
rect 4596 19631 6191 19665
rect 4630 19456 4664 19631
rect 4744 19617 4778 19631
rect 4790 19619 4791 19620
rect 4789 19618 4790 19619
rect 6192 19605 6320 19650
rect 6191 19604 6192 19605
rect 4766 19590 5038 19592
rect 4794 19562 5038 19564
rect 4982 19558 5038 19562
rect 6239 19558 6273 19603
rect 6341 19558 6375 20582
rect 9866 20208 18286 20652
rect 4806 19524 6375 19558
rect 6239 19456 6273 19524
rect 6341 19456 6375 19524
rect 9879 19558 9913 20208
rect 9981 19977 10015 20208
rect 10848 19961 10849 19962
rect 10847 19960 10848 19961
rect 10508 19949 10854 19955
rect 10860 19949 10894 20208
rect 13918 20048 13952 20208
rect 10905 19961 10906 19962
rect 10906 19960 10907 19961
rect 10900 19949 11190 19955
rect 13342 19949 13560 19960
rect 13884 19955 13890 20048
rect 13906 19961 13907 19962
rect 13905 19960 13906 19961
rect 13912 19955 13952 20048
rect 13918 19949 13952 19955
rect 14032 19949 14066 20208
rect 9934 19887 10015 19934
rect 10074 19915 14066 19949
rect 14910 19936 16410 19955
rect 16704 19949 16738 20208
rect 16806 20072 16840 20208
rect 18109 20057 18143 20208
rect 18062 20056 18143 20057
rect 18062 20044 18159 20056
rect 16759 19982 16840 20029
rect 16899 20010 18159 20044
rect 17762 19998 18159 20010
rect 17762 19992 18143 19998
rect 16806 19962 16840 19982
rect 18103 19977 18143 19992
rect 18103 19966 18118 19977
rect 18103 19965 18149 19966
rect 16670 19915 16738 19949
rect 16759 19961 16840 19962
rect 16759 19949 16887 19961
rect 18050 19955 18061 19960
rect 17762 19949 18062 19955
rect 16759 19938 18062 19949
rect 18211 19938 18245 20208
rect 20714 20092 20770 20106
rect 20714 20036 20770 20050
rect 19470 19992 19526 19994
rect 16759 19937 19526 19938
rect 16759 19936 18103 19937
rect 18149 19936 19526 19937
rect 16759 19915 18061 19936
rect 10847 19903 10848 19904
rect 10848 19902 10849 19903
rect 9981 19558 10015 19887
rect 10860 19617 10894 19915
rect 13918 19909 13952 19915
rect 10906 19903 10907 19904
rect 10905 19902 10906 19903
rect 13884 19826 13890 19909
rect 13905 19903 13906 19904
rect 13906 19902 13907 19903
rect 13912 19826 13952 19909
rect 13918 19810 13952 19826
rect 14032 19810 14066 19915
rect 16704 19826 16738 19915
rect 16790 19903 16887 19915
rect 16354 19810 16800 19826
rect 13484 19694 14104 19810
rect 14154 19758 14720 19792
rect 14154 19694 14188 19758
rect 13484 19663 14252 19694
rect 14525 19678 14536 19689
rect 10061 19605 10062 19606
rect 13484 19605 14290 19663
rect 14349 19644 14536 19678
rect 14537 19616 14618 19663
rect 10062 19604 10063 19605
rect 10832 19558 10879 19605
rect 13342 19578 14290 19605
rect 14584 19578 14618 19616
rect 13342 19558 14280 19578
rect 9879 19524 10879 19558
rect 10922 19552 14280 19558
rect 10922 19524 14252 19552
rect 14525 19550 14536 19561
rect 9879 19456 9913 19524
rect 9981 19456 10015 19524
rect 13484 19482 14252 19524
rect 14349 19516 14536 19550
rect 13484 19456 14104 19482
rect 4630 19422 14104 19456
rect 2010 19210 2458 19422
rect 2102 19200 2234 19210
rect -1916 19088 6300 19099
rect -1905 19076 6289 19088
rect -1916 19065 6300 19076
rect -1889 19019 -1855 19065
rect -980 19007 -524 19026
rect 6239 19019 6273 19065
rect -1796 18961 6180 19007
rect -1796 18951 6191 18961
rect -1889 18355 -1855 18945
rect -942 18936 -486 18951
rect 6239 18802 6273 18945
rect 6341 18802 6375 19422
rect 9879 18802 9913 19422
rect 13484 19388 14104 19422
rect 14154 19436 14188 19482
rect 14686 19436 14720 19758
rect 14154 19402 14720 19436
rect 11134 19322 11788 19324
rect 16704 19272 16738 19810
rect 16806 19414 16840 19903
rect 18062 19887 18143 19934
rect 18109 19399 18143 19887
rect 18062 19398 18143 19399
rect 18062 19386 18159 19398
rect 16899 19355 18159 19386
rect 16899 19352 18174 19355
rect 18062 19340 18174 19352
rect 16766 19272 18050 19306
rect 18109 19303 18143 19306
rect 18211 19272 18245 19936
rect 19470 19432 19526 19448
rect 20714 19432 20770 19448
rect 19470 19376 19526 19392
rect 20714 19376 20770 19392
rect 16704 19238 20160 19272
rect 13796 18836 14244 19048
rect 18211 18844 18245 19238
rect 14020 18826 14152 18836
rect 16704 18810 20160 18844
rect 4666 18768 14102 18802
rect 2010 18746 2458 18756
rect 2002 18544 2458 18746
rect 2002 18534 2450 18544
rect 4666 18360 4700 18768
rect 6239 18700 6273 18768
rect 6341 18700 6375 18768
rect 4842 18666 6375 18700
rect 6191 18619 6192 18620
rect 6192 18618 6193 18619
rect 4769 18607 4814 18618
rect 1144 18349 4700 18360
rect 4780 18370 4814 18607
rect 5060 18420 5116 18446
rect 4780 18349 5464 18370
rect 6180 18349 6191 18360
rect 6239 18355 6273 18666
rect -1796 18293 6191 18349
rect -1889 18265 -1855 18269
rect 4666 18235 4700 18293
rect 4780 18235 4814 18293
rect 4826 18281 4827 18282
rect 4825 18280 4826 18281
rect 4830 18272 5484 18293
rect 5060 18256 5116 18272
rect 6192 18265 6273 18312
rect 6239 18248 6273 18265
rect 6192 18235 6273 18248
rect 6341 18235 6375 18666
rect 9879 18725 9913 18768
rect 9952 18725 9975 18762
rect 10021 18725 10336 18762
rect 11194 18734 13726 18762
rect 11160 18725 13966 18734
rect 14068 18725 14102 18768
rect 16704 18725 16738 18810
rect 16744 18730 17812 18740
rect 18062 18730 18174 18742
rect 16744 18727 18174 18730
rect 16744 18725 18159 18727
rect 18211 18725 18245 18810
rect 9879 18691 18245 18725
rect 9879 18667 10915 18691
rect 10958 18672 13973 18691
rect 10942 18667 13973 18672
rect 9879 18666 13973 18667
rect -1927 18201 6375 18235
rect 4666 17669 4700 18201
rect 4780 17669 4814 18201
rect 5060 18200 5116 18201
rect 5060 17704 5116 17731
rect 6239 17697 6273 18201
rect 4825 17681 4826 17682
rect 4826 17680 4827 17681
rect 5060 17669 5116 17675
rect 6180 17669 6191 17680
rect 4632 17635 6191 17669
rect -1564 17530 -100 17546
rect 4666 17303 4700 17635
rect 4780 17303 4814 17635
rect 4826 17623 4827 17624
rect 4825 17622 4826 17623
rect 6192 17607 6273 17654
rect 6239 17308 6273 17607
rect -2787 17269 5483 17303
rect -20160 16868 -15716 16902
rect -18472 16788 -18438 16868
rect -18370 16822 -18336 16868
rect -15750 16810 -15716 16868
rect -18286 16788 -15716 16810
rect -18506 16776 -15716 16788
rect -18506 16764 -15902 16776
rect -18506 16754 -15891 16764
rect -20102 16748 -20028 16750
rect -20046 16692 -20028 16694
rect -18472 16130 -18438 16754
rect -18408 16748 -18298 16754
rect -18386 16742 -18298 16748
rect -18370 16180 -18336 16742
rect -15890 16726 -15818 16764
rect -15852 16164 -15818 16726
rect -15890 16152 -15802 16164
rect -15750 16152 -15716 16776
rect -18286 16130 -15716 16152
rect -18472 16118 -15716 16130
rect -18472 16096 -15902 16118
rect -18472 16038 -18438 16096
rect -15852 16068 -15818 16072
rect -15750 16038 -15716 16118
rect -18472 16004 -10220 16038
rect -15750 15669 -15716 16004
rect -18513 15464 -15680 15669
rect -20160 15438 -15680 15464
rect -22234 14162 -22222 14192
rect -22206 14162 -22194 14220
rect -22234 14084 -22222 14116
rect -22206 14056 -22194 14116
rect -18513 13314 -15680 15438
rect -18477 12979 -18443 13314
rect -10288 13174 -10075 15669
rect -10288 13163 -9179 13174
rect -10288 13151 -9190 13163
rect -10288 13140 -9179 13151
rect -10288 13071 -10075 13140
rect -10288 13060 -9279 13071
rect -23342 12966 -22668 12979
rect -23973 12945 -22668 12966
rect -20160 12945 -15703 12979
rect -23958 12803 -23338 12945
rect -23288 12911 -22754 12930
rect -23254 12896 -22756 12911
rect -23967 12764 -23338 12803
rect -24040 12678 -23338 12764
rect -23967 12526 -23338 12678
rect -23288 12871 -22722 12877
rect -23288 12865 -23254 12871
rect -22756 12865 -22722 12871
rect -18477 12865 -18443 12945
rect -18375 12899 -18341 12945
rect -15737 12887 -15703 12945
rect -18422 12865 -18341 12872
rect -18282 12865 -15703 12887
rect -23288 12862 -22722 12865
rect -23288 12790 -23254 12862
rect -23131 12850 -22879 12854
rect -23143 12831 -22867 12850
rect -22917 12816 -22906 12819
rect -23109 12801 -22901 12816
rect -23233 12790 -23152 12801
rect -23109 12797 -22824 12801
rect -23288 12748 -23248 12790
rect -23240 12754 -23152 12790
rect -23093 12782 -22906 12797
rect -22905 12754 -22824 12797
rect -23240 12748 -23220 12754
rect -23288 12574 -23254 12748
rect -23186 12716 -23152 12754
rect -22858 12716 -22824 12754
rect -22917 12688 -22906 12699
rect -23093 12654 -22906 12688
rect -22756 12574 -22722 12862
rect -18511 12853 -15703 12865
rect -18511 12841 -15898 12853
rect -18511 12831 -15887 12841
rect -23288 12540 -22722 12574
rect -23967 12472 -23933 12526
rect -23967 12235 -23338 12472
rect -23958 12050 -23338 12235
rect -23288 12420 -22722 12454
rect -23288 12207 -23254 12420
rect -22917 12340 -22906 12351
rect -23240 12213 -23238 12300
rect -23233 12278 -23152 12325
rect -23093 12306 -22906 12340
rect -22905 12278 -22824 12325
rect -23186 12224 -23152 12278
rect -22858 12241 -22824 12278
rect -22866 12232 -22814 12241
rect -22864 12228 -22818 12232
rect -22858 12224 -22824 12228
rect -23104 12219 -22906 12223
rect -23093 12207 -22917 12212
rect -22894 12207 -22786 12213
rect -22756 12207 -22722 12420
rect -23288 12173 -22722 12207
rect -23288 12098 -23254 12173
rect -22756 12098 -22722 12173
rect -23288 12064 -22722 12098
rect -18477 12207 -18443 12831
rect -18422 12825 -18294 12831
rect -18391 12819 -18294 12825
rect -18375 12257 -18341 12819
rect -15886 12803 -15805 12850
rect -15839 12241 -15805 12803
rect -15886 12229 -15789 12241
rect -15737 12229 -15703 12853
rect -18282 12207 -15703 12229
rect -18477 12195 -15703 12207
rect -18477 12173 -15898 12195
rect -15886 12183 -15758 12192
rect -18477 12115 -18443 12173
rect -15839 12145 -15805 12149
rect -15737 12115 -15703 12195
rect -10288 12115 -10075 13060
rect -10066 13026 -9279 13060
rect -18477 12081 -10075 12115
rect -23460 11446 -23260 11456
rect -23488 11418 -23232 11428
rect -17594 10980 -16130 10996
rect -18822 10851 -18766 10868
rect -18420 10851 -17538 10868
rect -16186 10851 -15886 10868
rect -18822 10795 -18766 10812
rect -15737 10598 -15703 12081
rect -10288 12045 -10075 12081
rect -14478 11322 -14472 11464
rect -14484 11300 -14472 11322
rect -14488 11274 -14472 11300
rect -14488 11244 -14462 11274
rect -14488 11140 -14462 11168
rect -14488 11112 -14466 11140
rect -14484 11104 -14466 11112
rect -14478 10646 -14466 11104
rect -18490 10562 -15667 10598
rect -10252 10562 -10218 12045
rect -10150 10562 -10116 12045
rect -9290 10656 -9279 10667
rect -10066 10622 -9279 10656
rect -18490 10528 -10202 10562
rect -10177 10555 -10106 10562
rect -10197 10542 -10106 10555
rect -9240 10542 -9206 13140
rect -18490 10448 -15667 10528
rect -18490 10414 -10292 10448
rect -10286 10420 -10276 10448
rect -10252 10420 -10218 10528
rect -10197 10508 -9172 10542
rect -10286 10414 -10218 10420
rect -18490 9575 -15667 10414
rect -14492 10408 -14422 10410
rect -10276 10398 -10218 10414
rect -10276 10386 -10202 10398
rect -14436 10352 -14422 10354
rect -10252 10316 -10184 10386
rect -10166 10344 -10150 10444
rect -10252 9868 -10170 10316
rect -14354 9800 -13982 9828
rect -10252 9818 -10184 9868
rect -10166 9840 -10142 10344
rect -10252 9806 -10202 9818
rect -14392 9762 -13944 9790
rect -10286 9762 -10276 9790
rect -10252 9762 -10218 9806
rect -10166 9802 -10150 9840
rect -10286 9756 -10218 9762
rect -10276 9740 -10218 9756
rect -10276 9728 -10202 9740
rect -20160 9541 -15667 9575
rect -18490 9391 -15667 9541
rect -10252 9664 -10184 9728
rect -10166 9692 -10150 9786
rect -10140 9692 -10106 10508
rect -10166 9664 -10106 9692
rect -20066 8668 -20064 8810
rect -20076 8646 -20064 8668
rect -20080 8620 -20064 8646
rect -20080 8590 -20054 8620
rect -19362 8520 -19330 8590
rect -20080 8486 -20054 8514
rect -19328 8486 -19296 8624
rect -20080 8458 -20058 8486
rect -20076 8450 -20058 8458
rect -21620 8020 -21468 8044
rect -21340 8034 -21194 8042
rect -21362 8020 -21194 8034
rect -21592 7992 -21496 8016
rect -21912 7944 -21878 7955
rect -21584 7944 -21550 7955
rect -22050 7908 -21412 7944
rect -21362 7908 -21328 8020
rect -21312 7992 -21222 8014
rect -21260 7922 -21226 7955
rect -20950 7922 -20916 7955
rect -20848 7908 -20814 8034
rect -20640 7960 -20636 8134
rect -20606 7994 -20602 8168
rect -20066 7992 -20058 8450
rect -18454 7908 -18420 9391
rect -10252 9268 -10106 9664
rect -9138 9268 -9104 15732
rect -11460 9198 -9068 9268
rect -17978 9160 -16576 9174
rect -22050 7874 -15698 7908
rect -22050 7726 -21412 7874
rect -21266 7806 -20910 7828
rect -21362 7780 -20814 7806
rect -18454 7794 -18420 7874
rect -18352 7856 -18312 7874
rect -18358 7832 -18312 7856
rect -18352 7828 -18318 7832
rect -15732 7816 -15698 7874
rect -18268 7794 -15698 7816
rect -18488 7782 -15698 7794
rect -18488 7770 -15884 7782
rect -18488 7760 -15873 7770
rect -23944 7148 -23910 7180
rect -23978 7114 -23876 7146
rect -18454 7136 -18420 7760
rect -18390 7754 -18280 7760
rect -18368 7748 -18280 7754
rect -18352 7186 -18318 7748
rect -15872 7732 -15800 7770
rect -15834 7170 -15800 7732
rect -15872 7158 -15784 7170
rect -15732 7158 -15698 7782
rect -18268 7136 -15698 7158
rect -18454 7124 -15698 7136
rect -18454 7102 -15884 7124
rect -23436 6680 -22256 7052
rect -18454 7044 -18420 7102
rect -15834 7074 -15800 7078
rect -15732 7044 -15698 7124
rect -11460 7854 -9058 9198
rect -11460 7818 -9068 7854
rect -11460 7044 -10070 7818
rect -18454 7010 -10070 7044
rect -23570 6506 -22168 6520
rect -19758 6478 -19080 6570
rect -18312 6538 -17764 6572
rect -18312 6510 -18278 6538
rect -17798 6510 -17764 6538
rect -18346 6478 -18244 6510
rect -17832 6478 -17730 6510
rect -17714 6478 -17076 6626
rect -19758 6444 -15884 6478
rect -19758 6236 -19080 6444
rect -18430 6406 -18344 6424
rect -20160 6094 -19080 6236
rect -18312 6256 -18278 6444
rect -18248 6414 -18176 6444
rect -18126 6432 -17950 6444
rect -18126 6424 -17939 6432
rect -17938 6414 -17866 6444
rect -18210 6380 -18176 6414
rect -17908 6410 -17904 6414
rect -17950 6370 -17939 6381
rect -17900 6380 -17866 6414
rect -18126 6336 -17939 6370
rect -17908 6360 -17904 6380
rect -17936 6332 -17904 6352
rect -17798 6256 -17764 6444
rect -18312 6222 -17764 6256
rect -17714 6164 -17076 6444
rect -20160 6024 -19724 6094
rect -18312 6062 -17764 6096
rect -18312 5780 -18278 6062
rect -17950 5982 -17939 5993
rect -18248 5938 -18176 5976
rect -18126 5948 -17939 5982
rect -17938 5938 -17866 5976
rect -18210 5904 -18176 5938
rect -18166 5904 -17910 5928
rect -17900 5904 -17866 5938
rect -17950 5900 -17939 5904
rect -18138 5876 -17938 5900
rect -18126 5860 -17939 5876
rect -17798 5814 -17764 6062
rect -18272 5786 -17764 5814
rect -17798 5780 -17764 5786
rect -18312 5746 -17764 5780
rect -17714 5688 -17076 6150
rect -17238 5668 -17182 5688
rect -27427 5350 -27219 5380
rect -15732 5367 -15698 7010
rect -11460 6974 -10070 7010
rect -27461 5316 -27185 5346
rect -24082 5331 -21847 5367
rect -17191 5336 -15662 5367
rect -25815 5297 -21847 5331
rect -29028 4026 -27848 4398
rect -25911 3531 -25877 5235
rect -25435 5229 -25401 5267
rect -25304 5229 -24124 5252
rect -24082 5229 -21847 5297
rect -25735 5195 -21847 5229
rect -25435 3531 -25401 5195
rect -25304 5147 -24124 5195
rect -25332 5136 -24124 5147
rect -25321 4880 -24124 5136
rect -25321 3916 -25276 4880
rect -25139 4320 -25094 4880
rect -24663 4320 -24618 4880
rect -25156 3916 -25086 4320
rect -24680 3916 -24610 4320
rect -25350 3864 -24610 3916
rect -25350 3632 -24672 3864
rect -25368 3556 -24672 3632
rect -25350 3531 -24672 3556
rect -24663 3531 -24618 3864
rect -24481 3531 -24436 4880
rect -24082 4390 -21847 5195
rect -20840 5331 -15662 5336
rect -12120 5331 -11699 5367
rect -20840 5302 -11699 5331
rect -20840 5162 -20806 5302
rect -20364 5272 -20330 5302
rect -17322 5272 -17288 5302
rect -17191 5297 -11699 5302
rect -17191 5272 -15662 5297
rect -20364 5234 -20326 5272
rect -20066 5234 -15662 5272
rect -20664 5229 -15662 5234
rect -15287 5229 -15253 5267
rect -13637 5245 -13626 5256
rect -13614 5245 -13603 5256
rect -13637 5229 -13603 5245
rect -12120 5229 -11699 5297
rect -20664 5200 -13227 5229
rect -20364 5174 -20330 5200
rect -18172 5194 -18144 5200
rect -17520 5194 -17492 5200
rect -18200 5174 -18172 5194
rect -18144 5174 -18116 5194
rect -17548 5174 -17520 5194
rect -17492 5174 -17464 5194
rect -17322 5174 -17288 5200
rect -17191 5195 -13227 5200
rect -12598 5195 -12569 5229
rect -17191 5174 -15662 5195
rect -20680 5162 -15662 5174
rect -20874 5128 -15662 5162
rect -20840 4504 -20806 5128
rect -20726 4504 -20692 5128
rect -20680 5116 -20679 5117
rect -20681 5115 -20680 5116
rect -20681 4516 -20680 4517
rect -20680 4515 -20679 4516
rect -20364 4504 -20330 5128
rect -20250 4504 -20216 5128
rect -20068 4714 -20023 5128
rect -19592 4802 -19547 5128
rect -19410 4802 -19365 5128
rect -18934 4802 -18889 5128
rect -18752 4802 -18707 5128
rect -18276 4802 -18231 5128
rect -18094 4802 -18049 5128
rect -17618 4802 -17573 5128
rect -17436 4802 -17391 5128
rect -17322 4802 -17288 5128
rect -17191 4802 -15662 5128
rect -19920 4770 -15662 4802
rect -15287 4770 -15253 5195
rect -15184 5136 -15128 5147
rect -15078 5136 -15022 5147
rect -14526 5136 -14470 5147
rect -14420 5136 -14364 5147
rect -13868 5136 -13812 5147
rect -13762 5136 -13706 5147
rect -15173 4770 -15128 5136
rect -15067 4770 -15022 5136
rect -19920 4736 -14794 4770
rect -19920 4715 -15662 4736
rect -15287 4715 -15253 4736
rect -15173 4715 -15128 4736
rect -15067 4715 -15022 4736
rect -20068 4504 -20034 4714
rect -19920 4668 -14923 4715
rect -19920 4634 -15581 4668
rect -15538 4634 -14923 4668
rect -19920 4504 -15662 4634
rect -15611 4575 -15555 4586
rect -20874 4470 -15662 4504
rect -20840 4390 -20806 4470
rect -20726 4390 -20692 4470
rect -20364 4390 -20330 4470
rect -20250 4390 -20205 4470
rect -20068 4398 -20023 4470
rect -19920 4398 -15662 4470
rect -20160 4396 -15662 4398
rect -20100 4390 -15662 4396
rect -24082 4356 -15662 4390
rect -24082 4320 -21847 4356
rect -24005 3531 -23960 4320
rect -23940 3954 -23912 3958
rect -23884 3954 -23856 3958
rect -23823 3954 -23778 4320
rect -23347 4304 -23302 4320
rect -23368 4182 -23298 4304
rect -23368 4110 -23272 4182
rect -23368 3954 -23298 4110
rect -23940 3848 -23298 3954
rect -23270 3936 -23242 3958
rect -23214 3936 -23186 3958
rect -23165 3936 -23120 4320
rect -23270 3902 -22704 3936
rect -23270 3858 -23236 3902
rect -23940 3532 -23302 3848
rect -23278 3808 -23236 3858
rect -23214 3864 -23186 3902
rect -23214 3808 -23174 3864
rect -23278 3802 -23230 3808
rect -23214 3807 -23202 3808
rect -23165 3807 -23120 3902
rect -23086 3822 -22888 3833
rect -23215 3802 -23118 3807
rect -23270 3682 -23230 3802
rect -23222 3794 -23118 3802
rect -23222 3760 -23100 3794
rect -23075 3788 -22888 3822
rect -22887 3760 -22759 3807
rect -23222 3682 -23202 3760
rect -23168 3733 -23100 3760
rect -23176 3722 -23100 3733
rect -22840 3722 -22759 3760
rect -23278 3626 -23230 3682
rect -23940 3531 -23912 3532
rect -23884 3531 -23856 3532
rect -23823 3531 -23778 3532
rect -27683 3497 -23751 3531
rect -25911 3482 -25877 3497
rect -25803 3482 -25757 3497
rect -25435 3482 -25401 3497
rect -25350 3482 -24672 3497
rect -24663 3482 -24618 3497
rect -24481 3482 -24436 3497
rect -24261 3482 -24227 3497
rect -26330 3476 -24106 3482
rect -24005 3476 -23960 3497
rect -23940 3478 -23912 3497
rect -23884 3478 -23856 3497
rect -23823 3478 -23751 3497
rect -23347 3478 -23302 3532
rect -23270 3608 -23230 3626
rect -23214 3608 -23202 3682
rect -23270 3580 -23236 3608
rect -23214 3580 -23174 3608
rect -23165 3580 -23120 3722
rect -23086 3694 -22888 3705
rect -23075 3660 -22888 3694
rect -22738 3580 -22704 3902
rect -23270 3572 -22704 3580
rect -22689 3572 -22644 4320
rect -22562 3844 -22534 3958
rect -22562 3572 -22534 3658
rect -22507 3572 -22462 4320
rect -22393 3572 -22359 4320
rect -23270 3546 -21847 3572
rect -23270 3486 -23242 3546
rect -23214 3486 -23186 3546
rect -23940 3476 -23302 3478
rect -26330 3467 -23302 3476
rect -27779 2677 -27745 3435
rect -27303 3429 -27269 3467
rect -26426 3448 -23302 3467
rect -23165 3460 -23120 3546
rect -22744 3536 -21847 3546
rect -20840 3536 -20806 4356
rect -20364 3536 -20330 4356
rect -20250 3536 -20205 4356
rect -20100 4328 -15662 4356
rect -20068 4274 -20023 4328
rect -19920 4320 -15662 4328
rect -19920 4274 -16776 4320
rect -20100 4232 -16776 4274
rect -20106 4226 -16776 4232
rect -20174 3536 -20146 3958
rect -20068 3536 -20023 4226
rect -19920 3864 -16776 4226
rect -19592 3536 -19547 3864
rect -19522 3536 -19494 3864
rect -19466 3536 -19438 3864
rect -19410 3536 -19365 3864
rect -18934 3536 -18889 3864
rect -18864 3536 -18836 3864
rect -18808 3536 -18780 3864
rect -18752 3536 -18707 3864
rect -22744 3502 -18680 3536
rect -22744 3460 -21847 3502
rect -26426 3429 -26392 3448
rect -25911 3429 -25877 3448
rect -25809 3429 -23302 3448
rect -27303 3418 -23302 3429
rect -23270 3434 -21847 3460
rect -21390 3440 -21362 3472
rect -21334 3440 -21306 3472
rect -20840 3434 -20806 3502
rect -20732 3472 -20686 3502
rect -20364 3472 -20330 3502
rect -20250 3472 -20205 3502
rect -20174 3472 -20146 3502
rect -20068 3472 -20023 3502
rect -19592 3472 -19547 3502
rect -19522 3472 -19494 3502
rect -19466 3472 -19438 3502
rect -19410 3472 -19365 3502
rect -19190 3472 -19156 3502
rect -18934 3472 -18889 3502
rect -18864 3472 -18836 3502
rect -20738 3434 -18818 3472
rect -23270 3426 -18818 3434
rect -27615 3389 -27548 3402
rect -27303 3395 -23313 3418
rect -31407 2643 -27475 2677
rect -31503 877 -31469 2581
rect -31027 2575 -30993 2613
rect -27985 2591 -27974 2602
rect -27962 2591 -27951 2602
rect -27985 2575 -27951 2591
rect -27779 2575 -27745 2643
rect -27665 2609 -27618 2622
rect -27665 2606 -27617 2609
rect -27677 2575 -27617 2606
rect -31327 2541 -27617 2575
rect -31027 877 -30993 2541
rect -30924 2482 -30868 2493
rect -30742 2482 -30686 2493
rect -30266 2482 -30210 2493
rect -30084 2482 -30028 2493
rect -29608 2482 -29563 2493
rect -29426 2482 -29381 2493
rect -28950 2482 -28905 2493
rect -28768 2482 -28723 2493
rect -28292 2482 -28247 2493
rect -28110 2482 -28065 2493
rect -30913 2226 -30192 2482
rect -30913 877 -30868 2226
rect -30852 877 -30824 2158
rect -30731 877 -30686 2226
rect -30255 877 -30210 2226
rect -30194 877 -30166 2158
rect -30138 877 -30110 2158
rect -30073 877 -30028 2482
rect -33275 843 -29819 877
rect -31503 -5655 -31469 843
rect -31027 822 -30993 843
rect -30913 840 -30868 843
rect -30913 822 -30879 840
rect -31389 806 -31342 822
rect -31401 775 -31342 806
rect -31311 781 -31264 822
rect -31328 775 -31264 781
rect -31027 775 -30980 822
rect -30913 775 -30866 822
rect -30852 794 -30824 843
rect -30731 840 -30686 843
rect -30255 840 -30210 843
rect -30731 822 -30697 840
rect -30255 822 -30221 840
rect -30731 775 -30684 822
rect -30653 775 -30606 822
rect -30255 775 -30208 822
rect -30194 794 -30166 843
rect -30138 794 -30110 843
rect -30073 840 -30028 843
rect -30073 822 -30039 840
rect -30073 775 -30026 822
rect -29995 775 -29948 822
rect -31401 741 -31264 775
rect -31221 741 -30606 775
rect -30563 741 -29948 775
rect -31401 735 -31299 741
rect -31401 694 -31343 735
rect -31272 707 -31271 741
rect -31389 450 -31355 694
rect -31294 682 -31249 693
rect -31389 -1014 -31349 450
rect -31332 -958 -31321 394
rect -31389 -5494 -31355 -1014
rect -31345 -5170 -31314 -3768
rect -31289 -5198 -31286 -3740
rect -31283 -5506 -31249 682
rect -31027 -5506 -30993 741
rect -30913 -5494 -30879 741
rect -30731 -5494 -30697 741
rect -30636 682 -30591 693
rect -30625 -1316 -30591 682
rect -30694 -1324 -30482 -1316
rect -30694 -1764 -30282 -1324
rect -30625 -5506 -30591 -1764
rect -30494 -1772 -30282 -1764
rect -30255 -5494 -30221 741
rect -30073 -5494 -30039 741
rect -29978 682 -29933 693
rect -29967 -1324 -29933 682
rect -29853 -1316 -29819 843
rect -29631 840 -29616 1946
rect -29853 -1324 -29636 -1316
rect -30018 -1764 -29636 -1324
rect -30018 -1772 -29806 -1764
rect -29967 -5506 -29933 -1772
rect -31295 -5553 -31236 -5506
rect -31027 -5553 -30980 -5506
rect -30637 -5553 -30578 -5506
rect -29979 -5553 -29921 -5506
rect -31327 -5587 -29921 -5553
rect -31395 -5649 -31372 -5593
rect -31295 -5603 -31237 -5587
rect -31283 -5655 -31249 -5621
rect -31027 -5655 -30993 -5587
rect -30690 -5600 -30579 -5587
rect -30637 -5602 -30579 -5600
rect -30662 -5603 -30579 -5602
rect -29979 -5603 -29921 -5587
rect -30662 -5655 -30631 -5603
rect -29936 -5618 -29921 -5603
rect -29853 -5553 -29819 -1772
rect -29597 -5494 -29563 2482
rect -29532 -3192 -29504 2158
rect -29476 -3192 -29448 2158
rect -29532 -5547 -29504 -3378
rect -29476 -5547 -29448 -3378
rect -29415 -5494 -29381 2482
rect -29164 -1324 -29160 -1316
rect -29152 -1764 -29148 -1324
rect -28939 -2458 -28905 2482
rect -28939 -2648 -28894 -2458
rect -28862 -2648 -28834 2158
rect -28806 -2648 -28778 2158
rect -28757 -2458 -28723 2482
rect -28281 918 -28247 2482
rect -28154 918 -28126 2158
rect -28099 918 -28065 2482
rect -27985 918 -27951 2541
rect -27779 918 -27745 2541
rect -27677 2532 -27635 2541
rect -27677 2494 -27631 2532
rect -27665 918 -27631 2494
rect -27623 2493 -27597 2498
rect -27623 918 -27589 2493
rect -27509 918 -27475 2643
rect -27303 918 -27269 3395
rect -27100 3389 -27072 3395
rect -26442 3389 -26392 3395
rect -27200 3336 -27155 3347
rect -27128 3346 -27100 3389
rect -27018 3336 -26973 3347
rect -26542 3336 -26497 3347
rect -26470 3346 -26442 3389
rect -26426 3346 -26386 3389
rect -25911 3380 -25877 3395
rect -25809 3380 -25750 3395
rect -25435 3380 -25401 3395
rect -25333 3380 -25274 3395
rect -25139 3380 -25092 3395
rect -24675 3380 -24616 3395
rect -24481 3380 -24434 3395
rect -24282 3380 -24227 3395
rect -26266 3361 -24227 3380
rect -26250 3357 -24227 3361
rect -25911 3348 -24227 3357
rect -27189 2692 -27155 3336
rect -27007 2692 -26973 3336
rect -26531 2692 -26497 3336
rect -26426 2718 -26392 3346
rect -26360 3336 -26315 3347
rect -26250 3346 -24227 3348
rect -26349 3298 -26315 3336
rect -26312 3298 -26281 3303
rect -25911 3299 -25827 3346
rect -26349 3287 -26278 3298
rect -26349 2718 -26315 3287
rect -26312 2718 -26278 3287
rect -25911 2718 -25877 3299
rect -25873 2802 -25839 3299
rect -25797 2802 -25763 3346
rect -25702 3336 -25657 3346
rect -25691 2802 -25657 3336
rect -25873 2718 -25828 2802
rect -25797 2718 -25752 2802
rect -25691 2718 -25646 2802
rect -25435 2718 -25401 3346
rect -25321 2802 -25287 3346
rect -25227 3299 -25169 3346
rect -25215 2802 -25181 3299
rect -25139 2802 -25105 3346
rect -25044 3336 -24999 3346
rect -25033 2802 -24999 3336
rect -24663 2802 -24629 3346
rect -24569 3299 -24511 3346
rect -24557 2802 -24523 3299
rect -24481 2802 -24447 3346
rect -24386 3336 -24341 3346
rect -24375 2802 -24341 3336
rect -24261 3298 -24227 3346
rect -24261 2802 -24220 3298
rect -25321 2718 -25276 2802
rect -25215 2718 -25170 2802
rect -25139 2718 -25094 2802
rect -25033 2718 -24988 2802
rect -24663 2718 -24618 2802
rect -24557 2718 -24512 2802
rect -24481 2718 -24436 2802
rect -24375 2718 -24330 2802
rect -24261 2718 -24209 2802
rect -24140 2718 -24106 3395
rect -24082 3088 -24072 3395
rect -24017 3348 -23313 3395
rect -24005 3346 -23313 3348
rect -24005 3088 -23960 3346
rect -24005 2802 -23971 3088
rect -23940 3056 -23313 3346
rect -23270 3402 -23236 3426
rect -23165 3418 -23120 3426
rect -23270 3388 -23214 3402
rect -23270 3346 -23236 3388
rect -23214 3346 -23186 3388
rect -23270 3332 -23214 3346
rect -23270 3104 -23236 3332
rect -23165 3331 -23131 3418
rect -22744 3400 -18818 3426
rect -22899 3346 -22888 3357
rect -23215 3318 -23118 3331
rect -23215 3284 -23100 3318
rect -23075 3312 -22888 3346
rect -22887 3284 -22806 3331
rect -23168 3257 -23100 3284
rect -23176 3246 -23100 3257
rect -22840 3246 -22806 3284
rect -23165 3104 -23131 3246
rect -22899 3218 -22888 3229
rect -23075 3184 -22888 3218
rect -22744 3104 -21847 3400
rect -21362 3394 -21334 3400
rect -21471 3350 -21415 3361
rect -23270 3070 -21847 3104
rect -23899 2802 -23865 3056
rect -23823 2802 -23789 3056
rect -23785 2802 -23751 3056
rect -24005 2718 -23960 2802
rect -23899 2718 -23854 2802
rect -23823 2718 -23751 2802
rect -23347 2802 -23313 3056
rect -23165 2802 -23131 3070
rect -23347 2718 -23302 2802
rect -23165 2718 -23120 2802
rect -22744 2718 -21847 3070
rect -26468 2713 -21847 2718
rect -21460 2713 -21415 3350
rect -21390 3346 -21362 3394
rect -21334 3346 -21306 3394
rect -20840 3361 -20806 3400
rect -20738 3394 -20676 3400
rect -20738 3362 -20680 3394
rect -21289 3350 -21233 3361
rect -21278 2713 -21233 3350
rect -20840 3350 -20757 3361
rect -20840 3094 -20806 3350
rect -20802 3094 -20757 3350
rect -20732 3346 -20681 3362
rect -20676 3361 -20630 3394
rect -20676 3350 -20575 3361
rect -20676 3346 -20630 3350
rect -20726 3094 -20681 3346
rect -20620 3094 -20575 3350
rect -20364 3094 -20330 3400
rect -20262 3362 -20204 3400
rect -20250 3094 -20205 3362
rect -20155 3350 -20099 3361
rect -20144 3094 -20099 3350
rect -20068 3094 -20023 3400
rect -19604 3362 -19546 3400
rect -19973 3350 -19917 3361
rect -19962 3094 -19917 3350
rect -19592 3094 -19547 3362
rect -19497 3350 -19441 3361
rect -19486 3094 -19441 3350
rect -19410 3094 -19365 3400
rect -19315 3350 -19259 3361
rect -19304 3094 -19259 3350
rect -19190 3094 -19156 3400
rect -18946 3362 -18836 3400
rect -18808 3362 -18780 3502
rect -18934 3361 -18836 3362
rect -18834 3361 -18780 3362
rect -18934 3350 -18780 3361
rect -18934 3346 -18836 3350
rect -18834 3346 -18780 3350
rect -18934 3094 -18889 3346
rect -18828 3094 -18783 3346
rect -18752 3094 -18680 3502
rect -18276 3100 -18231 3864
rect -18200 3346 -18172 3864
rect -18144 3346 -18116 3864
rect -18094 3100 -18049 3864
rect -17618 3100 -17573 3864
rect -17548 3410 -17520 3864
rect -17492 3346 -17464 3864
rect -17436 3100 -17391 3864
rect -17322 3100 -17288 3864
rect -17191 3531 -16776 3864
rect -16426 3531 -16420 3958
rect -16372 3565 -16338 4320
rect -16322 3830 -16298 3958
rect -16258 3599 -16213 4320
rect -16383 3534 -16338 3565
rect -16322 3534 -16298 3590
rect -15725 3587 -15680 4320
rect -15600 3599 -15555 4575
rect -15287 3587 -15253 4634
rect -15173 3632 -15128 4634
rect -15067 3632 -15022 4634
rect -14953 4575 -14897 4586
rect -15216 3587 -15022 3632
rect -14942 3599 -14897 4575
rect -16243 3540 -14923 3587
rect -16383 3531 -16298 3534
rect -16196 3531 -15581 3540
rect -15538 3531 -14923 3540
rect -14828 3531 -14794 4736
rect -14515 3958 -14470 5136
rect -14409 3958 -14364 5136
rect -13857 4768 -13812 5136
rect -13751 4768 -13706 5136
rect -13637 4768 -13603 5195
rect -12560 5157 -12531 5224
rect -12479 5195 -11699 5229
rect -14515 3531 -14430 3958
rect -14415 3531 -14364 3958
rect -14286 4734 -12708 4768
rect -14286 3531 -14252 4734
rect -13857 4713 -13812 4734
rect -13751 4713 -13706 4734
rect -13637 4713 -13603 4734
rect -14157 4666 -13495 4713
rect -13199 4682 -13152 4713
rect -13211 4666 -13152 4682
rect -12884 4666 -12837 4713
rect -14110 4632 -13495 4666
rect -13452 4634 -12837 4666
rect -13458 4632 -12837 4634
rect -14183 4573 -14127 4584
rect -14172 3597 -14127 4573
rect -13857 4234 -13812 4632
rect -13751 4282 -13706 4632
rect -13766 4234 -13696 4282
rect -13948 4080 -13696 4234
rect -13857 3585 -13812 4080
rect -13766 3826 -13696 4080
rect -13751 3585 -13706 3826
rect -13637 3585 -13603 4632
rect -13458 4598 -13400 4600
rect -13211 4585 -13153 4632
rect -13525 4573 -13469 4584
rect -13514 3597 -13469 4573
rect -13199 4422 -13165 4585
rect -12867 4573 -12822 4584
rect -12856 4422 -12822 4573
rect -13199 4304 -13154 4422
rect -13220 4230 -13150 4304
rect -13300 4084 -13050 4230
rect -13220 3848 -13150 4084
rect -13199 3585 -13154 3848
rect -12856 3597 -12811 4422
rect -14157 3538 -12837 3585
rect -14110 3531 -13495 3538
rect -17191 3504 -13495 3531
rect -13452 3504 -12837 3538
rect -17191 3497 -13603 3504
rect -17191 3476 -16776 3497
rect -16426 3490 -16420 3497
rect -16383 3476 -16338 3497
rect -15737 3490 -15679 3497
rect -15725 3482 -15691 3490
rect -15604 3482 -15560 3497
rect -15287 3482 -15253 3497
rect -15173 3482 -15128 3497
rect -15116 3496 -15105 3497
rect -15067 3482 -15022 3497
rect -14828 3482 -14794 3497
rect -14515 3490 -14430 3497
rect -14515 3482 -14470 3490
rect -14415 3482 -14364 3497
rect -14286 3482 -14252 3497
rect -16278 3476 -13958 3482
rect -17191 3448 -13958 3476
rect -17191 3438 -16244 3448
rect -15731 3438 -15713 3448
rect -15703 3438 -15685 3448
rect -15604 3444 -15560 3448
rect -15287 3438 -15253 3448
rect -15173 3445 -15128 3448
rect -15185 3438 -15127 3445
rect -15073 3438 -15022 3448
rect -14890 3438 -14190 3448
rect -17191 3436 -14190 3438
rect -13992 3436 -13958 3448
rect -13857 3445 -13812 3497
rect -13794 3466 -13789 3497
rect -13751 3463 -13706 3497
rect -13869 3436 -13811 3445
rect -13757 3436 -13706 3463
rect -13637 3436 -13603 3497
rect -13211 3488 -13153 3504
rect -12742 3436 -12708 4734
rect -17191 3429 -12708 3436
rect -17191 3427 -14364 3429
rect -17191 3418 -14362 3427
rect -14347 3418 -12708 3429
rect -17191 3404 -12708 3418
rect -17191 3395 -16343 3404
rect -16337 3402 -12708 3404
rect -16337 3395 -13706 3402
rect -17191 3100 -16776 3395
rect -16476 3389 -16399 3395
rect -16389 3361 -16343 3395
rect -16333 3389 -16244 3395
rect -20942 2713 -18634 3094
rect -18364 3064 -16776 3100
rect -16383 3064 -16349 3361
rect -16278 3064 -16244 3389
rect -15737 3380 -15678 3395
rect -15287 3380 -15253 3395
rect -15185 3380 -15126 3395
rect -15067 3380 -15020 3395
rect -14527 3380 -14468 3395
rect -14409 3380 -14362 3395
rect -14134 3380 -14087 3395
rect -16118 3361 -14087 3380
rect -16102 3346 -14087 3361
rect -15737 3299 -15679 3346
rect -16175 3287 -16130 3298
rect -16164 3144 -16130 3287
rect -16164 3064 -16119 3144
rect -18364 3030 -16092 3064
rect -18364 2962 -16776 3030
rect -16278 3009 -16244 3030
rect -16383 2978 -16336 3009
rect -16395 2962 -16336 2978
rect -16278 2962 -16231 3009
rect -18364 2928 -16231 2962
rect -18364 2718 -16776 2928
rect -16395 2881 -16337 2928
rect -16383 2802 -16349 2881
rect -16278 2880 -16244 2928
rect -16240 2880 -16210 2885
rect -16278 2869 -16206 2880
rect -16383 2718 -16338 2802
rect -16278 2718 -16244 2869
rect -16240 2802 -16206 2869
rect -16240 2718 -16195 2802
rect -16164 2718 -16092 3030
rect -15725 2802 -15691 3299
rect -15725 2718 -15680 2802
rect -15287 2718 -15253 3346
rect -15173 2802 -15139 3346
rect -15079 3299 -15021 3346
rect -15067 2802 -15033 3299
rect -15173 2718 -15128 2802
rect -15067 2718 -15022 2802
rect -14515 2718 -14481 3346
rect -14421 3299 -14363 3346
rect -14409 2718 -14375 3299
rect -14117 3287 -14072 3298
rect -14106 2718 -14072 3287
rect -13992 2718 -13958 3395
rect -13869 3348 -13811 3395
rect -13785 3389 -13767 3395
rect -13757 3361 -13706 3395
rect -13857 3156 -13812 3348
rect -13751 3156 -13706 3361
rect -13637 3156 -13603 3402
rect -13199 3156 -13165 3190
rect -12541 3156 -12507 5136
rect -12120 4806 -11699 5195
rect -11460 5336 -9022 5372
rect -8794 5336 -8760 17140
rect -8680 14582 -8646 17050
rect -8692 14548 -8176 14582
rect -8680 14518 -8646 14548
rect -8222 14518 -8188 14548
rect -8680 14480 -8296 14518
rect -8250 14480 -8188 14518
rect -8170 14510 -8154 14548
rect -8680 6922 -8646 14480
rect -8618 14446 -8188 14480
rect -8222 7062 -8188 14446
rect -8250 7024 -8188 7062
rect -8634 6990 -8188 7024
rect -8222 6922 -8188 6990
rect -8166 6922 -8154 6962
rect -8698 6888 -8176 6922
rect -8170 6888 -8154 6922
rect -8200 6800 -8188 6888
rect -8166 6834 -8154 6888
rect -8108 5336 -8074 17140
rect -2883 12268 -2849 17207
rect -1991 15752 -1957 17269
rect -1936 17189 -1808 17201
rect 4666 17200 4700 17269
rect 1144 17189 4700 17200
rect 4780 17189 4814 17269
rect 5288 17189 5299 17200
rect -1936 17155 5299 17189
rect -1905 17143 -1808 17155
rect -1951 17114 -1895 17128
rect -1908 17098 -1895 17114
rect -1936 17070 -1895 17072
rect -1889 17039 -1855 17143
rect 4666 17128 4700 17155
rect -1849 17098 4774 17128
rect 4666 17072 4700 17098
rect -1849 17070 4774 17072
rect 4666 17022 4700 17070
rect 1144 17011 4700 17022
rect 4780 17011 4814 17155
rect 4820 17098 5116 17128
rect 5300 17127 5381 17174
rect 4820 17070 5116 17072
rect 5060 17042 5116 17070
rect 5347 17024 5381 17127
rect 5300 17011 5381 17024
rect 5449 17022 5483 17269
rect 6239 17039 6320 17308
rect 5446 17011 6191 17022
rect -1936 16949 -1855 16996
rect -1796 16977 6191 17011
rect -1889 16544 -1855 16949
rect -1936 16543 -1855 16544
rect -1936 16531 -1808 16543
rect 4666 16542 4700 16977
rect 1144 16531 4700 16542
rect 4780 16531 4814 16977
rect 5347 16559 5381 16977
rect 5288 16531 5299 16542
rect -1936 16497 5299 16531
rect -1905 16485 -1808 16497
rect -1889 16381 -1855 16485
rect 4666 16470 4700 16497
rect -1849 16436 4774 16470
rect 4666 16414 4700 16436
rect -1849 16380 4774 16414
rect 4666 16364 4700 16380
rect 1144 16353 4700 16364
rect 4780 16353 4814 16497
rect 4820 16436 5116 16470
rect 5300 16469 5381 16516
rect 4820 16380 5116 16414
rect 5347 16366 5381 16469
rect 5300 16353 5381 16366
rect 5449 16364 5483 16977
rect 6192 16949 6320 16996
rect 6239 16381 6320 16949
rect 5446 16353 6191 16364
rect -1936 16291 -1855 16338
rect -1796 16319 6191 16353
rect -1889 15886 -1855 16291
rect -1936 15885 -1855 15886
rect -1936 15873 -1808 15885
rect 4666 15884 4700 16319
rect 1144 15873 4700 15884
rect 4780 15873 4814 16319
rect 5347 15901 5381 16319
rect 5288 15873 5299 15884
rect -1936 15839 5299 15873
rect -1905 15827 -1808 15839
rect -1908 15778 -1895 15780
rect -1991 15722 -1895 15752
rect -1889 15723 -1855 15827
rect 4666 15780 4700 15839
rect -1849 15778 4774 15780
rect 4666 15752 4700 15778
rect -1849 15722 4774 15752
rect -1991 15581 -1957 15722
rect 4666 15706 4700 15722
rect 1144 15695 4700 15706
rect 4780 15695 4814 15839
rect 5300 15811 5381 15858
rect 5060 15780 5116 15808
rect 4820 15778 5116 15780
rect 4820 15722 5116 15752
rect 5347 15708 5381 15811
rect 5300 15695 5381 15708
rect 5449 15706 5483 16319
rect 6192 16291 6320 16338
rect 6239 15723 6320 16291
rect 5446 15695 6191 15706
rect -1796 15661 6191 15695
rect 4666 15581 4700 15661
rect 4780 15581 4814 15661
rect 5347 15581 5381 15661
rect 5449 15581 5483 15661
rect 6341 15581 6375 18201
rect 7840 17894 7872 18316
rect 7878 17932 7910 18278
rect 9879 17861 9913 18666
rect 9981 18661 10015 18666
rect 10602 18660 10616 18666
rect 10816 18660 10880 18666
rect 9981 18645 10015 18654
rect 10588 18652 10602 18660
rect 10616 18652 10658 18660
rect 10118 18645 10738 18652
rect 10884 18645 11258 18666
rect 13670 18660 13938 18666
rect 10062 18639 13942 18645
rect 10062 18633 13966 18639
rect 14068 18633 14102 18691
rect 16704 18633 16738 18691
rect 16759 18668 16840 18691
rect 16887 18690 18245 18691
rect 19470 18690 19526 18694
rect 20714 18690 20770 18694
rect 18062 18684 18159 18690
rect 16806 18652 16840 18668
rect 16859 18662 17756 18684
rect 16778 18633 17234 18652
rect 18103 18649 18149 18684
rect 18109 18645 18143 18649
rect 18050 18633 18061 18644
rect 10058 18632 18061 18633
rect 9976 18618 10049 18620
rect 10062 18619 18061 18632
rect 18075 18621 18177 18638
rect 9934 18571 10062 18618
rect 10074 18577 18061 18619
rect 9981 17981 10062 18571
rect 10118 18230 10738 18577
rect 10788 18282 10822 18577
rect 10896 18509 10930 18577
rect 11159 18524 11170 18535
rect 10843 18496 10943 18509
rect 10843 18462 10958 18496
rect 10983 18490 11170 18524
rect 11171 18462 11252 18509
rect 10884 18424 10958 18462
rect 11218 18424 11252 18462
rect 10884 18408 10942 18424
rect 10896 18282 10930 18408
rect 11159 18396 11170 18407
rect 10983 18362 11170 18396
rect 11320 18282 11354 18577
rect 13954 18382 13988 18577
rect 14068 18382 14102 18577
rect 10788 18248 11354 18282
rect 13796 18372 14244 18382
rect 10118 17986 10738 18176
rect 10896 18162 10930 18248
rect 13796 18170 14252 18372
rect 10788 18128 11354 18162
rect 13804 18160 14252 18170
rect 10788 18054 10822 18128
rect 10788 18046 10890 18054
rect 10896 18046 10930 18128
rect 11159 18048 11170 18059
rect 10788 18016 10828 18046
rect 10896 18033 10936 18046
rect 10843 18026 10943 18033
rect 10836 18020 10943 18026
rect 10836 18016 10958 18020
rect 10778 18002 10786 18008
rect 10036 17975 10053 17981
rect 10063 17975 10738 17986
rect 10788 17996 10822 18016
rect 10843 17996 10958 18016
rect 10983 18014 11170 18048
rect 11171 17996 11252 18033
rect 11320 17996 11354 18128
rect 10788 17986 11444 17996
rect 10788 17975 11544 17986
rect 13954 17975 13988 18160
rect 14068 17975 14102 18160
rect 16704 17975 16738 18577
rect 16740 18562 17196 18577
rect 18062 18571 18143 18618
rect 16806 18100 16840 18562
rect 18109 18084 18143 18571
rect 18062 18072 18159 18084
rect 18211 18072 18245 18690
rect 19470 18634 19526 18638
rect 20714 18634 20770 18638
rect 19470 18132 19526 18134
rect 20714 18132 20770 18134
rect 19470 18076 19526 18078
rect 20714 18076 20770 18078
rect 16759 18050 16840 18057
rect 16759 18046 16874 18050
rect 16759 18022 16840 18046
rect 16899 18038 20160 18072
rect 18062 18037 18159 18038
rect 16887 18032 18159 18037
rect 17716 18026 18159 18032
rect 16759 18010 16846 18022
rect 17716 18020 18143 18026
rect 16800 17990 16846 18010
rect 16806 17987 16846 17990
rect 16790 17981 16887 17987
rect 16790 17976 17716 17981
rect 16790 17975 16887 17976
rect 18050 17975 18061 17986
rect 10036 17938 18061 17975
rect 18103 17981 18143 18020
rect 18103 17974 18118 17981
rect 9934 17891 10062 17938
rect 10074 17919 18061 17938
rect 9981 17874 10062 17891
rect 9934 17861 10062 17874
rect 10118 17861 10738 17919
rect 10770 17898 11424 17919
rect 13941 17907 13942 17908
rect 13942 17906 13943 17907
rect 10788 17861 10822 17898
rect 10896 17882 10930 17898
rect 10983 17895 11170 17898
rect 10967 17886 11175 17895
rect 10896 17864 10936 17882
rect 11194 17870 11250 17898
rect 11166 17864 11250 17870
rect 10896 17861 10930 17864
rect 11320 17861 11354 17898
rect 13954 17861 13988 17919
rect 14068 17861 14102 17919
rect 16704 17861 16738 17919
rect 16790 17907 16887 17919
rect 16806 17861 16840 17907
rect 18062 17891 18143 17938
rect 18109 17874 18143 17891
rect 18062 17861 18143 17874
rect 18211 17861 18245 18038
rect 9879 17827 18245 17861
rect -1991 15547 6375 15581
rect 4666 15328 4700 15547
rect -2794 15304 -2787 15328
rect -2741 15304 4774 15328
rect 4666 15215 4700 15304
rect 4780 15215 4814 15547
rect 4820 15304 5116 15328
rect 5060 15248 5116 15272
rect 5347 15243 5381 15547
rect 4825 15227 4826 15228
rect 4826 15226 4827 15227
rect 5288 15215 5299 15226
rect 4632 15181 5299 15215
rect 4666 14649 4700 15181
rect 4780 14649 4814 15181
rect 4826 15169 4827 15170
rect 4825 15168 4826 15169
rect 5300 15153 5381 15200
rect 5347 14649 5381 15153
rect 5449 14649 5483 15547
rect 7840 15240 7872 15662
rect 7878 15278 7910 15624
rect 9879 15207 9913 17827
rect 9981 17406 10062 17827
rect 10118 17754 10738 17827
rect 10788 17806 10822 17827
rect 10896 17806 10930 17827
rect 10936 17826 10970 17827
rect 11166 17808 11250 17827
rect 11320 17806 11354 17827
rect 10788 17772 11354 17806
rect 9981 17388 10015 17406
rect 10896 17388 10930 17772
rect 13954 17736 13988 17827
rect 14068 17736 14102 17827
rect 13796 17524 14244 17736
rect 13828 17388 14104 17524
rect 16704 17396 16738 17827
rect 16806 17442 16840 17827
rect 18109 17427 18143 17827
rect 18062 17426 18143 17427
rect 18062 17414 18159 17426
rect 16899 17396 18159 17414
rect 16434 17394 16800 17396
rect 16846 17394 18159 17396
rect 16704 17388 16738 17394
rect 16887 17388 18159 17394
rect 18211 17388 18245 17827
rect 19470 17468 19526 17476
rect 20714 17468 20770 17476
rect 19470 17412 19526 17420
rect 20714 17412 20770 17420
rect 9976 17280 18396 17388
rect 19470 17374 19526 17382
rect 20714 17374 20880 17402
rect 19470 17318 19526 17326
rect 20714 17318 20770 17346
rect 9934 17233 18396 17280
rect 9976 16622 18396 17233
rect 9934 16575 18396 16622
rect 9976 16572 18396 16575
rect 9976 15964 18281 16572
rect 9934 15917 18281 15964
rect 9976 15207 18281 15917
rect 9879 15173 18281 15207
rect -2808 14638 5483 14649
rect -2797 14626 5483 14638
rect -2808 14615 5483 14626
rect -2781 14569 -2747 14615
rect -2398 14578 -996 14594
rect -1992 14557 -1338 14578
rect 4666 14557 4700 14615
rect 4780 14557 4814 14615
rect 4825 14569 4826 14570
rect 5347 14569 5381 14615
rect 4826 14568 4827 14569
rect 5288 14557 5299 14568
rect -2688 14501 5299 14557
rect -2781 13905 -2747 14495
rect -1972 14480 -1318 14501
rect 1042 14306 1490 14316
rect 1034 14104 1490 14306
rect 1034 14094 1482 14104
rect 4058 13914 4464 14292
rect 3978 13910 4464 13914
rect 4666 13910 4700 14501
rect 1144 13899 4700 13910
rect 4780 13899 4814 14501
rect 5300 14495 5381 14542
rect 5288 13899 5299 13910
rect 5347 13905 5381 14495
rect -2688 13843 5299 13899
rect 4016 13824 4472 13843
rect -2781 13815 -2747 13819
rect 4058 13785 4464 13824
rect 4666 13785 4700 13843
rect 4780 13785 4814 13843
rect 4826 13831 4827 13832
rect 4825 13830 4826 13831
rect 5300 13815 5381 13862
rect 5347 13798 5381 13815
rect 5300 13785 5381 13798
rect 5449 13785 5483 14615
rect -2819 13751 5483 13785
rect 1258 13640 1390 13650
rect 1034 13428 1482 13640
rect 4666 13219 4700 13751
rect 4780 13219 4814 13751
rect 5347 13247 5381 13751
rect 4825 13231 4826 13232
rect 4826 13230 4827 13231
rect 5288 13219 5299 13230
rect 4632 13185 5299 13219
rect -274 13082 36 13088
rect 722 12994 1342 13088
rect 1392 13040 1958 13074
rect 1392 12994 1426 13040
rect 722 12945 1490 12994
rect 1576 12960 1774 12971
rect 722 12860 1575 12945
rect 1587 12926 1774 12960
rect 1775 12898 1903 12945
rect 1822 12860 1903 12898
rect 722 12834 1518 12860
rect 722 12782 1490 12834
rect 1576 12832 1774 12843
rect 1587 12798 1774 12832
rect 722 12666 1342 12782
rect 1392 12718 1426 12782
rect 1924 12718 1958 13040
rect 1392 12684 1958 12718
rect 4666 12666 4700 13185
rect 4780 12666 4814 13185
rect 4826 13173 4827 13174
rect 4825 13172 4826 13173
rect 5300 13157 5381 13204
rect 3592 12650 5056 12666
rect -2700 12521 580 12538
rect 2148 12521 3648 12540
rect 4666 12470 4700 12650
rect 4774 12619 4820 12650
rect 5300 12619 5301 12620
rect 5347 12619 5381 13157
rect 5299 12618 5300 12619
rect 4746 12595 4848 12610
rect 4746 12591 5322 12595
rect 4842 12573 5322 12591
rect 5347 12573 5381 12610
rect 4826 12572 5322 12573
rect 4826 12557 5300 12572
rect 5309 12557 5419 12572
rect 4826 12540 5439 12557
rect 5449 12540 5483 13751
rect 9976 15137 18281 15173
rect 9976 14698 14138 15137
rect 9976 14687 18285 14698
rect 9976 14675 18274 14687
rect 9976 14664 18285 14675
rect 9976 14606 14138 14664
rect 16786 14618 17244 14638
rect 18224 14618 18258 14664
rect 16746 14606 17244 14618
rect 9976 14560 18174 14606
rect 9976 14550 18185 14560
rect 9976 14370 14138 14550
rect 16746 14546 17244 14550
rect 16746 14526 17204 14546
rect 16490 14502 17594 14522
rect 16462 14474 17622 14494
rect 9976 14158 14334 14370
rect 9976 14130 14316 14158
rect 9976 13948 14138 14130
rect 18174 13948 18185 13959
rect 18224 13954 18258 14544
rect 9976 13938 18185 13948
rect 9976 13892 18174 13938
rect 9976 13834 14138 13892
rect 18224 13864 18258 13868
rect 9976 13800 18292 13834
rect 9976 13698 14138 13800
rect 9976 13486 14328 13698
rect 9976 13330 14138 13486
rect 9976 13296 14178 13330
rect 9976 13268 14138 13296
rect 14144 13268 14178 13296
rect 9976 13262 14178 13268
rect 9976 13230 14138 13262
rect 14144 13230 14178 13262
rect 9976 13228 14178 13230
rect 9976 13014 14138 13228
rect 14144 13014 14178 13228
rect 9976 12980 14178 13014
rect 9976 12571 14138 12980
rect 14228 12922 14866 13384
rect 4826 12530 5483 12540
rect 6708 12530 6764 12540
rect 4826 12522 5439 12530
rect 5000 12521 5300 12522
rect 5285 12515 5300 12521
rect 5347 12511 5381 12515
rect 5341 12484 5387 12511
rect 5449 12484 5483 12530
rect 9699 12500 14138 12571
rect 5300 12474 6764 12484
rect 5449 12470 5483 12474
rect 9699 12470 14262 12500
rect 4666 12436 14262 12470
rect 5449 12268 5483 12436
rect 9699 12400 14262 12436
rect 14130 12382 14262 12400
rect 13882 12317 14330 12382
rect 18326 12317 18360 16572
rect -2896 11061 5519 12268
rect 9976 11110 18391 12317
rect -2860 8570 -2826 11061
rect 1010 10996 1458 11061
rect 1258 10878 1390 10996
rect -2384 10830 -982 10844
rect 3916 10806 5336 10836
rect 5352 10814 5386 10853
rect 5454 10806 5488 11061
rect 10172 10842 13452 10857
rect 15020 10842 16520 10857
rect 17872 10842 18172 10857
rect 9953 10806 18391 10842
rect 3820 10772 18391 10806
rect -334 10458 60 10494
rect -274 10398 36 10434
rect 758 10364 1306 10398
rect 758 10082 792 10364
rect 1120 10284 1131 10295
rect 822 10240 894 10278
rect 944 10250 1131 10284
rect 1132 10240 1204 10278
rect 860 10206 894 10240
rect 904 10228 1160 10230
rect 1120 10202 1131 10207
rect 1170 10206 1204 10240
rect 932 10200 1132 10202
rect 1120 10196 1131 10200
rect 944 10178 1131 10196
rect 928 10162 1136 10178
rect 1166 10176 1256 10178
rect 932 10156 934 10162
rect 1128 10156 1132 10162
rect 1272 10150 1306 10364
rect 904 10144 934 10150
rect 1128 10148 1306 10150
rect 1128 10144 1160 10148
rect 894 10128 1170 10144
rect 906 10124 1158 10128
rect 1272 10116 1306 10148
rect 798 10110 1306 10116
rect 1272 10082 1306 10110
rect 758 10048 1306 10082
rect 1356 9994 1994 10456
rect 3820 10144 3854 10772
rect 5352 10744 5386 10756
rect 4664 10704 4702 10742
rect 5318 10710 5338 10716
rect 5346 10710 5386 10744
rect 5352 10704 5386 10710
rect 3996 10670 4702 10704
rect 4754 10670 5438 10704
rect 5313 10632 5314 10633
rect 5314 10631 5315 10632
rect 3923 10620 3968 10631
rect 4681 10620 4726 10631
rect 3934 10144 3968 10620
rect 3979 10156 3980 10157
rect 4680 10156 4681 10157
rect 3980 10155 3981 10156
rect 4679 10155 4680 10156
rect 4692 10144 4726 10620
rect 5352 10228 5386 10670
rect 5416 10228 5424 10660
rect 4737 10156 4738 10157
rect 4738 10155 4739 10156
rect 5302 10144 5313 10155
rect 3786 10110 5313 10144
rect 5318 10132 5338 10228
rect 5346 10172 5386 10228
rect 5444 10200 5452 10632
rect 5346 10160 5366 10172
rect 5318 10120 5338 10122
rect 1008 9680 1456 9892
rect 3820 9578 3854 10110
rect 3934 9578 3968 10110
rect 3980 10098 3981 10099
rect 4679 10098 4680 10099
rect 3979 10097 3980 10098
rect 4680 10097 4681 10098
rect 4692 9578 4726 10110
rect 4738 10098 4739 10099
rect 4737 10097 4738 10098
rect 5314 10082 5386 10120
rect 5318 10012 5338 10082
rect 5346 10012 5386 10082
rect 5352 9578 5386 10012
rect 5454 9578 5488 10772
rect 5496 10670 5535 10704
rect -2785 9567 5488 9578
rect -2774 9555 5488 9567
rect -2785 9544 5488 9555
rect -2758 9498 -2724 9544
rect -1992 9486 -1338 9504
rect 3820 9486 3854 9544
rect 3934 9486 3968 9544
rect 3979 9498 3980 9499
rect 4680 9498 4681 9499
rect 3980 9497 3981 9498
rect 4679 9497 4680 9498
rect 4692 9486 4726 9544
rect 4737 9498 4738 9499
rect 4738 9497 4739 9498
rect 5302 9486 5313 9497
rect -2674 9430 5313 9486
rect 5318 9474 5338 9544
rect 5346 9502 5386 9544
rect 5352 9498 5386 9502
rect 5318 9462 5338 9464
rect -2758 8834 -2724 9424
rect -1956 9406 -1302 9430
rect 996 9220 1444 9248
rect 996 9036 1462 9220
rect 1014 9008 1462 9036
rect 3820 8904 3854 9430
rect 3590 8884 3928 8904
rect 3820 8876 3854 8884
rect 3618 8856 3928 8876
rect 3820 8828 3854 8856
rect 3934 8852 3968 9430
rect 3974 8884 4076 8904
rect 4580 8884 4686 8904
rect 3974 8856 4076 8876
rect 4580 8856 4686 8876
rect 3874 8832 4332 8852
rect 3874 8828 4372 8832
rect 4692 8828 4726 9430
rect 5314 9424 5386 9462
rect 5318 9360 5338 9424
rect 5346 9360 5386 9424
rect 5444 9360 5446 9388
rect 5352 8884 5386 9360
rect 5416 9332 5418 9360
rect 5416 8884 5424 9332
rect 5302 8828 5313 8839
rect -2674 8772 5313 8828
rect 5318 8794 5338 8884
rect 5346 8834 5386 8884
rect 5444 8856 5452 9360
rect 5346 8822 5366 8834
rect 5318 8782 5338 8784
rect 2930 8766 3186 8772
rect -2758 8714 -2724 8748
rect 2958 8738 3158 8752
rect 3820 8714 3854 8772
rect 3874 8760 4372 8772
rect 4679 8760 4680 8761
rect 3914 8740 4372 8760
rect 4680 8759 4681 8760
rect 3934 8714 3968 8740
rect 4692 8714 4726 8772
rect 4738 8760 4739 8761
rect 4737 8759 4738 8760
rect 5314 8744 5386 8782
rect 5318 8718 5338 8744
rect 5346 8718 5386 8744
rect 5314 8714 5386 8718
rect 5454 8714 5488 9544
rect -2805 8680 5488 8714
rect -2758 8570 -2724 8680
rect -2860 8484 -2724 8570
rect -2860 8086 -2826 8484
rect -2758 8180 -2724 8484
rect -2718 8208 -2170 8242
rect -2718 8180 -2684 8208
rect -2204 8180 -2170 8208
rect -2764 8164 -2684 8180
rect -2718 8152 -2684 8164
rect -2792 8136 -2684 8152
rect -2238 8148 -2136 8180
rect -2120 8166 -1482 8296
rect -2120 8148 -1330 8166
rect 2930 8154 2944 8232
rect 2958 8154 2972 8232
rect 3820 8148 3854 8680
rect 3934 8148 3968 8680
rect 3979 8160 3980 8161
rect 4680 8160 4681 8161
rect 3980 8159 3981 8160
rect 4679 8159 4680 8160
rect 4692 8148 4726 8680
rect 5352 8232 5386 8680
rect 5416 8232 5428 8680
rect 4737 8160 4738 8161
rect 4738 8159 4739 8160
rect 5302 8148 5313 8159
rect -2860 8008 -2724 8086
rect -2860 7041 -2826 8008
rect -2758 7518 -2724 8008
rect -2718 7926 -2684 8136
rect -2674 8114 -2170 8148
rect -2654 8084 -2582 8114
rect -2532 8102 -2356 8114
rect -2532 8094 -2345 8102
rect -2344 8084 -2272 8114
rect -2616 8050 -2582 8084
rect -2356 8040 -2345 8051
rect -2306 8050 -2272 8084
rect -2532 8006 -2345 8040
rect -2314 8030 -2310 8050
rect -2342 8002 -2310 8022
rect -2204 7926 -2170 8114
rect -2718 7892 -2170 7926
rect -2120 8114 0 8148
rect 3786 8114 5313 8148
rect 5318 8136 5338 8232
rect 5346 8176 5386 8232
rect 5444 8204 5488 8680
rect 5346 8164 5366 8176
rect 5318 8124 5338 8126
rect -2120 8092 -1330 8114
rect -2120 7834 -1482 8092
rect -2718 7732 -2170 7766
rect -2718 7450 -2684 7732
rect -2356 7652 -2345 7663
rect -2654 7608 -2582 7646
rect -2532 7618 -2345 7652
rect -2344 7608 -2272 7646
rect -2616 7574 -2582 7608
rect -2572 7574 -2316 7598
rect -2306 7574 -2272 7608
rect -2356 7570 -2345 7574
rect -2544 7546 -2344 7570
rect -2532 7530 -2345 7546
rect -2204 7484 -2170 7732
rect -2678 7456 -2170 7484
rect -2204 7450 -2170 7456
rect -2718 7416 -2170 7450
rect -2120 7358 -1482 7820
rect 3820 7490 3854 8114
rect 3934 7490 3968 8114
rect 3980 8102 3981 8103
rect 4679 8102 4680 8103
rect 3979 8101 3980 8102
rect 4680 8101 4681 8102
rect 3979 7502 3980 7503
rect 4680 7502 4681 7503
rect 3980 7501 3981 7502
rect 4679 7501 4680 7502
rect 4692 7490 4726 8114
rect 4738 8102 4739 8103
rect 4737 8101 4738 8102
rect 5314 8086 5386 8124
rect 5318 8022 5338 8086
rect 5346 8022 5386 8086
rect 5352 7574 5386 8022
rect 5416 7674 5424 8022
rect 5444 7674 5452 8050
rect 4737 7502 4738 7503
rect 4738 7501 4739 7502
rect 5302 7490 5313 7501
rect 3786 7456 5313 7490
rect 5318 7478 5338 7574
rect 5346 7518 5392 7574
rect 5346 7506 5366 7518
rect 5380 7506 5392 7518
rect 5408 7478 5420 7574
rect 5318 7466 5338 7468
rect 3820 7041 3854 7456
rect 3934 7041 3968 7456
rect 3980 7444 3981 7445
rect 4679 7444 4680 7445
rect 3979 7443 3980 7444
rect 4680 7443 4681 7444
rect 4692 7041 4726 7456
rect 4738 7444 4739 7445
rect 4737 7443 4738 7444
rect 5314 7440 5386 7466
rect 5314 7428 5392 7440
rect 5318 7358 5338 7428
rect 5346 7358 5392 7428
rect 5408 7358 5420 7468
rect 5352 7041 5386 7358
rect -2896 7010 5419 7041
rect -11460 5302 -6760 5336
rect -11460 5234 -9022 5302
rect -8794 5234 -8760 5302
rect -8566 5272 -8532 5302
rect -8692 5234 -8434 5272
rect -8222 5265 -8184 5272
rect -8108 5268 -8074 5302
rect -8222 5250 -8176 5265
rect -8234 5234 -8176 5250
rect -11460 5200 -8176 5234
rect -8172 5200 -8140 5234
rect -11460 4806 -9022 5200
rect -8794 5184 -8760 5200
rect -8820 5161 -8760 5184
rect -8692 5162 -8634 5200
rect -8820 5150 -8741 5161
rect -8794 4806 -8726 5150
rect -8702 4806 -8690 4812
rect -8680 4806 -8635 5162
rect -12120 4770 -8594 4806
rect -12182 4736 -8594 4770
rect -12182 3156 -12148 4736
rect -12120 4408 -8594 4736
rect -8566 4408 -8532 5200
rect -8234 5162 -8176 5200
rect -8138 5184 -8074 5268
rect -8138 5166 -8060 5184
rect -8222 4596 -8188 5162
rect -8222 4422 -8182 4596
rect -8222 4420 -8177 4422
rect -8196 4408 -8182 4420
rect -12120 4336 -8212 4408
rect -8168 4380 -8154 4568
rect -12120 4268 -8594 4336
rect -8566 4268 -8532 4336
rect -8108 4330 -8060 5166
rect -8108 4268 -8074 4330
rect -12120 4234 -8074 4268
rect -12120 3536 -8594 4234
rect -8566 3536 -8532 4234
rect -12120 3502 -8532 3536
rect -12120 3156 -8594 3502
rect -8566 3402 -8532 3502
rect -13857 3122 -8594 3156
rect -13857 3104 -13782 3122
rect -13857 3074 -13823 3104
rect -13857 2718 -13817 3074
rect -13816 3018 -13782 3104
rect -13751 3104 -13706 3122
rect -13816 2718 -13761 3018
rect -13751 2718 -13717 3104
rect -13637 3054 -13603 3122
rect -12541 3101 -12507 3122
rect -12182 3114 -12148 3122
rect -12120 3114 -8594 3122
rect -13199 3070 -13152 3101
rect -13211 3054 -13152 3070
rect -13072 3054 -13025 3101
rect -12541 3070 -12494 3101
rect -12553 3054 -12494 3070
rect -12414 3054 -12367 3101
rect -12182 3064 -8594 3114
rect -12182 3058 -12148 3064
rect -12120 3058 -8594 3064
rect -12182 3054 -8594 3058
rect -13656 3020 -13025 3054
rect -12982 3020 -12367 3054
rect -12324 3020 -8594 3054
rect -13702 2972 -13683 2977
rect -13671 2972 -13668 2977
rect -13713 2961 -13668 2972
rect -13702 2718 -13668 2961
rect -13637 2718 -13603 3020
rect -13211 2973 -13153 3020
rect -13199 2718 -13165 2973
rect -13122 2968 -13112 3014
rect -13066 2968 -13056 3014
rect -12553 2973 -12495 3020
rect -13078 2776 -13056 2968
rect -13055 2961 -13010 2972
rect -13122 2718 -13112 2776
rect -13066 2718 -13056 2776
rect -13044 2718 -13010 2961
rect -12541 2718 -12507 2973
rect -12470 2718 -12450 3014
rect -12414 2972 -12394 3014
rect -12182 3008 -8594 3020
rect -12414 2961 -12352 2972
rect -12414 2718 -12394 2961
rect -12386 2718 -12352 2961
rect -18364 2713 -12220 2718
rect -27189 918 -27144 2692
rect -27128 1676 -27100 2158
rect -27128 1476 -27084 1676
rect -27128 918 -27100 1476
rect -27072 1448 -27056 1704
rect -27007 918 -26962 2692
rect -26531 918 -26486 2692
rect -26468 2426 -12220 2713
rect -12182 2426 -12148 3008
rect -12120 2426 -8594 3008
rect -8586 2534 -6628 3402
rect -6526 3268 -6512 3634
rect -6486 2994 -6470 3180
rect -5804 3160 -5770 3194
rect -5690 3160 -5656 3270
rect -5038 3160 -5004 3274
rect -3494 3238 -3460 3274
rect -4924 3160 -4890 3194
rect -4266 3160 -4232 3194
rect -3852 3160 -3460 3238
rect -2983 3272 -2949 6909
rect -2896 6860 5424 7010
rect -2896 6820 5420 6860
rect -2896 6810 5419 6820
rect -2896 6808 5420 6810
rect -2896 6202 5424 6808
rect 5444 6230 5446 6284
rect -2896 6060 5419 6202
rect 5454 6084 5488 8204
rect 5444 6060 5490 6084
rect 5496 6060 5514 6120
rect 6202 6060 6248 6084
rect -2896 6026 5488 6060
rect 7852 6032 7864 6084
rect 9953 6039 18391 10772
rect 19202 10768 19402 10770
rect 21312 10668 27232 20668
rect 27272 20628 27273 20629
rect 27271 20627 27272 20628
rect 21258 10664 27232 10668
rect 21312 10535 27232 10664
rect 19263 10504 27232 10535
rect 27520 20616 27598 22622
rect 27701 22218 27749 26373
rect 27829 26383 27863 26435
rect 28487 26414 28521 26435
rect 28445 26383 28521 26414
rect 28544 26414 28555 26432
rect 29145 26414 29179 26435
rect 29803 26414 29837 26435
rect 30066 26414 30278 26435
rect 30461 26414 30495 26435
rect 31119 26414 31153 26435
rect 27829 26286 27875 26383
rect 28445 26367 28533 26383
rect 28544 26367 31153 26414
rect 31232 26373 31303 26762
rect 27877 26340 28533 26367
rect 28535 26340 29191 26367
rect 27877 26333 29191 26340
rect 29193 26340 29849 26367
rect 29851 26340 30507 26367
rect 29193 26333 30507 26340
rect 30509 26333 31153 26367
rect 27904 26327 27932 26333
rect 28394 26327 28457 26333
rect 28481 26299 28485 26333
rect 28487 26327 28590 26333
rect 29052 26327 29104 26333
rect 28487 26286 28533 26327
rect 27829 26274 27863 26286
rect 28462 26274 28475 26285
rect 28487 26274 28521 26286
rect 27815 25630 27863 26274
rect 28473 25630 28521 26274
rect 28544 25630 28555 26327
rect 29145 26286 29191 26333
rect 29212 26327 29252 26333
rect 29714 26327 29773 26333
rect 29797 26299 29801 26333
rect 29803 26327 29922 26333
rect 29803 26286 29849 26327
rect 29120 26274 29133 26285
rect 29145 26274 29190 26286
rect 29778 26274 29791 26285
rect 29803 26274 29848 26286
rect 27815 24958 27874 25630
rect 28473 24958 28532 25630
rect 29131 24958 29190 26274
rect 29712 24958 29714 25096
rect 29740 24958 29742 25096
rect 29789 24958 29848 26274
rect 30066 26106 30278 26333
rect 30384 26327 30424 26333
rect 30461 26286 30507 26333
rect 30532 26327 30574 26333
rect 31036 26327 31089 26333
rect 31113 26299 31117 26333
rect 30436 26274 30449 26285
rect 30461 26274 30506 26286
rect 31094 26274 31107 26285
rect 31119 26274 31153 26333
rect 30052 25782 30392 26106
rect 30447 24958 30506 26274
rect 31034 24958 31036 25096
rect 31062 24958 31064 25096
rect 31105 24958 31153 26274
rect 27815 24911 31153 24958
rect 27815 24809 27874 24911
rect 27879 24877 28532 24911
rect 28549 24877 29190 24911
rect 27879 24871 27897 24877
rect 28461 24861 28532 24877
rect 29119 24861 29190 24877
rect 29195 24877 29848 24911
rect 29865 24877 30506 24911
rect 29195 24871 29213 24877
rect 28473 24809 28532 24861
rect 29131 24809 29190 24861
rect 29712 24809 29714 24871
rect 29740 24809 29742 24871
rect 29777 24861 29848 24877
rect 30435 24861 30506 24877
rect 30511 24877 31153 24911
rect 30511 24871 30529 24877
rect 29789 24809 29848 24861
rect 30447 24809 30506 24861
rect 31034 24809 31036 24871
rect 31062 24809 31064 24871
rect 31093 24861 31153 24877
rect 31105 24809 31153 24861
rect 31186 24809 31190 25016
rect 27803 24775 31190 24809
rect 27815 23815 27874 24775
rect 28473 23815 28532 24775
rect 29131 23815 29190 24775
rect 29712 24606 29714 24775
rect 29740 24634 29742 24775
rect 29789 23815 29848 24775
rect 30447 23815 30506 24775
rect 31034 24576 31036 24775
rect 31062 24604 31064 24775
rect 31105 23815 31153 24775
rect 31186 24604 31190 24775
rect 27803 23781 31187 23815
rect 27815 23778 27874 23781
rect 28473 23778 28532 23781
rect 27815 23713 27863 23778
rect 28473 23760 28521 23778
rect 28445 23713 28521 23760
rect 28544 23760 28555 23778
rect 29131 23760 29190 23781
rect 29789 23760 29848 23781
rect 30447 23760 30506 23781
rect 31105 23760 31153 23781
rect 28544 23713 31153 23760
rect 27815 23679 27874 23713
rect 27877 23679 28532 23713
rect 28535 23679 29190 23713
rect 29193 23679 29848 23713
rect 29851 23679 30506 23713
rect 30509 23679 31153 23713
rect 27815 22316 27863 23679
rect 28473 22316 28521 23679
rect 27815 22218 27849 22316
rect 28473 22304 28507 22316
rect 28510 22304 28521 22316
rect 28544 22304 28555 23679
rect 29131 22316 29190 23679
rect 29131 22304 29165 22316
rect 29712 22304 29714 23242
rect 29740 22304 29742 23242
rect 29789 22316 29848 23679
rect 30447 22316 30506 23679
rect 29789 22304 29823 22316
rect 30447 22304 30481 22316
rect 31034 22304 31036 23242
rect 31062 22304 31064 23242
rect 31105 22316 31153 23679
rect 31219 23538 31303 26373
rect 31382 24552 31416 27248
rect 31500 26418 31526 26424
rect 31528 26418 31554 26452
rect 31908 26360 32370 26998
rect 32786 26474 32820 27248
rect 32898 26474 32934 27248
rect 32944 26474 32945 27248
rect 33558 26952 33592 27248
rect 33556 26686 33598 26952
rect 33556 26572 33603 26686
rect 33612 26628 33626 26952
rect 33656 26686 33690 27248
rect 33558 26474 33603 26572
rect 33656 26474 33701 26686
rect 34216 26474 34261 27248
rect 34286 26474 34322 26952
rect 34342 26474 34378 26952
rect 34414 26474 34459 27248
rect 34874 26474 34919 27248
rect 35172 26474 35217 27248
rect 35532 26686 35566 27248
rect 35930 26686 35964 27248
rect 36190 26686 36224 27248
rect 35532 26474 35577 26686
rect 35930 26474 35975 26686
rect 36190 26474 36235 26686
rect 36304 26474 36338 27248
rect 38962 26505 38996 27248
rect 32772 26440 36338 26474
rect 31966 26276 32316 26310
rect 31966 25824 32000 26276
rect 32086 26242 32178 26246
rect 32086 26208 32192 26242
rect 32124 26174 32192 26208
rect 32128 26136 32174 26174
rect 32069 26124 32125 26135
rect 32080 25948 32125 26124
rect 32140 26124 32174 26136
rect 32186 26124 32213 26135
rect 32140 25948 32213 26124
rect 32140 25936 32174 25948
rect 32086 25932 32178 25936
rect 32086 25898 32192 25932
rect 32124 25864 32192 25898
rect 32128 25848 32174 25864
rect 32282 25824 32316 26276
rect 32772 25824 32820 26440
rect 32898 26410 32934 26440
rect 32944 26410 32945 26440
rect 33144 26410 33356 26440
rect 33558 26410 33603 26440
rect 33656 26410 33701 26440
rect 33810 26410 34022 26440
rect 34216 26410 34261 26440
rect 34272 26410 34322 26440
rect 34342 26410 34378 26440
rect 34414 26410 34670 26440
rect 34874 26410 34919 26440
rect 35172 26410 35217 26440
rect 35532 26410 35577 26440
rect 35930 26410 35975 26440
rect 32898 26372 33554 26410
rect 32898 26332 32945 26372
rect 32948 26338 33554 26372
rect 33558 26372 34212 26410
rect 33558 26340 33603 26372
rect 33606 26340 34212 26372
rect 33558 26338 34212 26340
rect 34216 26372 34870 26410
rect 32972 26332 32994 26338
rect 32875 26288 32886 26299
rect 32898 26288 32972 26332
rect 32886 26284 32972 26288
rect 32994 26284 33000 26332
rect 32886 25824 32945 26284
rect 33144 26186 33356 26338
rect 33558 26332 33702 26338
rect 33558 26299 33603 26332
rect 33644 26300 33702 26332
rect 33533 26288 33603 26299
rect 33544 26284 33603 26288
rect 33650 26284 33654 26300
rect 33544 26276 33650 26284
rect 33122 25824 33444 26186
rect 33544 25824 33603 26276
rect 33656 25824 33701 26300
rect 33810 26186 34022 26338
rect 34216 26328 34261 26372
rect 34264 26338 34870 26372
rect 34874 26372 35528 26410
rect 34322 26332 34328 26338
rect 34272 26328 34322 26332
rect 34198 26299 34322 26328
rect 34191 26288 34322 26299
rect 34198 26284 34322 26288
rect 34328 26284 34378 26332
rect 34402 26300 34670 26338
rect 34198 26186 34272 26284
rect 34322 26276 34328 26284
rect 33810 26014 34272 26186
rect 33912 25824 34272 26014
rect 34414 26198 34670 26300
rect 34874 26299 34919 26372
rect 34922 26338 35528 26372
rect 35532 26372 36186 26410
rect 35160 26300 35218 26338
rect 35532 26320 35577 26372
rect 35580 26338 36186 26372
rect 34849 26288 34919 26299
rect 34860 26198 34919 26288
rect 34414 26018 34960 26198
rect 34414 25824 34459 26018
rect 34638 25824 34960 26018
rect 35172 25824 35217 26300
rect 35514 26299 35588 26320
rect 35918 26300 35976 26338
rect 35507 26288 35588 26299
rect 35514 26220 35588 26288
rect 35384 25824 35706 26220
rect 35930 25824 35975 26300
rect 36190 26299 36235 26440
rect 36165 26288 36235 26299
rect 36176 25824 36235 26288
rect 36290 25824 36338 26440
rect 36421 25824 40045 26505
rect 41494 25824 41522 26508
rect 42762 26474 42786 27248
rect 42796 26474 42820 27248
rect 44575 26474 53013 27248
rect 31966 25762 41522 25824
rect 31994 25754 41522 25762
rect 41528 26440 53013 26474
rect 31338 24530 31458 24552
rect 31338 24404 31750 24530
rect 31344 24000 31750 24404
rect 31382 23690 31416 24000
rect 31994 23538 41502 25754
rect 41528 23820 41562 26440
rect 42762 26410 42786 26440
rect 42796 26410 42820 26440
rect 44268 26410 44302 26440
rect 44575 26410 53013 26440
rect 41994 26388 42032 26410
rect 41982 26372 42040 26388
rect 42272 26372 42310 26410
rect 42752 26388 42790 26410
rect 42796 26388 42968 26410
rect 42740 26372 42968 26388
rect 42982 26372 43626 26410
rect 43640 26372 53013 26410
rect 41704 26338 42310 26372
rect 42362 26338 42968 26372
rect 43020 26338 43626 26372
rect 41982 26300 42040 26338
rect 42740 26300 42820 26338
rect 43498 26332 43600 26338
rect 43666 26332 43672 26340
rect 43678 26338 44308 26372
rect 44196 26332 44308 26338
rect 44324 26338 53013 26372
rect 44324 26332 44400 26338
rect 43498 26300 43556 26332
rect 41631 26288 41676 26299
rect 41642 23820 41676 26288
rect 41994 23820 42028 26300
rect 42289 26288 42334 26299
rect 42300 23820 42334 26288
rect 42752 23820 42786 26300
rect 42796 25188 42820 26300
rect 42947 26288 43003 26299
rect 42958 25188 43003 26288
rect 42852 24368 42874 24672
rect 42908 24368 42930 24672
rect 42958 23820 42992 25188
rect 43510 25164 43555 26300
rect 43644 26299 43656 26300
rect 43605 26288 43661 26299
rect 43616 25164 43661 26288
rect 43672 26284 43684 26328
rect 44256 26304 44308 26332
rect 44256 26300 44262 26304
rect 44268 26288 44302 26304
rect 43510 23820 43544 25164
rect 43616 24602 43650 25164
rect 43582 23820 43594 24602
rect 43610 23820 43656 24602
rect 43672 24307 43684 24602
rect 44268 24307 44308 26288
rect 44314 24307 44319 26299
rect 44575 25133 53013 26338
rect 44932 24604 44966 25133
rect 44898 24307 44924 24604
rect 44926 24307 44972 24604
rect 44986 24307 45000 24604
rect 45046 24307 45080 25133
rect 50216 24307 50226 24502
rect 50244 24307 50254 24474
rect 43672 23820 52121 24307
rect 41528 23786 52121 23820
rect 41528 23538 41562 23786
rect 41642 23678 41676 23786
rect 41994 23756 42028 23786
rect 42300 23756 42334 23786
rect 41994 23718 42032 23756
rect 42272 23718 42334 23756
rect 42752 23756 42786 23786
rect 42958 23756 42992 23786
rect 42752 23718 42790 23756
rect 42930 23718 42992 23756
rect 43510 23756 43544 23786
rect 43610 23756 43656 23786
rect 43510 23718 43548 23756
rect 43588 23724 43656 23756
rect 43672 23724 52121 23786
rect 43582 23718 43656 23724
rect 43666 23718 52121 23724
rect 41688 23684 42334 23718
rect 42346 23684 42992 23718
rect 43004 23684 43656 23718
rect 43662 23684 52121 23718
rect 54880 23690 54914 27248
rect 56445 25046 58096 27248
rect 56445 25026 58174 25046
rect 56445 25018 58096 25026
rect 56445 24998 58146 25018
rect 56445 24943 58096 24998
rect 56445 24909 60480 24943
rect 56445 24759 58096 24909
rect 56756 24758 57304 24759
rect 57354 24704 57992 24759
rect 57286 24592 57290 24594
rect 57928 24374 57946 24532
rect 57966 24408 57984 24494
rect 58026 24374 58060 24759
rect 57928 24370 58146 24374
rect 57946 24356 58146 24370
rect 58026 24340 58060 24356
rect 57946 24322 58180 24340
rect 58026 24320 58060 24322
rect 56614 24286 60480 24320
rect 42300 23678 42334 23684
rect 42958 23678 42992 23684
rect 43582 23678 43600 23684
rect 43610 23678 43656 23684
rect 43666 23678 52121 23684
rect 41630 23640 41688 23678
rect 41966 23640 42004 23678
rect 42288 23640 42346 23678
rect 42724 23640 42762 23678
rect 42946 23640 43004 23678
rect 43482 23640 43520 23678
rect 43604 23646 43662 23678
rect 43672 23646 52121 23678
rect 41630 23606 42004 23640
rect 42056 23606 42762 23640
rect 42814 23606 43520 23640
rect 43560 23640 43662 23646
rect 43683 23640 52121 23646
rect 43560 23606 52121 23640
rect 53302 23622 53348 23646
rect 41630 23590 41688 23606
rect 42288 23590 42346 23606
rect 42946 23590 43004 23606
rect 43560 23600 43588 23606
rect 43604 23590 43662 23606
rect 41630 23575 41676 23590
rect 41642 23538 41676 23575
rect 42300 23538 42334 23590
rect 42958 23538 42992 23590
rect 43616 23538 43650 23590
rect 43683 23538 52121 23606
rect 53310 23600 53348 23622
rect 53366 23572 53376 23674
rect 56614 23640 56648 24286
rect 57154 24206 57188 24286
rect 57316 24206 57900 24217
rect 57912 24206 57946 24286
rect 58026 24206 58060 24286
rect 64788 24212 64804 24318
rect 56678 24144 56750 24182
rect 56800 24172 58094 24206
rect 57141 24160 57142 24161
rect 57142 24159 57143 24160
rect 56716 23640 56750 24144
rect 57154 23690 57188 24172
rect 57200 24160 57201 24161
rect 57899 24160 57900 24161
rect 57912 24160 57946 24172
rect 57199 24159 57200 24160
rect 57900 24159 57901 24160
rect 57912 23896 57957 24160
rect 58026 23896 58060 24172
rect 64778 24166 64804 24212
rect 64788 24088 64804 24166
rect 64806 24138 64816 24240
rect 64806 24094 64820 24116
rect 64778 24066 64820 24088
rect 56787 23678 56788 23679
rect 56788 23677 56789 23678
rect 57126 23640 57164 23678
rect 57462 23640 60428 23896
rect 56614 23606 57164 23640
rect 57216 23614 60428 23640
rect 56614 23538 56648 23606
rect 56716 23576 56750 23606
rect 57026 23600 57138 23606
rect 57204 23600 60428 23614
rect 57462 23586 60428 23600
rect 57054 23572 57166 23586
rect 57176 23572 60428 23586
rect 56716 23560 56750 23572
rect 56800 23538 60428 23572
rect 31219 23504 31321 23538
rect 31994 23504 60428 23538
rect 31219 23468 31303 23504
rect 31994 23468 41502 23504
rect 31105 22304 31139 22316
rect 27851 22218 27855 22291
rect 27879 22257 27883 22263
rect 28459 22257 31139 22304
rect 27875 22223 27883 22257
rect 27891 22223 28507 22257
rect 28533 22223 28541 22257
rect 28549 22223 29165 22257
rect 27879 22218 27883 22223
rect 28461 22218 28507 22223
rect 29119 22218 29165 22223
rect 29167 22218 29171 22257
rect 29195 22218 29199 22257
rect 29207 22223 29823 22257
rect 29865 22223 30481 22257
rect 27665 22155 29378 22218
rect 29712 22210 29714 22217
rect 29740 22182 29742 22217
rect 29777 22207 29823 22223
rect 30435 22207 30481 22223
rect 29789 22155 29823 22207
rect 30447 22155 30481 22207
rect 30483 22189 30487 22257
rect 30511 22217 30515 22257
rect 30523 22223 31139 22257
rect 31034 22210 31036 22217
rect 31062 22182 31064 22217
rect 31093 22207 31139 22223
rect 31105 22155 31139 22207
rect 31219 22217 31267 23468
rect 32030 22944 32064 23468
rect 32026 22910 32320 22944
rect 32030 22783 32064 22910
rect 32144 22889 32178 22910
rect 32010 22749 32064 22783
rect 32032 22573 32098 22749
rect 32110 22614 32120 22800
rect 32132 22761 32178 22889
rect 32138 22749 32178 22761
rect 32190 22749 32217 22760
rect 32138 22586 32217 22749
rect 32144 22573 32217 22586
rect 32030 22412 32064 22573
rect 32144 22561 32178 22573
rect 32132 22449 32178 22561
rect 32144 22412 32178 22449
rect 32286 22412 32320 22910
rect 32026 22378 32320 22412
rect 32736 22890 36374 23468
rect 36457 22890 36491 23468
rect 36571 23454 36616 23468
rect 36571 22942 36605 23454
rect 36758 23452 37148 23468
rect 36758 22954 36792 23452
rect 36972 23384 37019 23431
rect 36934 23350 37019 23384
rect 36861 23291 36906 23302
rect 36989 23291 37034 23302
rect 36872 23115 36906 23291
rect 37000 23115 37034 23291
rect 36972 23056 37019 23103
rect 36934 23022 37019 23056
rect 37114 22954 37148 23452
rect 36571 22918 36616 22942
rect 36758 22920 37148 22954
rect 37229 23452 37624 23468
rect 37229 23390 37274 23452
rect 37229 23016 37268 23390
rect 37440 23384 37495 23431
rect 37410 23350 37495 23384
rect 37337 23291 37382 23302
rect 37465 23291 37521 23302
rect 37348 23115 37382 23291
rect 37476 23115 37521 23291
rect 37440 23056 37495 23103
rect 37410 23022 37495 23056
rect 37229 22954 37274 23016
rect 37590 22954 37624 23452
rect 37229 22920 37624 22954
rect 37772 23332 38613 23468
rect 36512 22890 36616 22918
rect 36988 22890 37060 22918
rect 32736 22870 37082 22890
rect 37229 22870 37274 22920
rect 32736 22832 37162 22870
rect 37216 22832 37638 22870
rect 32030 22328 32064 22378
rect 27665 22121 31151 22155
rect 27520 10504 27584 20616
rect 27665 18286 29378 22121
rect 29789 18286 29823 20160
rect 30447 18286 30481 20160
rect 31105 18286 31139 20160
rect 27665 18239 31139 18286
rect 27665 18205 29829 18239
rect 27665 18137 29378 18205
rect 29755 18199 29773 18205
rect 29783 18171 29829 18205
rect 29839 18205 30487 18239
rect 29839 18199 29857 18205
rect 30413 18199 30431 18205
rect 30441 18171 30487 18205
rect 30497 18205 31139 18239
rect 30497 18199 30515 18205
rect 31071 18199 31089 18205
rect 31099 18171 31139 18205
rect 29789 18137 29823 18171
rect 30447 18137 30481 18171
rect 31105 18137 31139 18171
rect 27665 18103 31173 18137
rect 27665 15768 29378 18103
rect 31219 15545 31253 22217
rect 31994 22044 32338 22328
rect 32736 22250 37638 22832
rect 32736 22044 37534 22250
rect 37772 22044 38590 23332
rect 39203 22044 39248 23468
rect 39861 22942 39895 23468
rect 39861 22880 39906 22942
rect 39975 22880 40009 23468
rect 41318 23036 41352 23468
rect 41318 22954 41408 23036
rect 40686 22910 41076 22944
rect 39420 22330 40244 22880
rect 40686 22412 40720 22910
rect 40815 22842 40947 22889
rect 40862 22808 40947 22842
rect 40789 22749 40845 22760
rect 40917 22749 40973 22760
rect 40800 22573 40845 22749
rect 40928 22573 40973 22749
rect 40815 22514 40947 22561
rect 40862 22480 40947 22514
rect 41042 22412 41076 22910
rect 40686 22378 41076 22412
rect 39454 22044 39666 22330
rect 39846 22310 39916 22330
rect 39861 22044 39906 22310
rect 39975 22044 40009 22330
rect 40110 22244 40228 22330
rect 40672 22044 41094 22328
rect 41318 22044 41352 22954
rect 31994 22010 41364 22044
rect 31994 21989 32338 22010
rect 32736 21989 37534 22010
rect 37772 21989 38590 22010
rect 39203 21989 39248 22010
rect 31994 21942 39486 21989
rect 39861 21942 39895 22010
rect 39975 21942 40009 22010
rect 40672 21942 41094 22010
rect 41318 21989 41352 22010
rect 41290 21942 41352 21989
rect 31994 21908 41352 21942
rect 31994 21708 32338 21908
rect 32030 21192 32064 21708
rect 32030 20924 32302 21192
rect 32002 20802 32302 20924
rect 32030 20748 32302 20802
rect 32030 20290 32064 20748
rect 32026 20256 32320 20290
rect 32030 20160 32064 20256
rect 32036 20129 32064 20160
rect 32010 20095 32064 20129
rect 32132 20219 32144 20235
rect 32132 20204 32147 20219
rect 32132 20160 32160 20204
rect 32132 20107 32178 20160
rect 32144 20095 32178 20107
rect 32190 20095 32217 20106
rect 32032 19919 32098 20095
rect 32144 19919 32217 20095
rect 32030 19758 32064 19919
rect 32144 19907 32178 19919
rect 32132 19795 32178 19907
rect 32144 19758 32178 19795
rect 32286 19758 32320 20256
rect 32026 19724 32320 19758
rect 32030 19674 32064 19724
rect 31994 19605 32338 19674
rect 32736 19605 37534 21908
rect 37772 21902 38590 21908
rect 37772 19605 38613 21902
rect 39203 19605 39248 21908
rect 31994 19558 39486 19605
rect 39861 19558 39895 21908
rect 39975 19558 40009 21908
rect 40672 21708 41094 21908
rect 41318 20382 41352 21908
rect 41318 20300 41400 20382
rect 40686 20256 41076 20290
rect 40686 19758 40720 20256
rect 40900 20188 40947 20235
rect 40862 20154 40947 20188
rect 40789 20095 40834 20106
rect 40917 20095 40962 20106
rect 40800 19919 40834 20095
rect 40928 19919 40962 20095
rect 40900 19860 40947 19907
rect 40862 19826 40947 19860
rect 41042 19758 41076 20256
rect 40686 19724 41076 19758
rect 40672 19558 41094 19674
rect 41318 19605 41352 20300
rect 41290 19558 41352 19605
rect 31994 19524 41352 19558
rect 31994 19456 32338 19524
rect 32736 19468 37534 19524
rect 37772 19518 38590 19524
rect 32736 19456 37610 19468
rect 37772 19456 38613 19518
rect 39203 19456 39248 19524
rect 39861 19456 39895 19524
rect 39975 19456 40009 19524
rect 40672 19456 41094 19524
rect 41318 19456 41352 19524
rect 31994 19422 41364 19456
rect 41370 19422 41386 19456
rect 31994 19054 32338 19422
rect 32736 18936 37534 19422
rect 37576 18936 37610 19422
rect 32736 18902 37610 18936
rect 32030 18802 32064 18856
rect 32736 18852 37534 18902
rect 32128 18802 32178 18836
rect 32736 18802 37624 18852
rect 37772 18802 38613 19422
rect 39203 18802 39248 19422
rect 39861 18802 39895 19422
rect 39975 18802 40009 19422
rect 40672 19054 41094 19422
rect 41318 18802 41352 19422
rect 32066 18768 32118 18802
rect 32132 18768 41364 18802
rect 32032 18706 32064 18740
rect 32066 10842 32100 18768
rect 32132 18645 32154 18768
rect 32736 18747 37624 18768
rect 37772 18747 38613 18768
rect 39203 18747 39248 18768
rect 32195 18700 39486 18747
rect 39861 18700 39895 18768
rect 39975 18700 40009 18768
rect 41318 18747 41352 18768
rect 41318 18716 41364 18747
rect 41306 18700 41364 18716
rect 32242 18666 41364 18700
rect 32132 15873 32178 18645
rect 32190 18607 32225 18618
rect 32132 15861 32154 15873
rect 32180 15861 32225 18607
rect 32736 18286 37624 18666
rect 37772 18660 38590 18666
rect 37772 18286 38613 18660
rect 39203 18286 39248 18666
rect 39861 18286 39895 18666
rect 32736 18239 39486 18286
rect 39833 18239 39895 18286
rect 32736 18205 39248 18239
rect 39265 18205 39895 18239
rect 32736 18137 37534 18205
rect 37772 18137 38613 18205
rect 39203 18137 39248 18205
rect 39861 18137 39895 18205
rect 39975 18137 40009 18666
rect 41306 18657 41342 18666
rect 41306 18619 41352 18657
rect 32736 18103 40009 18137
rect 32736 17440 37534 18103
rect 37772 17758 38613 18103
rect 32736 16200 36360 17440
rect 36457 16200 36491 17440
rect 36571 17004 36605 17440
rect 37229 17004 37263 17440
rect 36571 16782 36616 17004
rect 37229 16814 37274 17004
rect 36571 16200 36605 16782
rect 36744 16780 37134 16814
rect 36744 16282 36778 16780
rect 36958 16712 37005 16759
rect 36920 16678 37005 16712
rect 36847 16619 36892 16630
rect 36975 16619 37020 16630
rect 36858 16443 36892 16619
rect 36986 16443 37020 16619
rect 36958 16384 37005 16431
rect 36920 16350 37005 16384
rect 37100 16282 37134 16780
rect 37220 16780 37610 16814
rect 37220 16752 37263 16780
rect 37220 16355 37288 16752
rect 37434 16712 37481 16759
rect 37396 16678 37481 16712
rect 37323 16619 37368 16630
rect 37451 16619 37507 16630
rect 37334 16443 37368 16619
rect 37462 16443 37507 16619
rect 37434 16384 37481 16431
rect 37218 16344 37288 16355
rect 37396 16350 37481 16384
rect 36744 16248 37134 16282
rect 37220 16282 37263 16344
rect 37576 16282 37610 16780
rect 37220 16248 37610 16282
rect 37772 16570 38590 17758
rect 37229 16200 37263 16248
rect 32736 16198 37544 16200
rect 32736 16166 37624 16198
rect 32736 16086 36360 16166
rect 36457 16156 36514 16166
rect 36457 16138 36491 16156
rect 36508 16138 36514 16156
rect 36412 16100 36491 16138
rect 36452 16086 36491 16100
rect 36571 16086 36605 16166
rect 36726 16086 37148 16166
rect 37202 16086 37624 16166
rect 32736 16052 37624 16086
rect 32736 15861 36360 16052
rect 36452 16048 36491 16052
rect 36452 15986 36454 16048
rect 32168 15814 36360 15861
rect 36457 15814 36491 16048
rect 36508 15986 36510 16048
rect 36571 15861 36605 16052
rect 36571 15814 36618 15861
rect 36726 15814 37148 16052
rect 37202 15814 37624 16052
rect 37772 15861 38613 16570
rect 39203 15861 39248 18103
rect 39861 15861 39895 18103
rect 37654 15814 39486 15861
rect 39861 15814 39908 15861
rect 39975 15814 40009 18103
rect 40584 18154 40974 18188
rect 40584 17656 40618 18154
rect 40798 18086 40845 18133
rect 40760 18052 40845 18086
rect 40687 17993 40732 18004
rect 40815 17993 40860 18004
rect 40698 17817 40732 17993
rect 40826 17817 40860 17993
rect 40798 17758 40845 17805
rect 40760 17724 40845 17758
rect 40940 17656 40974 18154
rect 40584 17622 40974 17656
rect 40566 16952 40988 17572
rect 41318 17564 41352 18619
rect 41354 18607 41386 18623
rect 41354 17564 41388 18607
rect 41432 17624 41466 23468
rect 41492 22942 41502 23468
rect 41492 22010 41522 22942
rect 41492 18838 41502 22010
rect 41528 18838 41562 23504
rect 41492 18768 41562 18838
rect 41468 17624 41562 18768
rect 41642 18296 41676 23504
rect 41680 22344 41682 22400
rect 41680 22088 41682 22144
rect 41680 21944 41682 22000
rect 41680 21688 41682 21744
rect 41680 19690 41714 19746
rect 41708 19490 41714 19690
rect 41736 19490 41742 19690
rect 41680 19434 41714 19490
rect 41680 19290 41714 19346
rect 41708 19090 41714 19290
rect 41736 19090 41742 19290
rect 41680 19034 41714 19090
rect 42300 18300 42334 23504
rect 42958 18300 42992 23504
rect 43576 21948 43588 23052
rect 43616 18300 43650 23504
rect 43683 23468 52121 23504
rect 43683 21508 45116 23468
rect 56614 22188 56648 23504
rect 56716 23470 56750 23502
rect 57462 22958 60428 23504
rect 60974 22462 62624 23900
rect 63060 22460 64710 23898
rect 64788 23762 64804 24066
rect 64826 23576 64860 24144
rect 64866 24094 64920 24116
rect 64866 24066 64892 24088
rect 64788 23456 64804 23460
rect 56440 22182 58748 22188
rect 54490 22152 58748 22182
rect 54540 22000 54554 22102
rect 54568 22028 54610 22074
rect 56214 22034 56436 22054
rect 56252 21996 56398 22016
rect 43683 21491 50408 21508
rect 43683 21474 45116 21491
rect 43683 21440 50470 21474
rect 43683 21360 45116 21440
rect 45594 21360 50286 21371
rect 43683 21326 50286 21360
rect 43683 20867 45116 21326
rect 50287 21298 50415 21345
rect 46884 21040 47330 21146
rect 46748 20964 47330 21040
rect 46884 20904 47330 20964
rect 45690 20878 48010 20890
rect 50334 20880 50415 21298
rect 50287 20878 50415 20880
rect 45594 20867 50415 20878
rect 50436 20867 50470 21440
rect 56440 21242 58748 22152
rect 59018 21246 61326 22194
rect 61488 21666 61744 21668
rect 61516 21638 61716 21640
rect 64788 21580 64804 21684
rect 64778 21534 64804 21580
rect 59018 21242 62624 21246
rect 43683 20833 50504 20867
rect 43683 20753 45116 20833
rect 45690 20753 45724 20833
rect 47834 20788 47881 20833
rect 45866 20787 47881 20788
rect 45850 20754 47881 20787
rect 46028 20753 46084 20754
rect 47578 20753 47634 20754
rect 47976 20753 48010 20833
rect 50287 20826 50415 20833
rect 50287 20821 50399 20826
rect 50216 20753 50328 20758
rect 50374 20753 50376 20758
rect 50436 20753 50470 20833
rect 56440 20756 62624 21242
rect 43683 20719 51989 20753
rect 56440 20750 60440 20756
rect 43683 20708 45116 20719
rect 45690 20718 45724 20719
rect 45218 20714 45852 20718
rect 45218 20708 47850 20714
rect 47862 20708 47896 20711
rect 47976 20708 48010 20719
rect 50244 20708 50328 20719
rect 43683 20707 50328 20708
rect 43683 20702 46084 20707
rect 47578 20702 50328 20707
rect 43683 20696 50328 20702
rect 50374 20696 50432 20719
rect 43683 20685 50291 20696
rect 43683 20683 45116 20685
rect 44068 19272 45116 20683
rect 45690 20668 48050 20685
rect 45690 20044 45724 20668
rect 45804 20044 45838 20668
rect 47794 20662 47856 20668
rect 45850 20656 45851 20657
rect 45849 20655 45850 20656
rect 47822 20634 47856 20660
rect 47862 20618 47896 20668
rect 47902 20662 48050 20668
rect 47976 20660 48010 20662
rect 47902 20634 48022 20660
rect 47976 20618 48010 20634
rect 47860 20570 48010 20618
rect 47850 20500 48010 20570
rect 46894 20246 47340 20488
rect 47850 20268 47910 20500
rect 47014 20160 47254 20246
rect 46028 20092 46084 20106
rect 47724 20092 47780 20106
rect 45849 20056 45850 20057
rect 47850 20056 47851 20057
rect 47862 20056 47896 20268
rect 45850 20055 45851 20056
rect 46028 20044 46084 20050
rect 47324 20044 47944 20056
rect 47976 20044 48010 20500
rect 50436 20160 50470 20719
rect 56708 20566 56742 20750
rect 57462 20732 60428 20750
rect 60974 20732 62624 20756
rect 63060 20732 64710 21244
rect 64788 21108 64804 21534
rect 64806 21506 64816 21608
rect 64826 21602 64860 22170
rect 64826 20944 64860 21512
rect 65108 21108 65118 21332
rect 65108 20802 65118 20806
rect 58448 20704 58744 20732
rect 59792 20704 60088 20732
rect 61010 20618 61044 20732
rect 61366 20730 61618 20732
rect 61400 20696 61622 20700
rect 61112 20618 61142 20636
rect 56500 20532 57324 20566
rect 45690 20042 48010 20044
rect 45690 20010 48560 20042
rect 45690 19468 45724 20010
rect 45804 19658 45838 20010
rect 45850 19998 45851 19999
rect 45849 19997 45850 19998
rect 47324 19794 47944 20010
rect 46894 19776 47944 19794
rect 46638 19662 47944 19776
rect 45804 19468 45849 19658
rect 46894 19634 47944 19662
rect 47976 20008 48560 20010
rect 47976 19686 48028 20008
rect 48526 19994 48560 20008
rect 48366 19984 49406 19994
rect 48365 19928 48376 19939
rect 48049 19866 48130 19913
rect 48189 19894 48376 19928
rect 48377 19866 48458 19913
rect 48096 19828 48130 19866
rect 48424 19828 48458 19866
rect 48365 19800 48376 19811
rect 48189 19766 48376 19800
rect 48526 19686 48560 19984
rect 47976 19652 48560 19686
rect 49250 19718 50506 19754
rect 54394 19718 54428 20160
rect 49250 19684 54606 19718
rect 46894 19552 47340 19634
rect 45500 19434 45890 19468
rect 45500 19386 45534 19434
rect 45690 19400 45724 19434
rect 45642 19399 45724 19400
rect 45629 19386 45724 19399
rect 45804 19386 45838 19434
rect 45849 19398 45850 19399
rect 45850 19397 45851 19398
rect 45856 19386 45890 19434
rect 45976 19434 46366 19468
rect 45976 19386 46010 19434
rect 46118 19399 46224 19400
rect 46105 19386 46237 19399
rect 46332 19386 46366 19434
rect 47850 19398 47851 19399
rect 47849 19397 47850 19398
rect 47182 19386 47400 19397
rect 47730 19386 47780 19392
rect 47862 19386 47896 19634
rect 47976 19386 48010 19652
rect 49250 19386 50506 19684
rect 45500 19352 50506 19386
rect 45500 19280 45534 19352
rect 45645 19340 45748 19352
rect 45690 19332 45748 19340
rect 45804 19339 45838 19352
rect 45302 19272 45592 19280
rect 45614 19272 45648 19306
rect 45690 19272 45724 19332
rect 45792 19313 45842 19339
rect 45778 19312 45842 19313
rect 45770 19306 45778 19312
rect 45742 19285 45778 19306
rect 45742 19280 45782 19285
rect 45792 19280 45842 19312
rect 45856 19280 45890 19352
rect 45976 19280 46010 19352
rect 46028 19312 46084 19336
rect 46152 19332 46237 19352
rect 46090 19284 46124 19306
rect 46218 19284 46252 19306
rect 46079 19280 46124 19284
rect 45742 19272 45776 19280
rect 45778 19272 45842 19280
rect 45844 19273 46124 19280
rect 46207 19273 46252 19284
rect 45844 19272 46084 19273
rect 46090 19272 46124 19273
rect 46218 19272 46252 19273
rect 46332 19272 46366 19352
rect 47182 19286 47400 19306
rect 47862 19272 47896 19352
rect 47976 19272 48010 19352
rect 49250 19272 50506 19352
rect 44068 19238 50506 19272
rect 44068 19236 45116 19238
rect 45500 19236 45534 19238
rect 45690 19236 45724 19238
rect 45742 19236 45758 19238
rect 45766 19236 45776 19238
rect 45792 19236 45842 19238
rect 45856 19236 45890 19238
rect 45976 19236 46010 19238
rect 46090 19236 46124 19238
rect 46218 19236 46252 19238
rect 46332 19236 46366 19238
rect 47976 19236 48010 19238
rect 49250 19236 50506 19238
rect 44068 19202 50506 19236
rect 44274 19200 44308 19202
rect 44932 19200 44966 19202
rect 45046 19200 45080 19202
rect 45464 19200 48046 19202
rect 49286 19200 49320 19202
rect 49400 19200 49434 19202
rect 43742 19166 52090 19200
rect 43742 18300 43776 19166
rect 44184 19092 44196 19150
rect 44212 19092 44224 19122
rect 44274 19086 44308 19166
rect 44932 19086 44966 19166
rect 45046 19086 45080 19166
rect 43806 19024 43878 19062
rect 43928 19052 45080 19086
rect 43844 18456 43878 19024
rect 44184 18986 44196 19046
rect 44212 19014 44224 19046
rect 44261 19040 44262 19041
rect 44262 19039 44263 19040
rect 44274 18880 44308 19052
rect 44320 19040 44321 19041
rect 44919 19040 44920 19041
rect 44319 19039 44320 19040
rect 44920 19039 44921 19040
rect 44932 18880 44966 19052
rect 45046 18880 45080 19052
rect 45464 18880 48046 19166
rect 49286 19086 49320 19166
rect 49400 19086 49434 19166
rect 49446 19086 51915 19097
rect 49286 19052 51915 19086
rect 49286 18880 49320 19052
rect 49400 19040 49434 19052
rect 49446 19040 49447 19041
rect 49400 19039 49446 19040
rect 49400 18880 49445 19039
rect 51916 19024 52026 19062
rect 44068 18744 50506 18880
rect 51916 18744 51917 18745
rect 51954 18744 52026 19024
rect 44068 18706 51916 18744
rect 51954 18706 51988 18744
rect 52056 18706 52090 19166
rect 44068 18672 52090 18706
rect 44068 18604 50506 18672
rect 51954 18604 51988 18672
rect 52056 18604 52090 18672
rect 54394 18604 54428 19684
rect 54430 19582 54462 19616
rect 54480 19544 54488 19674
rect 54496 19544 54530 19570
rect 54465 19532 54530 19544
rect 54458 19038 54530 19532
rect 54458 19007 54504 19038
rect 54458 19000 54492 19007
rect 54458 18986 54462 19000
rect 54458 18948 54504 18986
rect 54458 18756 54530 18948
rect 54540 18942 54554 19044
rect 54572 19016 54606 19684
rect 56500 19534 56534 20532
rect 56618 20480 56656 20522
rect 56580 20392 56606 20414
rect 56626 20396 56646 20480
rect 56660 20470 56698 20480
rect 56660 20448 56702 20470
rect 56708 20448 56742 20532
rect 56660 20424 56742 20448
rect 56638 20392 56640 20396
rect 56660 20392 56698 20424
rect 56580 20380 56678 20392
rect 56602 19534 56674 20380
rect 56708 19534 56742 20424
rect 57654 20304 58646 20602
rect 58964 20304 59956 20610
rect 60132 20304 60428 20618
rect 60974 20352 61142 20618
rect 61292 20540 62624 20622
rect 63060 20540 64710 20622
rect 61236 20518 62750 20540
rect 62942 20518 64718 20540
rect 61236 20516 62770 20518
rect 62780 20516 64744 20518
rect 61236 20508 62750 20516
rect 62942 20508 64718 20516
rect 60830 20350 61142 20352
rect 61292 20490 62624 20508
rect 63060 20490 64710 20508
rect 61292 20488 62742 20490
rect 62808 20488 64716 20490
rect 61292 20484 62624 20488
rect 63060 20484 64710 20488
rect 61292 20480 62750 20484
rect 62942 20480 64746 20484
rect 60830 20316 61158 20350
rect 61292 20316 62624 20480
rect 60178 20298 60202 20304
rect 60294 20298 60316 20304
rect 60232 20264 60256 20298
rect 60270 20264 60780 20298
rect 60198 20202 60202 20236
rect 57758 20132 57844 20160
rect 57672 20116 57844 20132
rect 57672 19978 57826 20116
rect 60232 19982 60266 20264
rect 60270 20178 60320 20264
rect 60407 20184 60605 20195
rect 60270 20140 60406 20178
rect 60418 20150 60605 20184
rect 60606 20140 60716 20178
rect 60270 20090 60328 20140
rect 60334 20106 60406 20140
rect 60407 20096 60605 20107
rect 60644 20106 60716 20140
rect 60270 19982 60320 20090
rect 60418 20062 60605 20096
rect 60746 19982 60780 20264
rect 60232 19948 60256 19982
rect 60270 19948 60780 19982
rect 60830 20282 62624 20316
rect 60830 20202 61158 20282
rect 61237 20202 61248 20213
rect 60830 20168 61248 20202
rect 61292 20187 62624 20282
rect 60830 20074 61158 20168
rect 61170 20156 61171 20157
rect 61169 20155 61170 20156
rect 61249 20140 62624 20187
rect 61169 20086 61170 20087
rect 61170 20085 61171 20086
rect 61237 20074 61248 20085
rect 60830 20040 61248 20074
rect 60830 20039 61158 20040
rect 60830 20028 61124 20039
rect 60830 20027 61142 20028
rect 60830 19932 61124 20027
rect 61292 19994 62624 20140
rect 61186 19980 62624 19994
rect 61292 19960 62624 19980
rect 61159 19949 62624 19960
rect 61170 19932 62624 19949
rect 60830 19926 62624 19932
rect 60830 19890 61124 19926
rect 60974 19808 61124 19890
rect 61292 19808 62624 19926
rect 59000 19540 59034 19558
rect 56440 19249 57456 19534
rect 57654 19249 58646 19534
rect 59000 19504 59956 19540
rect 58678 19249 58712 19402
rect 59018 19285 59956 19504
rect 58964 19249 59956 19285
rect 60132 19316 61124 19540
rect 61136 19316 61140 19321
rect 60132 19249 61140 19316
rect 61142 19249 61176 19283
rect 61256 19249 61290 19408
rect 61292 19285 61326 19540
rect 61328 19285 61344 19558
rect 61442 19285 61476 19808
rect 63060 19806 64710 20480
rect 63424 19792 64220 19806
rect 65200 19539 65234 23768
rect 66008 23676 66012 23681
rect 66008 23490 66036 23676
rect 66008 21210 66012 23490
rect 67940 21210 67944 23681
rect 68464 22352 68712 22372
rect 68484 22161 68485 22352
rect 68692 22161 68712 22352
rect 68484 22160 68712 22161
rect 65302 21176 68650 21210
rect 65314 21142 65348 21176
rect 65972 21170 66006 21176
rect 66008 21170 66012 21176
rect 65966 21155 66012 21170
rect 66630 21155 66664 21176
rect 67288 21155 67322 21176
rect 67940 21170 67944 21176
rect 67946 21170 67980 21176
rect 67940 21155 67986 21170
rect 68604 21155 68638 21176
rect 65314 21040 65354 21142
rect 65944 21114 66012 21155
rect 65364 21108 65382 21114
rect 65938 21108 66012 21114
rect 66022 21108 66040 21114
rect 66602 21108 66664 21155
rect 67260 21108 67322 21155
rect 67918 21114 67986 21155
rect 68576 21114 68638 21155
rect 67912 21108 67986 21114
rect 67996 21108 68014 21114
rect 68570 21108 68638 21114
rect 65360 21074 66012 21108
rect 66018 21074 66664 21108
rect 66676 21074 67322 21108
rect 67334 21074 67986 21108
rect 67992 21074 68638 21108
rect 65364 21068 65382 21074
rect 65938 21068 65956 21074
rect 65314 19668 65348 21040
rect 65966 21022 66012 21074
rect 66022 21068 66040 21074
rect 65972 21012 66036 21022
rect 65972 19696 66006 21012
rect 66008 20836 66036 21012
rect 66008 20654 66012 20836
rect 66008 19696 66012 20516
rect 65966 19681 66012 19696
rect 66630 19681 66664 21074
rect 67288 19681 67322 21074
rect 67912 21068 67930 21074
rect 67940 21012 67986 21074
rect 67996 21068 68014 21074
rect 68570 21068 68588 21074
rect 68598 21040 68638 21074
rect 67940 19894 67944 21012
rect 65314 19566 65354 19668
rect 65944 19640 66012 19681
rect 65364 19634 65382 19640
rect 65938 19634 66012 19640
rect 66022 19634 66040 19640
rect 66602 19634 66664 19681
rect 67260 19634 67322 19681
rect 67754 19634 67830 19804
rect 67834 19634 67890 19864
rect 67918 19696 67944 19894
rect 67946 19696 67980 21012
rect 68604 19718 68638 21040
rect 68464 19698 68712 19718
rect 67918 19686 67980 19696
rect 67940 19681 67986 19686
rect 67918 19640 67986 19681
rect 67912 19634 67986 19640
rect 67996 19634 68014 19640
rect 68484 19634 68485 19698
rect 68604 19681 68638 19698
rect 68576 19640 68638 19681
rect 68570 19634 68638 19640
rect 65360 19600 66012 19634
rect 66018 19600 66664 19634
rect 66676 19600 67322 19634
rect 67334 19600 67986 19634
rect 67992 19600 68638 19634
rect 65364 19594 65382 19600
rect 65938 19594 65956 19600
rect 61292 19249 64916 19285
rect 56440 19215 64916 19249
rect 56440 19182 57456 19215
rect 57654 19182 58646 19215
rect 56440 19146 56778 19182
rect 56440 19135 57236 19146
rect 57248 19135 57282 19182
rect 57294 19135 57894 19146
rect 57906 19135 57940 19182
rect 57952 19135 58552 19146
rect 58564 19135 58598 19182
rect 58678 19135 58712 19215
rect 54568 18970 54610 19016
rect 56122 18976 56248 19048
rect 54465 18744 54530 18756
rect 54430 18672 54462 18706
rect 54480 18656 54488 18744
rect 54496 18718 54530 18744
rect 54572 18604 54606 18970
rect 56066 18944 56248 18976
rect 56440 19022 56778 19135
rect 56786 19101 58712 19135
rect 56844 19022 57096 19101
rect 57235 19089 57236 19090
rect 57248 19089 57282 19101
rect 57862 19095 57900 19101
rect 57294 19089 57295 19090
rect 57893 19089 57894 19090
rect 57906 19089 57940 19101
rect 57946 19095 58004 19101
rect 57952 19089 57953 19090
rect 58551 19089 58552 19090
rect 58564 19089 58598 19101
rect 57236 19088 57237 19089
rect 57248 19088 57294 19089
rect 57894 19088 57895 19089
rect 57906 19088 57952 19089
rect 58552 19088 58553 19089
rect 57248 19046 57293 19088
rect 57906 19082 57951 19088
rect 57890 19067 57900 19082
rect 57906 19067 58004 19082
rect 57218 19026 57242 19046
rect 57248 19026 57312 19046
rect 56066 18806 56234 18944
rect 56246 18792 56250 18814
rect 56246 18736 56306 18758
rect 56440 18750 57128 19022
rect 57248 19018 57293 19026
rect 57190 18998 57242 19018
rect 57248 18998 57340 19018
rect 44068 18570 54606 18604
rect 44068 18472 50506 18570
rect 44068 18450 51340 18472
rect 44068 18428 50506 18450
rect 43806 18366 43878 18404
rect 43928 18394 50506 18428
rect 41642 18194 41682 18296
rect 41692 18262 41710 18268
rect 42272 18262 42334 18300
rect 42680 18262 43780 18300
rect 43844 18262 43878 18366
rect 44068 18262 50506 18394
rect 41688 18228 42334 18262
rect 42346 18228 43656 18262
rect 41692 18222 41710 18228
rect 41642 18160 41676 18194
rect 42300 18160 42334 18228
rect 42932 18190 42992 18228
rect 43582 18222 43600 18228
rect 43610 18194 43656 18228
rect 43666 18260 50506 18262
rect 52056 18260 52090 18570
rect 54394 18260 54428 18570
rect 56440 18488 56778 18750
rect 57248 18490 57293 18998
rect 57906 18590 57951 19067
rect 57954 18946 58336 19018
rect 57954 18840 58422 18946
rect 57954 18780 58336 18840
rect 57884 18496 57964 18590
rect 57236 18489 57237 18490
rect 57248 18489 57294 18490
rect 57235 18488 57236 18489
rect 56440 18477 57236 18488
rect 57248 18477 57282 18489
rect 57294 18488 57295 18489
rect 57482 18488 58136 18496
rect 58552 18489 58553 18490
rect 58564 18489 58609 19089
rect 58551 18488 58552 18489
rect 57294 18477 58552 18488
rect 58564 18477 58598 18489
rect 58678 18477 58712 19101
rect 58964 19146 59956 19215
rect 60132 19146 61140 19215
rect 58964 19141 61140 19146
rect 58964 19135 61124 19141
rect 61142 19135 61176 19215
rect 61256 19135 61290 19215
rect 61292 19135 64916 19215
rect 58964 19124 64916 19135
rect 58964 19101 61290 19124
rect 58758 18946 58764 19098
rect 58786 18968 58820 19098
rect 58964 18682 59956 19101
rect 60132 18682 61124 19101
rect 61129 19089 61130 19090
rect 61130 19088 61131 19089
rect 61136 19018 61140 19095
rect 58964 18672 60012 18682
rect 60076 18678 61124 18682
rect 60132 18674 61124 18678
rect 58964 18590 59956 18672
rect 60132 18598 61134 18674
rect 56440 18438 56778 18477
rect 56786 18443 58712 18477
rect 54469 18427 56778 18438
rect 57235 18431 57236 18432
rect 57248 18431 57282 18443
rect 57294 18431 57295 18432
rect 57236 18430 57237 18431
rect 57248 18430 57294 18431
rect 54480 18415 56778 18427
rect 54469 18404 56778 18415
rect 54496 18260 54530 18404
rect 56440 18335 56778 18404
rect 54569 18324 56036 18335
rect 56146 18324 56778 18335
rect 57248 18327 57293 18430
rect 57482 18422 58136 18443
rect 58551 18431 58552 18432
rect 58564 18431 58598 18443
rect 58552 18430 58553 18431
rect 57884 18338 57964 18422
rect 57906 18327 57951 18338
rect 58564 18327 58609 18431
rect 54580 18315 56778 18324
rect 54580 18290 58583 18315
rect 56440 18268 58583 18290
rect 43666 18228 56014 18260
rect 43666 18222 43684 18228
rect 42958 18160 42992 18190
rect 43616 18160 43650 18194
rect 43742 18160 43776 18228
rect 43844 18164 43878 18228
rect 44068 18226 56014 18228
rect 44068 18180 50506 18226
rect 52056 18180 52090 18226
rect 44068 18172 51954 18180
rect 51988 18172 54272 18180
rect 43844 18160 43916 18164
rect 44068 18160 50506 18172
rect 41624 18146 50506 18160
rect 51916 18146 52019 18158
rect 52056 18146 52090 18172
rect 54394 18146 54428 18226
rect 55326 18172 55878 18180
rect 54465 18157 54568 18158
rect 54465 18150 55326 18157
rect 54458 18146 55326 18150
rect 55828 18146 55839 18157
rect 41624 18138 54272 18146
rect 54360 18138 55844 18146
rect 41624 18126 52004 18138
rect 41424 17564 41564 17624
rect 41228 17478 41564 17564
rect 41228 17176 41562 17478
rect 41318 15873 41352 17176
rect 41320 15861 41352 15873
rect 41290 15857 41352 15861
rect 41290 15814 41337 15857
rect 41354 15835 41388 17176
rect 41354 15823 41386 15835
rect 32190 15780 41337 15814
rect 32190 15764 32226 15780
rect 32736 15712 36360 15780
rect 36457 15712 36491 15780
rect 36571 15712 36605 15780
rect 36726 15712 37148 15780
rect 37202 15712 37624 15780
rect 37772 15712 38590 15780
rect 39203 15712 39248 15780
rect 39861 15712 39895 15780
rect 39975 15712 40009 15780
rect 41432 15712 41466 17176
rect 32126 15678 32134 15712
rect 32168 15678 41400 15712
rect 41434 15678 41466 15712
rect 32736 15436 36360 15678
rect 36457 15654 36491 15678
rect 36571 15654 36605 15678
rect 36726 15654 37148 15678
rect 37202 15654 37624 15678
rect 36378 15644 37624 15654
rect 36457 15483 36491 15644
rect 36726 15632 37148 15644
rect 37202 15632 37624 15644
rect 37772 15644 38590 15678
rect 39203 15644 39248 15678
rect 39861 15644 39895 15678
rect 37772 15632 38585 15644
rect 36586 15585 37624 15632
rect 37654 15585 39486 15632
rect 39833 15585 39880 15632
rect 36633 15578 38564 15585
rect 36633 15551 37248 15578
rect 37291 15551 38564 15578
rect 38607 15551 39222 15585
rect 39265 15551 39880 15585
rect 37408 15483 37489 15551
rect 37510 15483 37544 15551
rect 37772 15483 38564 15551
rect 39975 15483 40009 15678
rect 36457 15449 40009 15483
rect 41468 15568 41562 17176
rect 42300 15658 42334 18126
rect 42958 15658 42992 18126
rect 43742 15682 43776 18126
rect 43844 17798 43916 18126
rect 44068 18112 52004 18126
rect 52022 18112 52090 18138
rect 54360 18112 55839 18138
rect 44068 17781 50506 18112
rect 51916 18100 52004 18112
rect 51954 17798 51988 18100
rect 43917 17770 50506 17781
rect 51904 17770 51915 17781
rect 43806 17708 43916 17746
rect 43928 17736 51915 17770
rect 43844 17252 43916 17708
rect 44068 17688 50506 17736
rect 51916 17708 51988 17746
rect 51954 17700 51988 17708
rect 51916 17688 52004 17700
rect 52056 17688 52090 18112
rect 54394 17688 54428 18112
rect 54480 18100 54568 18112
rect 54496 17700 54568 18100
rect 55840 18084 55912 18122
rect 55878 17716 55912 18084
rect 54480 17699 54568 17700
rect 54480 17692 55326 17699
rect 54458 17688 55326 17692
rect 55828 17688 55839 17699
rect 44068 17672 52004 17688
rect 52022 17672 52090 17688
rect 44068 17654 52090 17672
rect 54360 17654 55839 17688
rect 44068 17648 52054 17654
rect 44068 17644 50506 17648
rect 51916 17644 52019 17648
rect 44068 17642 52026 17644
rect 44068 17620 51948 17642
rect 51994 17620 52026 17642
rect 44068 17574 50506 17620
rect 52056 17574 52090 17654
rect 54394 17574 54428 17654
rect 54465 17642 54568 17654
rect 55980 17574 56014 18226
rect 56440 18234 57267 18268
rect 57310 18234 57925 18268
rect 57968 18234 58583 18268
rect 56440 18166 56778 18234
rect 58678 18166 58712 18443
rect 56440 18132 58712 18166
rect 59054 18477 59088 18590
rect 59168 18490 59213 18590
rect 59826 18490 59871 18590
rect 60484 18584 60529 18598
rect 59168 18489 59214 18490
rect 59814 18489 59815 18490
rect 59826 18489 59872 18490
rect 59168 18477 59202 18489
rect 59214 18488 59215 18489
rect 59813 18488 59814 18489
rect 59214 18477 59814 18488
rect 59826 18477 59860 18489
rect 59872 18488 59873 18489
rect 60392 18488 60422 18570
rect 60448 18488 60450 18570
rect 60472 18489 60473 18490
rect 60471 18488 60472 18489
rect 59872 18477 60472 18488
rect 60480 18488 60800 18584
rect 61108 18488 61134 18598
rect 60480 18477 61134 18488
rect 61136 18483 61140 18570
rect 61142 18477 61176 19101
rect 61256 18477 61290 19101
rect 61292 18477 64916 19124
rect 59054 18443 64916 18477
rect 59054 18172 59088 18443
rect 59168 18431 59202 18443
rect 59214 18431 59215 18432
rect 59813 18431 59814 18432
rect 59826 18431 59860 18443
rect 59872 18431 59873 18432
rect 59168 18430 59214 18431
rect 59814 18430 59815 18431
rect 59826 18430 59872 18431
rect 59168 18333 59213 18430
rect 59826 18333 59871 18430
rect 60392 18366 60422 18437
rect 60448 18380 60450 18437
rect 60471 18431 60472 18432
rect 60472 18430 60473 18431
rect 60480 18406 60800 18443
rect 60392 18324 60450 18366
rect 60484 18333 60529 18406
rect 60556 18380 60588 18394
rect 60556 18324 60588 18366
rect 61108 18321 61134 18443
rect 61136 18380 61140 18437
rect 61142 18333 61176 18443
rect 61142 18321 61168 18333
rect 59183 18317 61168 18321
rect 59183 18274 61161 18317
rect 59230 18240 59845 18274
rect 59888 18240 60503 18274
rect 60546 18240 61161 18274
rect 61256 18172 61290 18443
rect 59054 18138 61290 18172
rect 56440 18096 56778 18132
rect 56555 17948 56778 18096
rect 56555 17912 57456 17948
rect 44068 17540 56014 17574
rect 56500 17878 57456 17912
rect 43844 17140 43878 17252
rect 44068 17112 50506 17540
rect 51920 17170 51938 17196
rect 51948 17142 51966 17196
rect 43928 17098 50506 17112
rect 43806 17050 43878 17088
rect 43928 17078 51904 17098
rect 43844 16482 43878 17050
rect 44068 17064 50506 17078
rect 52056 17064 52090 17540
rect 54394 17064 54428 17540
rect 44068 17030 54606 17064
rect 44068 17016 51322 17030
rect 44068 17000 50506 17016
rect 44068 16962 51916 17000
rect 51954 16962 51988 17030
rect 52056 16962 52090 17030
rect 44068 16928 52090 16962
rect 44068 16454 50506 16928
rect 51915 16890 51916 16891
rect 51954 16890 51988 16928
rect 51916 16889 51917 16890
rect 51954 16582 52026 16890
rect 51954 16482 51988 16582
rect 51904 16454 51915 16465
rect 43806 16392 43878 16430
rect 43928 16420 51915 16454
rect 43844 15824 43878 16392
rect 44068 16052 50506 16420
rect 51916 16392 51988 16430
rect 51916 16090 51917 16091
rect 51915 16089 51916 16090
rect 51954 16052 51988 16392
rect 52056 16052 52090 16928
rect 44068 16018 52090 16052
rect 44068 15950 50506 16018
rect 51954 15950 51988 16018
rect 52056 15950 52090 16018
rect 54394 15950 54428 17030
rect 54430 16928 54462 16962
rect 54480 16890 54488 17020
rect 54496 16890 54530 17030
rect 54465 16878 54530 16890
rect 54458 16102 54530 16878
rect 54465 16090 54530 16102
rect 54430 16018 54462 16052
rect 54480 16002 54488 16090
rect 54496 15950 54530 16090
rect 54572 15963 54606 17030
rect 56500 16598 56534 17878
rect 56555 16598 57456 17878
rect 56500 16564 57456 16598
rect 56555 16528 57456 16564
rect 57654 16528 58646 17948
rect 56555 16515 56778 16528
rect 56555 16457 56796 16515
rect 56555 15963 56778 16457
rect 58758 16286 58764 17968
rect 58786 16314 58820 17968
rect 54569 15952 55936 15963
rect 56458 15952 56778 15963
rect 54572 15950 56778 15952
rect 44068 15918 56778 15950
rect 58964 15936 59956 17956
rect 60132 15944 61124 17964
rect 44068 15916 54606 15918
rect 44068 15844 50506 15916
rect 44068 15824 51324 15844
rect 44068 15796 50506 15824
rect 43928 15762 50506 15796
rect 44068 15682 50506 15762
rect 52056 15744 52090 15916
rect 43742 15660 50506 15682
rect 43742 15648 52090 15660
rect 42842 15634 43780 15642
rect 42842 15620 42950 15634
rect 44068 15612 50506 15648
rect 42808 15586 42946 15608
rect 43004 15600 43604 15608
rect 43662 15600 43814 15608
rect 43728 15574 43890 15576
rect 41468 15472 41556 15568
rect 43766 15536 43852 15538
rect 44068 15518 45116 15612
rect 45152 15608 45314 15612
rect 45482 15606 50506 15612
rect 54394 15606 54428 15916
rect 56555 15857 56778 15918
rect 56555 15845 56796 15857
rect 61292 15845 64916 18443
rect 56555 15838 64916 15845
rect 54449 15811 64916 15838
rect 54449 15804 56796 15811
rect 56555 15799 56796 15804
rect 56555 15661 56778 15799
rect 61292 15661 64916 15811
rect 64923 15731 64934 19215
rect 65164 16808 65247 19539
rect 65314 19532 65348 19566
rect 65966 19538 66012 19600
rect 66022 19594 66040 19600
rect 65972 19532 66006 19538
rect 66008 19532 66012 19538
rect 66630 19532 66664 19600
rect 67288 19532 67322 19600
rect 67754 19552 67830 19600
rect 67754 19532 67832 19552
rect 67834 19532 67892 19600
rect 67912 19594 67930 19600
rect 67940 19538 67986 19600
rect 67996 19594 68014 19600
rect 67940 19532 67944 19538
rect 67946 19532 67980 19538
rect 68484 19532 68485 19600
rect 68570 19594 68588 19600
rect 68598 19566 68638 19600
rect 68604 19532 68638 19566
rect 65296 19507 68650 19532
rect 68656 19507 68672 19532
rect 68692 19507 68712 19698
rect 65296 19506 68712 19507
rect 65296 19498 68650 19506
rect 68656 19498 68672 19506
rect 66008 17027 66012 19498
rect 66630 17039 66664 19498
rect 67754 19468 67832 19498
rect 67834 19468 67892 19498
rect 67833 18992 67838 19256
rect 67833 18896 67844 18992
rect 67940 18832 67944 19498
rect 67874 18264 67984 18832
rect 67940 17240 67944 18264
rect 67918 17032 67944 17240
rect 67940 17027 67944 17032
rect 68718 16940 68752 23768
rect 68958 18612 69256 18628
rect 68974 18372 69256 18612
rect 45190 15570 45276 15582
rect 45482 15578 56014 15606
rect 45630 15572 56014 15578
rect 45152 15518 45176 15560
rect 45190 15518 45214 15570
rect 37408 15436 37489 15449
rect 35178 15058 35212 15436
rect 35238 15058 35361 15436
rect 37408 15071 37442 15436
rect 37361 15058 37442 15071
rect 37510 15058 37544 15449
rect 37772 15058 38564 15449
rect 41468 15436 41538 15472
rect 44068 15458 45374 15518
rect 45630 15458 50506 15572
rect 54394 15492 54428 15572
rect 54465 15503 54568 15504
rect 54465 15496 55326 15503
rect 54458 15492 55326 15496
rect 55828 15492 55839 15503
rect 54360 15458 55839 15492
rect 55844 15468 55946 15470
rect 55840 15462 55946 15468
rect 45812 15436 45816 15458
rect 45840 15452 45844 15458
rect 32168 15024 41400 15058
rect 32180 15003 32214 15024
rect 35178 15003 35212 15024
rect 32180 14956 35212 15003
rect 32180 12619 32214 14956
rect 32242 14922 35212 14956
rect 35178 13914 35212 14922
rect 35238 15003 35361 15024
rect 35238 14956 36338 15003
rect 37408 14956 37442 15024
rect 37510 14956 37544 15024
rect 37772 15003 38564 15024
rect 41354 15003 41388 15024
rect 37654 14956 39486 15003
rect 41326 14956 41388 15003
rect 35238 14922 41388 14956
rect 35238 14598 35361 14922
rect 35238 14056 35314 14598
rect 37408 14056 37442 14922
rect 35238 14040 35306 14056
rect 35238 13914 35272 14040
rect 37349 14028 37360 14039
rect 35373 13994 37360 14028
rect 37510 13914 37544 14922
rect 35178 13880 37544 13914
rect 35238 12619 35272 13880
rect 37772 13820 38564 14922
rect 38296 12619 38330 13820
rect 41354 12619 41388 14922
rect 32180 12572 33498 12619
rect 35210 12606 35272 12619
rect 38268 12606 38330 12619
rect 35210 12578 35278 12606
rect 38268 12578 38336 12606
rect 35204 12572 35278 12578
rect 35288 12572 35306 12578
rect 38262 12572 38336 12578
rect 38346 12572 38364 12578
rect 38580 12572 39494 12619
rect 41326 12578 41388 12619
rect 41320 12572 41388 12578
rect 32180 12504 32220 12572
rect 32230 12538 35278 12572
rect 35284 12538 38336 12572
rect 38342 12538 41388 12572
rect 32230 12532 32248 12538
rect 35204 12532 35222 12538
rect 35232 12504 35278 12538
rect 35288 12532 35306 12538
rect 38262 12532 38280 12538
rect 38290 12504 38336 12538
rect 38346 12532 38364 12538
rect 41320 12532 41338 12538
rect 41348 12504 41388 12538
rect 32180 12470 32214 12504
rect 35238 12470 35272 12504
rect 38296 12470 38330 12504
rect 41354 12470 41388 12504
rect 32162 12436 41422 12470
rect 41468 10842 41502 15436
rect 41526 14598 41536 15436
rect 44068 15100 44468 15136
rect 44518 15100 44552 15132
rect 44713 15100 44889 15134
rect 45050 15100 45084 15132
rect 45630 15100 50506 15136
rect 44068 15066 50506 15100
rect 44068 14824 44468 15066
rect 44518 14986 44552 15066
rect 44620 15014 44654 15024
rect 44948 15014 44982 15024
rect 44589 14986 44701 14998
rect 44901 14986 45013 14998
rect 45050 14986 45084 15066
rect 45094 14998 45176 15024
rect 44518 14960 45214 14986
rect 44518 14952 45084 14960
rect 44518 14872 44552 14952
rect 45050 14950 45084 14952
rect 44896 14946 45084 14950
rect 45050 14872 45084 14946
rect 44518 14838 45084 14872
rect 45630 14920 50506 15066
rect 54394 15034 54428 15458
rect 54480 15446 54568 15458
rect 54496 15294 54568 15446
rect 55840 15442 55912 15462
rect 55840 15430 55918 15442
rect 55872 15406 55918 15430
rect 55872 15396 55912 15406
rect 55878 15278 55912 15396
rect 54569 15266 55326 15277
rect 55840 15266 55928 15278
rect 54458 15204 54568 15242
rect 54580 15232 55928 15266
rect 54496 15046 54568 15204
rect 55326 15198 55330 15228
rect 55840 15220 55928 15232
rect 55878 15096 55912 15220
rect 55872 15070 55912 15096
rect 55872 15050 55918 15070
rect 54480 15045 54568 15046
rect 54480 15038 55330 15045
rect 54458 15034 55330 15038
rect 55828 15034 55839 15045
rect 54360 15000 55839 15034
rect 54394 14920 54428 15000
rect 54465 14988 54568 15000
rect 55980 14920 56014 15572
rect 69367 15545 69401 26373
rect 69531 26327 69598 26340
rect 70046 26327 70123 26340
rect 70189 26327 70256 26340
rect 70704 26327 70781 26340
rect 70847 26327 70918 26340
rect 71366 26327 71439 26340
rect 71505 26327 71588 26340
rect 72036 26327 72097 26340
rect 72163 26327 72240 26340
rect 72688 26327 72755 26340
rect 72113 23815 72147 26274
rect 69469 23781 72817 23815
rect 69481 23747 69515 23781
rect 70139 23760 70173 23781
rect 70797 23760 70831 23781
rect 71455 23760 71489 23781
rect 72113 23760 72147 23781
rect 72771 23760 72805 23781
rect 70111 23747 70173 23760
rect 70769 23747 70831 23760
rect 71427 23747 71489 23760
rect 72085 23747 72147 23760
rect 69481 23645 69521 23747
rect 70111 23719 70179 23747
rect 70769 23719 70837 23747
rect 71427 23719 71495 23747
rect 72085 23719 72153 23747
rect 72743 23719 72805 23760
rect 69531 23713 69549 23719
rect 70105 23713 70179 23719
rect 70189 23713 70207 23719
rect 70763 23713 70837 23719
rect 70847 23713 70865 23719
rect 71421 23713 71495 23719
rect 71505 23713 71523 23719
rect 72079 23713 72153 23719
rect 72163 23713 72181 23719
rect 72737 23713 72805 23719
rect 69527 23679 70179 23713
rect 70185 23679 70837 23713
rect 70843 23679 71495 23713
rect 71501 23679 72153 23713
rect 72159 23679 72805 23713
rect 69531 23673 69549 23679
rect 70105 23673 70123 23679
rect 70133 23645 70179 23679
rect 70189 23673 70207 23679
rect 70763 23673 70781 23679
rect 70791 23645 70837 23679
rect 70847 23673 70865 23679
rect 71421 23673 71439 23679
rect 71449 23645 71495 23679
rect 71505 23673 71523 23679
rect 72079 23673 72097 23679
rect 72107 23645 72153 23679
rect 72163 23673 72181 23679
rect 72737 23673 72755 23679
rect 72765 23645 72805 23679
rect 69481 18273 69515 23645
rect 70139 18286 70173 23645
rect 70797 18286 70831 23645
rect 71455 18286 71489 23645
rect 72113 18286 72147 23645
rect 72771 18286 72805 23645
rect 70111 18273 70173 18286
rect 70769 18273 70831 18286
rect 71427 18273 71489 18286
rect 72085 18273 72147 18286
rect 69481 18171 69521 18273
rect 70111 18245 70179 18273
rect 70769 18245 70837 18273
rect 71427 18245 71495 18273
rect 72085 18245 72153 18273
rect 72743 18245 72805 18286
rect 69531 18239 69549 18245
rect 70105 18239 70179 18245
rect 70189 18239 70207 18245
rect 70763 18239 70837 18245
rect 70847 18239 70865 18245
rect 71421 18239 71495 18245
rect 71505 18239 71523 18245
rect 72079 18239 72153 18245
rect 72163 18239 72181 18245
rect 72737 18239 72805 18245
rect 69527 18205 70179 18239
rect 70185 18205 70837 18239
rect 70843 18205 71495 18239
rect 71501 18205 72153 18239
rect 72159 18205 72805 18239
rect 69531 18199 69549 18205
rect 70105 18199 70123 18205
rect 70133 18171 70179 18205
rect 70189 18199 70207 18205
rect 70763 18199 70781 18205
rect 70791 18171 70837 18205
rect 70847 18199 70865 18205
rect 71421 18199 71439 18205
rect 71449 18171 71495 18205
rect 71505 18199 71523 18205
rect 72079 18199 72097 18205
rect 72107 18171 72153 18205
rect 72163 18199 72181 18205
rect 72737 18199 72755 18205
rect 72765 18171 72805 18205
rect 69481 18137 69515 18171
rect 70139 18137 70173 18171
rect 70797 18137 70831 18171
rect 71455 18137 71489 18171
rect 72113 18137 72147 18171
rect 72771 18137 72805 18171
rect 69463 18103 72817 18137
rect 72823 18103 72839 18137
rect 72885 15545 72919 26373
rect 74303 25167 74337 31839
rect 74417 31777 74451 31938
rect 75075 31926 75109 31938
rect 75733 31926 75767 31938
rect 74453 31811 74457 31913
rect 74481 31879 74485 31885
rect 75061 31879 75109 31926
rect 75719 31879 75767 31926
rect 74477 31845 74485 31879
rect 74493 31845 75109 31879
rect 75135 31845 75143 31879
rect 75151 31845 75767 31879
rect 74481 31839 74485 31845
rect 75063 31829 75109 31845
rect 75721 31829 75767 31845
rect 75075 31777 75109 31829
rect 75733 31777 75767 31829
rect 75769 31811 75773 31913
rect 76314 31885 76316 32982
rect 76342 31885 76344 32954
rect 76391 31938 76439 33242
rect 77049 31938 77097 33242
rect 76391 31926 76425 31938
rect 77049 31926 77083 31938
rect 75797 31879 75801 31885
rect 76377 31879 76425 31926
rect 77035 31879 77083 31926
rect 75793 31845 75801 31879
rect 75809 31845 76425 31879
rect 76451 31845 76459 31879
rect 76467 31845 77083 31879
rect 75797 31839 75801 31845
rect 76314 31832 76316 31839
rect 76342 31804 76344 31839
rect 76379 31829 76425 31845
rect 77037 31829 77083 31845
rect 76391 31777 76425 31829
rect 77049 31777 77083 31829
rect 77085 31811 77089 31913
rect 77636 31885 77638 32952
rect 77664 31885 77666 32924
rect 77707 31938 77755 33242
rect 77707 31926 77741 31938
rect 77113 31879 77117 31885
rect 77693 31879 77741 31926
rect 77109 31845 77117 31879
rect 77125 31845 77741 31879
rect 77113 31839 77117 31845
rect 77636 31832 77638 31839
rect 77664 31804 77666 31839
rect 77695 31829 77741 31845
rect 77707 31777 77741 31829
rect 77821 31839 77869 33341
rect 79374 31862 79422 33346
rect 79502 33356 79536 33408
rect 80118 33374 80156 33378
rect 79502 33268 79548 33356
rect 80118 33340 80158 33374
rect 79550 33306 80158 33340
rect 80126 33300 80130 33306
rect 80154 33272 80158 33306
rect 80160 33356 80194 33408
rect 80160 33268 80206 33356
rect 80776 33340 80814 33378
rect 80208 33306 80814 33340
rect 80818 33346 80884 33408
rect 80908 33346 80912 33408
rect 80818 33300 80864 33346
rect 81434 33340 81472 33378
rect 80866 33306 81472 33340
rect 81476 33356 81510 33408
rect 82070 33378 82096 33408
rect 82098 33378 82168 33408
rect 82070 33356 82168 33378
rect 82750 33374 82788 33378
rect 79502 33256 79536 33268
rect 80135 33256 80148 33267
rect 80160 33256 80194 33268
rect 80793 33256 80806 33267
rect 80818 33256 80884 33300
rect 79488 31952 79536 33256
rect 74405 31743 77753 31777
rect 77821 26759 77855 31839
rect 77821 26510 77891 26759
rect 74402 25035 77891 26510
rect 79374 26505 79408 31862
rect 79488 31800 79522 31952
rect 79524 31834 79528 31936
rect 80074 31908 80082 32720
rect 80102 31908 80110 32692
rect 80146 31952 80194 33256
rect 80804 32242 80884 33256
rect 80146 31940 80180 31952
rect 80804 31940 80858 32242
rect 80908 32214 80912 33300
rect 81476 33268 81522 33356
rect 82070 33346 82180 33356
rect 82092 33340 82130 33346
rect 81524 33306 82130 33340
rect 82134 33300 82180 33346
rect 82750 33340 82790 33374
rect 82182 33306 82790 33340
rect 82758 33300 82762 33306
rect 81451 33256 81464 33267
rect 81476 33256 81510 33268
rect 81462 31952 81510 33256
rect 82070 32178 82096 33300
rect 82098 33268 82180 33300
rect 82786 33272 82790 33306
rect 82098 32206 82168 33268
rect 82767 33256 82780 33267
rect 82792 33256 82826 33408
rect 82906 33346 82940 36356
rect 90876 36352 90896 36472
rect 90904 36346 90924 36500
rect 96108 36302 96128 36456
rect 96136 36308 96156 36428
rect 83558 34992 91534 35026
rect 84140 34410 85244 34430
rect 82086 32132 82096 32178
rect 82114 32132 82168 32206
rect 82702 32132 82708 32704
rect 82730 32132 82736 32676
rect 82120 31994 82168 32132
rect 81462 31940 81496 31952
rect 79552 31902 79556 31908
rect 80132 31902 80180 31940
rect 80790 31908 80844 31940
rect 80790 31902 80838 31908
rect 79548 31868 79556 31902
rect 79564 31868 80180 31902
rect 80206 31868 80214 31902
rect 80222 31868 80838 31902
rect 79552 31862 79556 31868
rect 80074 31856 80082 31862
rect 80102 31828 80110 31862
rect 80134 31852 80180 31868
rect 80792 31862 80838 31868
rect 80840 31862 80844 31908
rect 80868 31902 80872 31908
rect 81448 31902 81496 31940
rect 82086 31908 82096 31994
rect 82114 31952 82168 31994
rect 82114 31940 82154 31952
rect 82106 31902 82154 31940
rect 80864 31868 80872 31902
rect 80880 31868 81496 31902
rect 81522 31868 81530 31902
rect 81538 31868 82154 31902
rect 80868 31862 80872 31868
rect 80792 31852 80844 31862
rect 81450 31852 81496 31868
rect 80146 31800 80180 31852
rect 80804 31806 80844 31852
rect 80804 31800 80838 31806
rect 81462 31800 81496 31852
rect 82086 31800 82096 31862
rect 82108 31852 82154 31868
rect 82114 31800 82154 31852
rect 82156 31834 82160 31936
rect 82702 31908 82708 31994
rect 82730 31908 82736 31994
rect 82778 31952 82826 33256
rect 82778 31940 82812 31952
rect 82184 31902 82188 31908
rect 82764 31902 82812 31940
rect 82180 31868 82188 31902
rect 82196 31868 82812 31902
rect 82184 31862 82188 31868
rect 82702 31850 82708 31862
rect 82730 31828 82736 31862
rect 82766 31852 82812 31868
rect 82778 31800 82812 31852
rect 82892 31862 82940 33346
rect 83336 33332 86647 33473
rect 91618 33442 91620 33476
rect 83219 33301 86647 33332
rect 83336 33298 86647 33301
rect 83139 32920 83162 33282
rect 83185 33267 86647 33298
rect 83167 32920 83190 33254
rect 83336 32280 86647 33267
rect 88130 33408 91665 33442
rect 88130 33052 88164 33408
rect 88874 33340 88912 33378
rect 89532 33340 89570 33378
rect 90190 33340 90228 33378
rect 90848 33340 90886 33378
rect 91506 33340 91544 33378
rect 88306 33306 88912 33340
rect 88964 33306 89570 33340
rect 89622 33306 90228 33340
rect 90280 33306 90886 33340
rect 90938 33306 91544 33340
rect 91584 33296 91602 33306
rect 88233 33256 88278 33267
rect 88891 33256 88936 33267
rect 89549 33256 89594 33267
rect 90207 33256 90252 33267
rect 90865 33256 90910 33267
rect 88244 33052 88278 33256
rect 88289 33064 88290 33065
rect 88890 33064 88891 33065
rect 88290 33063 88291 33064
rect 88889 33063 88890 33064
rect 88902 33052 88936 33256
rect 88947 33064 88948 33065
rect 89548 33064 89549 33065
rect 88948 33063 88949 33064
rect 89547 33063 89548 33064
rect 89560 33052 89594 33256
rect 89605 33064 89606 33065
rect 90206 33064 90207 33065
rect 89606 33063 89607 33064
rect 90205 33063 90206 33064
rect 90218 33052 90252 33256
rect 90263 33064 90264 33065
rect 90864 33064 90865 33065
rect 90264 33063 90265 33064
rect 90863 33063 90864 33064
rect 90876 33052 90910 33256
rect 91500 33144 91518 33296
rect 91578 33294 91602 33296
rect 91550 33268 91568 33272
rect 91578 33268 91606 33294
rect 91528 33267 91606 33268
rect 91523 33256 91606 33267
rect 91528 33116 91606 33256
rect 91534 33080 91606 33116
rect 91534 33068 91602 33080
rect 90921 33064 90922 33065
rect 91522 33064 91523 33065
rect 90922 33063 90923 33064
rect 91521 33063 91522 33064
rect 91534 33052 91580 33068
rect 91584 33064 91602 33068
rect 91614 33064 91618 33408
rect 91648 33080 91665 33408
rect 88096 33049 91580 33052
rect 88096 33040 91574 33049
rect 88096 33030 91568 33040
rect 91648 33037 91652 33080
rect 88096 33028 91574 33030
rect 88096 33018 91580 33028
rect 88130 32394 88164 33018
rect 88244 32394 88278 33018
rect 88290 33006 88291 33007
rect 88889 33006 88890 33007
rect 88289 33005 88290 33006
rect 88890 33005 88891 33006
rect 88289 32406 88290 32407
rect 88890 32406 88891 32407
rect 88290 32405 88291 32406
rect 88889 32405 88890 32406
rect 88902 32394 88936 33018
rect 88948 33006 88949 33007
rect 89547 33006 89548 33007
rect 88947 33005 88948 33006
rect 89548 33005 89549 33006
rect 88947 32406 88948 32407
rect 89548 32406 89549 32407
rect 88948 32405 88949 32406
rect 89547 32405 89548 32406
rect 89560 32394 89594 33018
rect 89606 33006 89607 33007
rect 90205 33006 90206 33007
rect 89605 33005 89606 33006
rect 90206 33005 90207 33006
rect 89605 32406 89606 32407
rect 90206 32406 90207 32407
rect 89606 32405 89607 32406
rect 90205 32405 90206 32406
rect 90218 32394 90252 33018
rect 90264 33006 90265 33007
rect 90863 33006 90864 33007
rect 90263 33005 90264 33006
rect 90864 33005 90865 33006
rect 90263 32406 90264 32407
rect 90864 32406 90865 32407
rect 90264 32405 90265 32406
rect 90863 32405 90864 32406
rect 90876 32394 90910 33018
rect 90922 33006 90923 33007
rect 91521 33006 91522 33007
rect 90921 33005 90922 33006
rect 91522 33005 91523 33006
rect 91534 33002 91580 33018
rect 91584 33002 91602 33006
rect 91534 32990 91602 33002
rect 91534 32940 91606 32990
rect 90921 32406 90922 32407
rect 91522 32406 91523 32407
rect 90922 32405 90923 32406
rect 91521 32405 91522 32406
rect 91534 32394 91580 32940
rect 91584 32422 91606 32940
rect 91584 32406 91602 32422
rect 91614 32406 91618 33006
rect 91648 32422 91665 33037
rect 88096 32391 91580 32394
rect 88096 32360 91568 32391
rect 91648 32372 91652 32422
rect 88130 32280 88164 32360
rect 88244 32280 88278 32360
rect 88902 32280 88936 32360
rect 89560 32280 89594 32360
rect 90218 32280 90252 32360
rect 90876 32280 90910 32360
rect 91534 32280 91568 32360
rect 83336 32246 91580 32280
rect 91648 32246 91658 32314
rect 91686 32280 91720 33496
rect 113115 33045 113149 39409
rect 115861 35962 115895 39310
rect 115861 35610 115901 35962
rect 113229 33141 113263 33175
rect 113887 33141 113921 33175
rect 114545 33141 114579 33175
rect 115203 33141 115237 33175
rect 115861 33141 115895 35610
rect 116519 33437 116553 33471
rect 116633 33437 116667 39409
rect 118958 33473 118992 39324
rect 118150 33437 119557 33473
rect 121590 33442 121624 33476
rect 121704 33442 121738 39414
rect 115969 33403 119557 33437
rect 115969 33141 116003 33403
rect 116098 33335 116565 33382
rect 116145 33301 116565 33335
rect 116507 33254 116565 33301
rect 116072 33242 116128 33253
rect 116083 33141 116128 33242
rect 116519 33175 116564 33254
rect 116519 33141 116573 33175
rect 116633 33141 116667 33403
rect 118150 33182 119557 33403
rect 113179 33107 113183 33141
rect 113195 33107 116667 33141
rect 83336 32210 86647 32246
rect 79476 31766 82824 31800
rect 80146 26505 80180 31766
rect 80804 26505 80838 31766
rect 82086 31398 82096 31766
rect 82114 31398 82152 31766
rect 81528 30892 82120 30906
rect 82154 30892 82308 30906
rect 81562 30858 82120 30872
rect 82154 30858 82308 30872
rect 82086 28938 82096 30210
rect 82114 28938 82152 30210
rect 82086 27438 82096 27750
rect 82114 27438 82152 27750
rect 80846 26512 80870 26972
rect 80852 26505 80870 26512
rect 74438 15568 74472 25035
rect 74540 23786 77888 23820
rect 74552 18296 74586 23786
rect 75210 23756 75244 23786
rect 75868 23756 75902 23786
rect 76526 23756 76560 23786
rect 77184 23756 77218 23786
rect 77842 23756 77876 23786
rect 75182 23718 75244 23756
rect 75840 23718 75902 23756
rect 76498 23718 76560 23756
rect 77156 23718 77218 23756
rect 77814 23718 77876 23756
rect 74598 23684 75244 23718
rect 75256 23684 75902 23718
rect 75914 23684 76560 23718
rect 76572 23684 77218 23718
rect 77230 23684 77876 23718
rect 74618 19462 74624 19718
rect 74646 19490 74652 19690
rect 74618 19062 74624 19318
rect 74646 19090 74652 19290
rect 75210 18300 75244 23684
rect 75868 18300 75902 23684
rect 76526 18300 76560 23684
rect 77184 18300 77218 23684
rect 77842 18300 77876 23684
rect 75182 18296 75244 18300
rect 75840 18296 75902 18300
rect 76498 18296 76560 18300
rect 77156 18296 77218 18300
rect 74552 18194 74592 18296
rect 75182 18268 75250 18296
rect 75840 18268 75908 18296
rect 76498 18268 76566 18296
rect 77156 18268 77224 18296
rect 77814 18268 77876 18300
rect 74602 18262 74620 18268
rect 75176 18262 75250 18268
rect 75260 18262 75278 18268
rect 75834 18262 75908 18268
rect 75918 18262 75936 18268
rect 76492 18262 76566 18268
rect 76576 18262 76594 18268
rect 77150 18262 77224 18268
rect 77234 18262 77252 18268
rect 77808 18262 77876 18268
rect 74598 18228 75250 18262
rect 75256 18228 75908 18262
rect 75914 18228 76566 18262
rect 76572 18228 77224 18262
rect 77230 18228 77876 18262
rect 74602 18222 74620 18228
rect 75176 18222 75194 18228
rect 75204 18194 75250 18228
rect 75260 18222 75278 18228
rect 75834 18222 75852 18228
rect 75862 18194 75908 18228
rect 75918 18222 75936 18228
rect 76492 18222 76510 18228
rect 76520 18194 76566 18228
rect 76576 18222 76594 18228
rect 77150 18222 77168 18228
rect 77178 18194 77224 18228
rect 77234 18222 77252 18228
rect 77808 18222 77826 18228
rect 77836 18194 77876 18228
rect 74552 18160 74586 18194
rect 75210 18160 75244 18194
rect 75868 18160 75902 18194
rect 76526 18160 76560 18194
rect 77184 18160 77218 18194
rect 77842 18160 77876 18194
rect 74534 18126 77910 18160
rect 75210 15862 75244 18126
rect 76540 17252 77328 17270
rect 76540 17140 76560 17252
rect 77184 17236 77232 17252
rect 76574 17202 77294 17236
rect 75178 15828 75244 15862
rect 75868 15828 75902 15862
rect 75116 15794 76264 15828
rect 75116 15506 75150 15794
rect 75210 15690 75244 15794
rect 75868 15714 75902 15794
rect 76078 15714 76089 15725
rect 75180 15668 75252 15690
rect 75302 15680 76089 15714
rect 75855 15668 75856 15669
rect 75180 15652 75256 15668
rect 75856 15667 75857 15668
rect 75868 15658 75902 15680
rect 75914 15668 75915 15669
rect 75913 15667 75914 15668
rect 76090 15652 76162 15690
rect 75198 15646 75256 15652
rect 75289 15646 75290 15647
rect 76090 15646 76091 15647
rect 75202 15642 75252 15646
rect 75290 15645 75291 15646
rect 75184 15608 75194 15614
rect 75202 15608 75258 15642
rect 75260 15608 75286 15614
rect 75840 15608 75878 15646
rect 76089 15645 76090 15646
rect 76128 15608 76162 15652
rect 76230 15608 76264 15794
rect 76574 15642 76608 17202
rect 77118 17134 77156 17172
rect 76750 17100 77156 17134
rect 77196 17100 77218 17164
rect 77150 17061 77180 17066
rect 76677 17050 76722 17061
rect 77135 17050 77180 17061
rect 76688 15646 76722 17050
rect 77146 15646 77180 17050
rect 77184 15646 77218 17100
rect 76554 15608 76608 15642
rect 75180 15574 75198 15608
rect 75202 15574 75878 15608
rect 75930 15574 76264 15608
rect 75184 15568 75194 15574
rect 75202 15558 75258 15574
rect 75260 15568 75286 15574
rect 75212 15540 75258 15558
rect 75218 15506 75252 15540
rect 76128 15506 76162 15574
rect 76230 15506 76264 15574
rect 76574 15506 76608 15608
rect 76676 15608 76734 15646
rect 77134 15642 77218 15646
rect 77134 15608 77190 15642
rect 77230 15608 77252 17164
rect 76676 15574 77190 15608
rect 76676 15558 76734 15574
rect 77134 15558 77172 15574
rect 76676 15543 76691 15558
rect 77260 15506 77294 17202
rect 77956 15568 77990 26378
rect 78123 15545 78157 26373
rect 78287 26327 78354 26340
rect 78802 26327 78879 26340
rect 78945 26327 79012 26340
rect 79338 25058 81711 26505
rect 82246 26284 82248 26992
rect 82892 25190 82926 31862
rect 83135 31790 83136 31876
rect 83173 31752 83174 31914
rect 83342 31872 83764 32210
rect 83818 31872 84240 32210
rect 86577 30727 86611 32210
rect 86612 31830 86647 32084
rect 86866 31368 86901 31830
rect 87322 31658 87424 31670
rect 88130 30763 88164 32246
rect 88206 32018 88220 32104
rect 88244 31980 88258 32142
rect 113083 31235 113149 33045
rect 113225 33055 113229 33073
rect 113225 33039 113275 33055
rect 113286 33045 113304 33060
rect 113314 33045 113332 33058
rect 113827 33039 113874 33086
rect 113883 33055 113887 33073
rect 113883 33039 113933 33055
rect 114485 33045 114532 33086
rect 114476 33039 114532 33045
rect 114541 33055 114545 33073
rect 114541 33039 114591 33055
rect 114606 33045 114612 33048
rect 114634 33045 114640 33058
rect 115143 33039 115190 33086
rect 115199 33055 115203 33073
rect 115199 33039 115249 33055
rect 115801 33045 115848 33086
rect 115861 33073 115895 33107
rect 115796 33039 115848 33045
rect 115857 33055 115895 33073
rect 115900 33055 115901 33107
rect 115969 33086 116003 33107
rect 116083 33104 116128 33107
rect 116519 33104 116564 33107
rect 116083 33086 116117 33104
rect 115857 33039 115907 33055
rect 115969 33039 116016 33086
rect 116083 33055 116130 33086
rect 116071 33039 116130 33055
rect 116459 33039 116506 33086
rect 113229 33005 113874 33039
rect 113887 33005 114532 33039
rect 114545 33005 115190 33039
rect 115203 33005 115848 33039
rect 115861 33005 116506 33039
rect 113229 32958 113275 33005
rect 113185 32946 113203 32958
rect 113229 32946 113263 32958
rect 113185 31322 113263 32946
rect 113286 31658 113304 32999
rect 113314 31630 113332 32999
rect 113887 32958 113933 33005
rect 114476 32999 114497 33005
rect 114504 32971 114525 33005
rect 114545 32958 114591 33005
rect 113844 32946 113875 32957
rect 113887 32946 113921 32958
rect 114502 32946 114533 32957
rect 114545 32946 114579 32958
rect 113784 31322 113794 32680
rect 113812 31322 113822 32652
rect 113855 31322 113921 32946
rect 114513 31322 114579 32946
rect 114606 31646 114612 32999
rect 114634 31618 114640 32999
rect 115203 32958 115249 33005
rect 115796 32999 115813 33005
rect 115824 32971 115841 33005
rect 115861 32999 115907 33005
rect 115861 32958 115932 32999
rect 115160 32946 115191 32957
rect 115203 32946 115237 32958
rect 115818 32946 115849 32957
rect 115861 32946 115895 32958
rect 115094 31322 115114 32686
rect 115122 31322 115142 32658
rect 115171 31322 115237 32946
rect 115829 31337 115895 32946
rect 115900 31624 115932 32958
rect 115900 31337 115901 31624
rect 115956 31596 115960 32999
rect 115829 31322 115901 31337
rect 115969 31322 116003 33005
rect 116071 32958 116129 33005
rect 116083 31322 116117 32958
rect 116519 32957 116553 33104
rect 116476 32946 116553 32957
rect 116487 31334 116553 32946
rect 116487 31322 116532 31334
rect 113185 31318 115550 31322
rect 113185 31308 113231 31318
rect 113244 31308 115550 31318
rect 113185 31284 115550 31308
rect 113083 30832 113117 31235
rect 113185 31173 113231 31284
rect 113244 31275 115550 31284
rect 115817 31275 115876 31322
rect 115969 31275 116016 31322
rect 116083 31275 116130 31322
rect 116487 31275 116534 31322
rect 113291 31241 113902 31275
rect 113937 31272 114560 31275
rect 113949 31241 114560 31272
rect 114607 31241 115218 31275
rect 115265 31241 115876 31275
rect 115923 31241 116534 31275
rect 113843 31225 113889 31241
rect 114501 31225 114547 31241
rect 115159 31225 115205 31241
rect 115817 31235 115863 31241
rect 115817 31225 115869 31235
rect 115829 31179 115869 31225
rect 115829 31173 115863 31179
rect 115969 31173 116003 31241
rect 116083 31173 116117 31241
rect 116487 31173 116521 31241
rect 116601 31173 116667 33107
rect 118118 33146 119557 33182
rect 121040 33408 124496 33442
rect 119616 33146 119650 33180
rect 120274 33146 120308 33180
rect 120932 33146 120966 33180
rect 121040 33146 121074 33408
rect 121590 33371 121628 33378
rect 121590 33356 121636 33371
rect 121578 33340 121636 33356
rect 121216 33306 121636 33340
rect 121578 33268 121636 33306
rect 121143 33256 121188 33267
rect 121154 33146 121188 33256
rect 121590 33180 121624 33268
rect 121590 33146 121644 33180
rect 121704 33146 121738 33408
rect 118118 33112 121738 33146
rect 118118 33082 119557 33112
rect 118118 33040 119594 33082
rect 119610 33060 119624 33106
rect 119610 33050 119662 33060
rect 119612 33044 119662 33050
rect 120214 33044 120252 33082
rect 120270 33060 120274 33078
rect 120270 33044 120320 33060
rect 120872 33044 120910 33082
rect 120928 33060 120932 33078
rect 120970 33060 120972 33112
rect 121040 33082 121074 33112
rect 121154 33082 121188 33112
rect 120928 33044 120978 33060
rect 121040 33044 121078 33082
rect 121154 33060 121192 33082
rect 121142 33044 121200 33060
rect 121530 33044 121568 33082
rect 118118 33010 119596 33040
rect 118118 33004 119568 33010
rect 116698 31596 116704 32948
rect 117464 31940 117502 32140
rect 117520 31912 117530 32168
rect 113185 31139 116667 31173
rect 118118 31298 119557 33004
rect 119574 32976 119596 33010
rect 119616 33010 120252 33044
rect 120274 33010 120910 33044
rect 120932 33010 121568 33044
rect 119574 32971 119588 32976
rect 119616 32972 119662 33010
rect 120274 32972 120320 33010
rect 120932 33004 120978 33010
rect 121040 33004 121074 33010
rect 120932 32972 121004 33004
rect 119573 32960 119604 32971
rect 119616 32960 119650 32972
rect 120231 32960 120262 32971
rect 120274 32960 120308 32972
rect 120889 32960 120920 32971
rect 120932 32960 120966 32972
rect 119574 31638 119650 32960
rect 119578 31348 119650 31638
rect 119578 31336 119618 31348
rect 119572 31298 119622 31336
rect 120174 31304 120190 32236
rect 120202 31304 120218 32236
rect 120242 31348 120308 32960
rect 120318 31546 120338 32236
rect 120900 31360 120966 32960
rect 120970 31602 121004 32972
rect 120970 31360 120972 31602
rect 121026 31546 121074 33004
rect 121142 32972 121200 33010
rect 120242 31336 120276 31348
rect 120900 31336 120972 31360
rect 121040 31336 121074 31546
rect 121154 31336 121188 32972
rect 121590 32971 121624 33112
rect 121547 32960 121624 32971
rect 121558 31348 121624 32960
rect 120230 31298 120280 31336
rect 120888 31304 120940 31336
rect 120888 31298 120938 31304
rect 121040 31298 121078 31336
rect 121154 31298 121192 31336
rect 121558 31332 121603 31348
rect 121558 31298 121596 31332
rect 118118 31264 119622 31298
rect 119678 31264 120280 31298
rect 120336 31264 120938 31298
rect 120994 31264 121596 31298
rect 118118 31196 119557 31264
rect 119572 31248 119618 31264
rect 120230 31248 120276 31264
rect 120888 31258 120934 31264
rect 120888 31248 120940 31258
rect 120900 31202 120940 31248
rect 120900 31196 120934 31202
rect 121040 31196 121074 31264
rect 121154 31200 121188 31264
rect 121558 31200 121592 31264
rect 121154 31196 121199 31200
rect 121558 31196 121603 31200
rect 121672 31196 121738 33112
rect 121774 32692 121790 32694
rect 121768 31588 121790 32692
rect 121812 32596 121846 33256
rect 121812 32514 121912 32596
rect 121774 31304 121790 31504
rect 118118 31162 121738 31196
rect 113197 30832 113231 30866
rect 113855 30832 113889 30866
rect 114513 30832 114547 30866
rect 115171 30832 115205 30866
rect 111898 30798 115354 30832
rect 88094 30727 91718 30763
rect 83377 30693 91718 30727
rect 83377 27209 83411 30693
rect 83831 30692 83865 30693
rect 83831 30619 83871 30692
rect 83890 30619 83899 30664
rect 83831 30613 83865 30619
rect 84489 30613 84523 30693
rect 85147 30613 85181 30693
rect 85805 30613 85839 30693
rect 86463 30613 86497 30693
rect 86577 30613 86611 30693
rect 83432 30551 83513 30598
rect 83572 30579 86611 30613
rect 83831 30573 83865 30579
rect 83818 30567 83819 30568
rect 83819 30566 83820 30567
rect 83479 29983 83513 30551
rect 83831 30508 83871 30573
rect 83877 30567 83878 30568
rect 83876 30566 83877 30567
rect 83890 30536 83899 30573
rect 84476 30567 84477 30568
rect 84477 30566 84478 30567
rect 83819 29967 83820 29968
rect 83818 29966 83819 29967
rect 83831 29955 83865 30508
rect 83876 29967 83877 29968
rect 84477 29967 84478 29968
rect 83877 29966 83878 29967
rect 84476 29966 84477 29967
rect 84489 29955 84523 30579
rect 84535 30567 84536 30568
rect 85134 30567 85135 30568
rect 84534 30566 84535 30567
rect 85135 30566 85136 30567
rect 84534 29967 84535 29968
rect 85135 29967 85136 29968
rect 84535 29966 84536 29967
rect 85134 29966 85135 29967
rect 85147 29955 85181 30579
rect 85193 30567 85194 30568
rect 85792 30567 85793 30568
rect 85192 30566 85193 30567
rect 85793 30566 85794 30567
rect 85192 29967 85193 29968
rect 85793 29967 85794 29968
rect 85193 29966 85194 29967
rect 85792 29966 85793 29967
rect 85805 29955 85839 30579
rect 85851 30567 85852 30568
rect 86450 30567 86451 30568
rect 85850 30566 85851 30567
rect 86451 30566 86452 30567
rect 85850 29967 85851 29968
rect 86451 29967 86452 29968
rect 85851 29966 85852 29967
rect 86450 29966 86451 29967
rect 86463 29955 86497 30579
rect 86577 29955 86611 30579
rect 88094 29955 91736 30693
rect 104936 30668 104940 30673
rect 104866 30640 104912 30645
rect 104866 30633 104934 30640
rect 104872 30630 104934 30633
rect 83432 29893 83513 29940
rect 83572 29921 91736 29955
rect 83818 29909 83819 29910
rect 83819 29908 83820 29909
rect 83479 29325 83513 29893
rect 83819 29309 83820 29310
rect 83818 29308 83819 29309
rect 83831 29297 83865 29921
rect 83877 29909 83878 29910
rect 84476 29909 84477 29910
rect 83876 29908 83877 29909
rect 84477 29908 84478 29909
rect 84489 29312 84523 29921
rect 84535 29909 84536 29910
rect 85134 29909 85135 29910
rect 84534 29908 84535 29909
rect 85135 29908 85136 29909
rect 84714 29312 84926 29444
rect 83876 29309 83877 29310
rect 83877 29308 83878 29309
rect 84404 29297 84926 29312
rect 85135 29309 85136 29310
rect 85134 29308 85135 29309
rect 85147 29297 85181 29921
rect 85193 29909 85194 29910
rect 85792 29909 85793 29910
rect 85192 29908 85193 29909
rect 85793 29908 85794 29909
rect 85192 29309 85193 29310
rect 85793 29309 85794 29310
rect 85193 29308 85194 29309
rect 85792 29308 85793 29309
rect 85805 29297 85839 29921
rect 85851 29909 85852 29910
rect 86450 29909 86451 29910
rect 85850 29908 85851 29909
rect 86451 29908 86452 29909
rect 85850 29309 85851 29310
rect 86451 29309 86452 29310
rect 85851 29308 85852 29309
rect 86450 29308 86451 29309
rect 86463 29297 86497 29921
rect 86577 29297 86611 29921
rect 87288 29878 87678 29912
rect 86642 29396 86898 29402
rect 87288 29380 87322 29878
rect 87502 29810 87549 29857
rect 87464 29776 87549 29810
rect 87391 29717 87436 29728
rect 87519 29717 87564 29728
rect 87402 29541 87436 29717
rect 87530 29541 87564 29717
rect 87502 29482 87549 29529
rect 87464 29448 87549 29482
rect 87644 29380 87678 29878
rect 87798 29396 88054 29414
rect 86670 29368 86870 29374
rect 87288 29346 87678 29380
rect 87826 29368 88026 29386
rect 83432 29235 83513 29282
rect 83572 29263 86611 29297
rect 83818 29251 83819 29252
rect 83819 29250 83820 29251
rect 83479 28667 83513 29235
rect 83819 28651 83820 28652
rect 83818 28650 83819 28651
rect 83831 28639 83865 29263
rect 83877 29251 83878 29252
rect 83876 29250 83877 29251
rect 84404 29242 84926 29263
rect 85134 29251 85135 29252
rect 85135 29250 85136 29251
rect 83871 29214 83948 29230
rect 84396 29214 84483 29230
rect 83876 28651 83877 28652
rect 84477 28651 84478 28652
rect 83877 28650 83878 28651
rect 84476 28650 84477 28651
rect 84489 28639 84523 29242
rect 84529 29214 84610 29230
rect 84714 28996 84926 29242
rect 85058 29214 85141 29230
rect 84534 28651 84535 28652
rect 85135 28651 85136 28652
rect 84535 28650 84536 28651
rect 85134 28650 85135 28651
rect 85147 28639 85181 29263
rect 85193 29251 85194 29252
rect 85792 29251 85793 29252
rect 85192 29250 85193 29251
rect 85793 29250 85794 29251
rect 85187 29214 85212 29230
rect 85192 28651 85193 28652
rect 85793 28651 85794 28652
rect 85193 28650 85194 28651
rect 85792 28650 85793 28651
rect 85805 28639 85839 29263
rect 85851 29251 85852 29252
rect 86450 29251 86451 29252
rect 85850 29250 85851 29251
rect 86451 29250 86452 29251
rect 85850 28651 85851 28652
rect 86451 28651 86452 28652
rect 85851 28650 85852 28651
rect 86450 28650 86451 28651
rect 86463 28639 86497 29263
rect 86577 28639 86611 29263
rect 86870 29182 87130 29202
rect 86870 29154 87130 29174
rect 87274 28676 87696 29296
rect 87826 29186 88026 29202
rect 87798 29158 88054 29174
rect 88094 28639 91736 29921
rect 102714 29219 103150 29242
rect 102748 29185 103116 29208
rect 103621 29120 103655 30587
rect 104880 30448 104934 30630
rect 104880 30160 104912 30448
rect 104872 30157 104912 30160
rect 104866 30145 104912 30157
rect 104936 30420 104962 30668
rect 106182 30642 106228 30645
rect 106164 30633 106228 30642
rect 112610 30644 112614 30649
rect 106164 30630 106222 30633
rect 106164 30456 106180 30630
rect 112610 30458 112638 30644
rect 104936 30117 104940 30420
rect 106182 30157 106222 30160
rect 106182 30145 106228 30157
rect 104934 30064 105502 30098
rect 107706 29798 107930 29818
rect 109898 29802 110118 29822
rect 107726 29646 107727 29798
rect 107910 29646 107930 29798
rect 109918 29646 109919 29802
rect 110098 29646 110118 29802
rect 112610 29606 112614 30458
rect 103078 29086 105218 29120
rect 96888 28682 96944 28684
rect 83432 28577 83513 28624
rect 83572 28605 91736 28639
rect 83818 28593 83819 28594
rect 83819 28592 83820 28593
rect 83479 28009 83513 28577
rect 83819 27993 83820 27994
rect 83818 27992 83819 27993
rect 83831 27981 83865 28605
rect 83877 28593 83878 28594
rect 84476 28593 84477 28594
rect 83876 28592 83877 28593
rect 84477 28592 84478 28593
rect 83876 27993 83877 27994
rect 84477 27993 84478 27994
rect 83877 27992 83878 27993
rect 84476 27992 84477 27993
rect 84489 27981 84523 28605
rect 84535 28593 84536 28594
rect 85134 28593 85135 28594
rect 84534 28592 84535 28593
rect 85135 28592 85136 28593
rect 84534 27993 84535 27994
rect 85135 27993 85136 27994
rect 84535 27992 84536 27993
rect 85134 27992 85135 27993
rect 85147 27981 85181 28605
rect 85193 28593 85194 28594
rect 85792 28593 85793 28594
rect 85192 28592 85193 28593
rect 85793 28592 85794 28593
rect 85192 27993 85193 27994
rect 85793 27993 85794 27994
rect 85193 27992 85194 27993
rect 85792 27992 85793 27993
rect 85805 27981 85839 28605
rect 85851 28593 85852 28594
rect 86450 28593 86451 28594
rect 85850 28592 85851 28593
rect 86451 28592 86452 28593
rect 85850 27993 85851 27994
rect 86451 27993 86452 27994
rect 85851 27992 85852 27993
rect 86450 27992 86451 27993
rect 86463 27981 86497 28605
rect 86577 27981 86611 28605
rect 87838 28534 87880 28540
rect 88018 28534 88046 28540
rect 87810 28506 87880 28512
rect 88018 28506 88074 28512
rect 88094 27981 91736 28605
rect 103078 28595 103112 29086
rect 103519 29018 103553 29086
rect 103621 29018 103655 29086
rect 103254 28984 103655 29018
rect 103471 28937 103472 28938
rect 103472 28936 103473 28937
rect 103181 28925 103226 28936
rect 103192 28595 103226 28925
rect 103519 28623 103553 28984
rect 103237 28607 103238 28608
rect 103238 28606 103239 28607
rect 103460 28595 103471 28606
rect 103044 28561 103471 28595
rect 96888 28520 96944 28524
rect 96888 28464 96944 28468
rect 83432 27919 83513 27966
rect 83572 27947 91736 27981
rect 83818 27935 83819 27936
rect 83819 27934 83820 27935
rect 83479 27351 83513 27919
rect 83819 27335 83820 27336
rect 83818 27334 83819 27335
rect 83831 27323 83865 27947
rect 83877 27935 83878 27936
rect 84476 27935 84477 27936
rect 83876 27934 83877 27935
rect 84477 27934 84478 27935
rect 83876 27335 83877 27336
rect 84477 27335 84478 27336
rect 83877 27334 83878 27335
rect 84476 27334 84477 27335
rect 84489 27323 84523 27947
rect 84535 27935 84536 27936
rect 85134 27935 85135 27936
rect 84534 27934 84535 27935
rect 85135 27934 85136 27935
rect 84534 27335 84535 27336
rect 85135 27335 85136 27336
rect 84535 27334 84536 27335
rect 85134 27334 85135 27335
rect 85147 27323 85181 27947
rect 85193 27935 85194 27936
rect 85792 27935 85793 27936
rect 85192 27934 85193 27935
rect 85793 27934 85794 27935
rect 85192 27335 85193 27336
rect 85793 27335 85794 27336
rect 85193 27334 85194 27335
rect 85792 27334 85793 27335
rect 85805 27323 85839 27947
rect 85851 27935 85852 27936
rect 86450 27935 86451 27936
rect 85850 27934 85851 27935
rect 86451 27934 86452 27935
rect 85850 27335 85851 27336
rect 86451 27335 86452 27336
rect 85851 27334 85852 27335
rect 86450 27334 86451 27335
rect 86463 27323 86497 27947
rect 86577 27323 86611 27947
rect 87276 27941 87532 27947
rect 87304 27913 87504 27932
rect 83572 27289 86611 27323
rect 83831 27209 83865 27289
rect 84489 27209 84523 27289
rect 85147 27209 85181 27289
rect 85805 27209 85839 27289
rect 86463 27209 86497 27289
rect 86577 27209 86611 27289
rect 88094 27209 91736 27947
rect 103078 27937 103112 28561
rect 103192 27949 103226 28561
rect 103238 28549 103239 28550
rect 103237 28548 103238 28549
rect 103472 28533 103553 28580
rect 103237 27949 103238 27950
rect 103238 27948 103239 27949
rect 103256 27948 103258 27971
rect 103519 27965 103553 28533
rect 103256 27937 103286 27943
rect 103460 27937 103471 27948
rect 103044 27903 103146 27937
rect 103154 27924 103472 27937
rect 103154 27911 103476 27924
rect 103204 27903 103476 27911
rect 103078 27788 103112 27903
rect 103214 27897 103472 27903
rect 103238 27891 103472 27897
rect 103242 27890 103294 27891
rect 103621 27890 103655 28984
rect 106396 28728 106420 28938
rect 104550 28212 104574 28220
rect 104550 27960 104576 28212
rect 104550 27948 104574 27960
rect 103238 27869 103655 27890
rect 103254 27856 103655 27869
rect 103519 27788 103553 27856
rect 103621 27788 103655 27856
rect 83377 27175 91718 27209
rect 86577 26860 86611 27175
rect 88094 27139 91718 27175
rect 83336 26824 86647 26860
rect 88130 26824 88164 27139
rect 90248 26874 90252 27036
rect 90286 26912 90290 26998
rect 83336 26790 91580 26824
rect 91648 26790 91658 26858
rect 83234 26510 83248 26648
rect 83336 26510 86647 26790
rect 88130 26710 88164 26790
rect 88244 26710 88278 26790
rect 88290 26710 88890 26721
rect 88902 26710 88936 26790
rect 88948 26710 89548 26721
rect 89560 26710 89594 26790
rect 89606 26710 90206 26721
rect 90218 26710 90252 26790
rect 90264 26710 90864 26721
rect 90876 26710 90910 26790
rect 90922 26710 91522 26721
rect 91534 26710 91568 26790
rect 91652 26728 91682 26762
rect 88096 26688 91568 26710
rect 88096 26686 91574 26688
rect 88096 26676 91580 26686
rect 83158 26474 86647 26510
rect 83158 26440 86746 26474
rect 83158 26052 86647 26440
rect 86712 26052 86746 26440
rect 87416 26306 87864 26468
rect 87340 26256 87864 26306
rect 87340 26152 87494 26256
rect 88130 26052 88164 26676
rect 88244 26664 88278 26676
rect 88290 26664 88291 26665
rect 88889 26664 88890 26665
rect 88902 26664 88936 26676
rect 88948 26664 88949 26665
rect 89547 26664 89548 26665
rect 89560 26664 89594 26676
rect 89606 26664 89607 26665
rect 90205 26664 90206 26665
rect 90218 26664 90252 26676
rect 90264 26664 90265 26665
rect 90863 26664 90864 26665
rect 90876 26664 90910 26676
rect 90922 26664 90923 26665
rect 91521 26664 91522 26665
rect 88244 26663 88290 26664
rect 88890 26663 88891 26664
rect 88902 26663 88948 26664
rect 89548 26663 89549 26664
rect 89560 26663 89606 26664
rect 90206 26663 90207 26664
rect 90218 26663 90264 26664
rect 90864 26663 90865 26664
rect 90876 26663 90922 26664
rect 91522 26663 91523 26664
rect 88244 26505 88289 26663
rect 88902 26505 88947 26663
rect 89560 26505 89605 26663
rect 90218 26505 90263 26663
rect 90876 26505 90921 26663
rect 91534 26660 91580 26676
rect 91534 26648 91602 26660
rect 91534 26592 91606 26648
rect 91534 26505 91580 26592
rect 91584 26505 91606 26592
rect 91648 26505 91665 26695
rect 91686 26505 91720 26790
rect 88235 26052 91756 26505
rect 91812 26472 91859 26505
rect 83158 26018 86746 26052
rect 88096 26018 91756 26052
rect 83158 25394 86647 26018
rect 86712 25394 86746 26018
rect 88130 25394 88164 26018
rect 88235 25394 91756 26018
rect 83158 25360 86746 25394
rect 88096 25360 91756 25394
rect 80211 23815 80245 25058
rect 80869 23815 80903 25058
rect 78225 23781 81573 23815
rect 78237 18286 78271 23781
rect 78895 23760 78929 23781
rect 79553 23760 79587 23781
rect 80211 23760 80245 23781
rect 80869 23760 80903 23781
rect 81527 23760 81561 23781
rect 78867 23713 78929 23760
rect 79525 23713 79587 23760
rect 80183 23713 80245 23760
rect 80841 23713 80903 23760
rect 81499 23713 81561 23760
rect 78283 23679 78929 23713
rect 78941 23679 79587 23713
rect 79599 23679 80245 23713
rect 80257 23679 80903 23713
rect 80915 23679 81561 23713
rect 78895 19468 78929 23679
rect 78410 19434 78800 19468
rect 78410 18936 78444 19434
rect 78624 19366 78671 19413
rect 78586 19332 78671 19366
rect 78513 19273 78558 19284
rect 78641 19273 78686 19284
rect 78524 19097 78558 19273
rect 78652 19097 78686 19273
rect 78624 19038 78671 19085
rect 78586 19004 78671 19038
rect 78766 18936 78800 19434
rect 78410 18902 78800 18936
rect 78886 19434 79276 19468
rect 78886 18936 78929 19434
rect 79100 19366 79147 19413
rect 79062 19332 79147 19366
rect 78989 19273 79034 19284
rect 79117 19273 79162 19284
rect 79000 19097 79034 19273
rect 79128 19097 79162 19273
rect 79100 19038 79147 19085
rect 79062 19004 79147 19038
rect 79242 18936 79276 19434
rect 78886 18902 79276 18936
rect 78895 18852 78929 18902
rect 78392 18286 78814 18852
rect 78868 18286 79290 18852
rect 79553 18286 79587 23679
rect 80211 18286 80245 23679
rect 80776 18532 80792 20046
rect 80869 18286 80903 23679
rect 81527 18286 81561 23679
rect 78237 18239 79290 18286
rect 79525 18273 79587 18286
rect 80183 18273 80245 18286
rect 79525 18245 79593 18273
rect 80183 18245 80251 18273
rect 80841 18245 80903 18286
rect 79519 18239 79593 18245
rect 79603 18239 79621 18245
rect 80177 18239 80251 18245
rect 80261 18239 80279 18245
rect 80807 18239 80903 18245
rect 81499 18239 81561 18286
rect 78237 18171 78277 18239
rect 78287 18232 79593 18239
rect 78287 18205 78935 18232
rect 78287 18199 78305 18205
rect 78861 18199 78879 18205
rect 78889 18171 78935 18205
rect 78945 18205 79593 18232
rect 79599 18205 80251 18239
rect 80257 18205 80903 18239
rect 80915 18205 81561 18239
rect 81562 18220 81595 21898
rect 78945 18199 78963 18205
rect 79519 18199 79537 18205
rect 79547 18171 79593 18205
rect 79603 18199 79621 18205
rect 80177 18199 80195 18205
rect 80205 18171 80251 18205
rect 80261 18199 80279 18205
rect 80807 18199 80853 18205
rect 80863 18171 80903 18205
rect 78237 18137 78271 18171
rect 78895 18137 78929 18171
rect 79553 18137 79587 18171
rect 80211 18137 80245 18171
rect 80869 18137 80903 18171
rect 81527 18137 81561 18205
rect 78219 18103 81573 18137
rect 81579 18103 81595 18137
rect 78410 16780 78800 16814
rect 78410 16282 78444 16780
rect 78624 16712 78671 16759
rect 78586 16678 78671 16712
rect 78513 16619 78558 16630
rect 78641 16619 78686 16630
rect 78524 16443 78558 16619
rect 78652 16443 78686 16619
rect 78624 16384 78671 16431
rect 78586 16350 78671 16384
rect 78766 16282 78800 16780
rect 78410 16248 78800 16282
rect 78886 16780 79276 16814
rect 78886 16752 78920 16780
rect 78886 16344 78954 16752
rect 79100 16712 79147 16759
rect 79062 16678 79147 16712
rect 78989 16619 79034 16630
rect 79117 16619 79162 16630
rect 79000 16443 79034 16619
rect 79128 16443 79162 16619
rect 79100 16384 79147 16431
rect 79062 16350 79147 16384
rect 78886 16282 78920 16344
rect 79242 16282 79276 16780
rect 79512 16430 79516 16570
rect 78886 16248 79276 16282
rect 78392 15585 78814 16198
rect 78299 15551 78867 15585
rect 78868 15578 79290 16198
rect 80896 15934 80940 16570
rect 80896 15647 80909 15934
rect 80952 15906 80968 16570
rect 80869 15644 80909 15647
rect 80863 15632 80909 15644
rect 81641 15545 81675 25058
rect 83158 25035 86647 25360
rect 83194 18198 83228 25035
rect 83338 23820 83342 25035
rect 83372 23820 83406 25035
rect 83474 24764 83508 25035
rect 83954 24748 83955 24749
rect 83953 24747 83954 24748
rect 83966 24736 84000 25035
rect 84011 24748 84012 24749
rect 84612 24748 84613 24749
rect 84012 24747 84013 24748
rect 84611 24747 84612 24748
rect 84624 24736 84658 25035
rect 84669 24748 84670 24749
rect 85270 24748 85271 24749
rect 84670 24747 84671 24748
rect 85269 24747 85270 24748
rect 85282 24736 85316 25035
rect 85327 24748 85328 24749
rect 85928 24748 85929 24749
rect 85328 24747 85329 24748
rect 85927 24747 85928 24748
rect 85940 24736 85974 25035
rect 85985 24748 85986 24749
rect 86586 24748 86587 24749
rect 85986 24747 85987 24748
rect 86585 24747 86586 24748
rect 86598 24736 86632 25035
rect 86712 24736 86746 25360
rect 88130 25128 88164 25360
rect 88235 25128 91756 25360
rect 88130 25094 91756 25128
rect 83436 24674 83508 24712
rect 83558 24702 86746 24736
rect 83953 24690 83954 24691
rect 83954 24689 83955 24690
rect 83474 24106 83508 24674
rect 83954 24090 83955 24091
rect 83953 24089 83954 24090
rect 83966 24078 84000 24702
rect 84012 24690 84013 24691
rect 84611 24690 84612 24691
rect 84011 24689 84012 24690
rect 84612 24689 84613 24690
rect 84011 24090 84012 24091
rect 84612 24090 84613 24091
rect 84012 24089 84013 24090
rect 84611 24089 84612 24090
rect 84624 24078 84658 24702
rect 84670 24690 84671 24691
rect 85269 24690 85270 24691
rect 84669 24689 84670 24690
rect 85270 24689 85271 24690
rect 84669 24090 84670 24091
rect 85270 24090 85271 24091
rect 84670 24089 84671 24090
rect 85269 24089 85270 24090
rect 85282 24078 85316 24702
rect 85328 24690 85329 24691
rect 85927 24690 85928 24691
rect 85327 24689 85328 24690
rect 85928 24689 85929 24690
rect 85327 24090 85328 24091
rect 85928 24090 85929 24091
rect 85328 24089 85329 24090
rect 85927 24089 85928 24090
rect 85940 24078 85974 24702
rect 85986 24690 85987 24691
rect 86585 24690 86586 24691
rect 85985 24689 85986 24690
rect 86586 24689 86587 24690
rect 85985 24090 85986 24091
rect 86586 24090 86587 24091
rect 85986 24089 85987 24090
rect 86585 24089 86586 24090
rect 86598 24078 86632 24702
rect 86712 24078 86746 24702
rect 83436 24016 83508 24054
rect 83558 24044 86746 24078
rect 83953 24032 83954 24033
rect 83954 24031 83955 24032
rect 83474 23820 83508 24016
rect 83966 23820 84000 24044
rect 84012 24032 84013 24033
rect 84611 24032 84612 24033
rect 84011 24031 84012 24032
rect 84612 24031 84613 24032
rect 84624 23820 84658 24044
rect 84670 24032 84671 24033
rect 85269 24032 85270 24033
rect 84669 24031 84670 24032
rect 85270 24031 85271 24032
rect 85282 23820 85316 24044
rect 85328 24032 85329 24033
rect 85927 24032 85928 24033
rect 85327 24031 85328 24032
rect 85928 24031 85929 24032
rect 85940 23820 85974 24044
rect 85986 24032 85987 24033
rect 86585 24032 86586 24033
rect 85985 24031 85986 24032
rect 86586 24031 86587 24032
rect 86598 23820 86632 24044
rect 86712 23820 86746 24044
rect 83296 23786 86746 23820
rect 83308 21789 83342 23786
rect 83372 23756 83406 23786
rect 83372 23718 83410 23756
rect 83474 23718 83508 23786
rect 83966 23756 84000 23786
rect 84624 23756 84658 23786
rect 85282 23756 85316 23786
rect 85940 23756 85974 23786
rect 86598 23756 86632 23786
rect 83938 23718 84000 23756
rect 84596 23718 84658 23756
rect 85254 23718 85316 23756
rect 85912 23718 85974 23756
rect 86570 23718 86632 23756
rect 83354 23684 84000 23718
rect 84012 23684 84658 23718
rect 84670 23684 85316 23718
rect 85328 23684 85974 23718
rect 85986 23684 86632 23718
rect 83372 23306 83406 23684
rect 83474 23448 83508 23684
rect 83954 23432 83955 23433
rect 83953 23431 83954 23432
rect 83966 23420 84000 23684
rect 84011 23432 84012 23433
rect 84612 23432 84613 23433
rect 84012 23431 84013 23432
rect 84611 23431 84612 23432
rect 84624 23420 84658 23684
rect 84669 23432 84670 23433
rect 85270 23432 85271 23433
rect 84670 23431 84671 23432
rect 85269 23431 85270 23432
rect 85282 23420 85316 23684
rect 85327 23432 85328 23433
rect 85928 23432 85929 23433
rect 85328 23431 85329 23432
rect 85927 23431 85928 23432
rect 85940 23420 85974 23684
rect 85985 23432 85986 23433
rect 86586 23432 86587 23433
rect 85986 23431 85987 23432
rect 86585 23431 86586 23432
rect 86598 23420 86632 23684
rect 86712 23420 86746 23786
rect 83558 23386 86746 23420
rect 83966 23306 84000 23386
rect 84624 23306 84658 23386
rect 85282 23306 85316 23386
rect 85940 23306 85974 23386
rect 86598 23306 86632 23386
rect 86712 23306 86746 23386
rect 88235 23306 91756 25094
rect 83372 23272 91756 23306
rect 86684 22990 86686 23020
rect 86712 21789 86746 23272
rect 88235 23236 91756 23272
rect 83308 21753 86782 21789
rect 88271 21753 88305 23236
rect 89026 22620 89077 22804
rect 88922 22502 89077 22620
rect 89026 22348 89077 22502
rect 91675 21753 91681 21787
rect 83308 21719 91721 21753
rect 83308 18342 86782 21719
rect 88271 21639 88305 21719
rect 88385 21639 88419 21719
rect 89043 21639 89077 21719
rect 89701 21639 89735 21719
rect 90359 21639 90393 21719
rect 91017 21639 91051 21719
rect 91709 21691 91721 21719
rect 91675 21657 91721 21691
rect 91548 21639 91559 21650
rect 88271 21605 91559 21639
rect 88271 20981 88305 21605
rect 88385 20981 88419 21605
rect 88431 21593 88432 21594
rect 89030 21593 89031 21594
rect 88430 21592 88431 21593
rect 89031 21592 89032 21593
rect 88430 20993 88431 20994
rect 89031 20993 89032 20994
rect 88431 20992 88432 20993
rect 89030 20992 89031 20993
rect 89043 20981 89077 21605
rect 89089 21593 89090 21594
rect 89688 21593 89689 21594
rect 89088 21592 89089 21593
rect 89689 21592 89690 21593
rect 89088 20993 89089 20994
rect 89689 20993 89690 20994
rect 89089 20992 89090 20993
rect 89688 20992 89689 20993
rect 89701 20981 89735 21605
rect 89747 21593 89748 21594
rect 90346 21593 90347 21594
rect 89746 21592 89747 21593
rect 90347 21592 90348 21593
rect 89746 20993 89747 20994
rect 90347 20993 90348 20994
rect 89747 20992 89748 20993
rect 90346 20992 90347 20993
rect 90359 20981 90393 21605
rect 90405 21593 90406 21594
rect 91004 21593 91005 21594
rect 90404 21592 90405 21593
rect 91005 21592 91006 21593
rect 90404 20993 90405 20994
rect 91005 20993 91006 20994
rect 90405 20992 90406 20993
rect 91004 20992 91005 20993
rect 91017 20981 91051 21605
rect 91063 21593 91064 21594
rect 91062 21592 91063 21593
rect 91560 21589 91641 21624
rect 91669 21615 91675 21617
rect 91560 21577 91647 21589
rect 91573 21522 91592 21577
rect 91601 21522 91647 21577
rect 91669 21550 91679 21615
rect 91607 21074 91654 21522
rect 91062 20993 91063 20994
rect 91063 20992 91064 20993
rect 91548 20981 91559 20992
rect 88271 20947 91559 20981
rect 91573 20969 91592 21074
rect 91601 21009 91647 21074
rect 91601 20997 91620 21009
rect 91641 20997 91647 21009
rect 91669 21046 91682 21550
rect 91669 20971 91679 21046
rect 91669 20969 91675 20971
rect 88271 20323 88305 20947
rect 88385 20323 88419 20947
rect 88431 20935 88432 20936
rect 89030 20935 89031 20936
rect 88430 20934 88431 20935
rect 89031 20934 89032 20935
rect 88430 20335 88431 20336
rect 89031 20335 89032 20336
rect 88431 20334 88432 20335
rect 89030 20334 89031 20335
rect 89043 20323 89077 20947
rect 89089 20935 89090 20936
rect 89688 20935 89689 20936
rect 89088 20934 89089 20935
rect 89689 20934 89690 20935
rect 89088 20335 89089 20336
rect 89689 20335 89690 20336
rect 89089 20334 89090 20335
rect 89688 20334 89689 20335
rect 89701 20323 89735 20947
rect 89747 20935 89748 20936
rect 90346 20935 90347 20936
rect 89746 20934 89747 20935
rect 90347 20934 90348 20935
rect 89746 20335 89747 20336
rect 90347 20335 90348 20336
rect 89747 20334 89748 20335
rect 90346 20334 90347 20335
rect 90359 20323 90393 20947
rect 90405 20935 90406 20936
rect 91004 20935 91005 20936
rect 90404 20934 90405 20935
rect 91005 20934 91006 20935
rect 90404 20335 90405 20336
rect 91005 20335 91006 20336
rect 90405 20334 90406 20335
rect 91004 20334 91005 20335
rect 91017 20323 91051 20947
rect 91063 20935 91064 20936
rect 91062 20934 91063 20935
rect 91560 20931 91641 20966
rect 91669 20957 91675 20959
rect 91560 20919 91647 20931
rect 91573 20870 91592 20919
rect 91601 20870 91647 20919
rect 91669 20898 91679 20957
rect 91607 20422 91654 20870
rect 91062 20335 91063 20336
rect 91063 20334 91064 20335
rect 91548 20323 91559 20334
rect 88271 20289 91559 20323
rect 91573 20311 91592 20422
rect 91601 20351 91647 20422
rect 91601 20339 91620 20351
rect 91641 20339 91647 20351
rect 91669 20394 91682 20898
rect 91669 20313 91679 20394
rect 91669 20311 91675 20313
rect 88271 19665 88305 20289
rect 88385 19665 88419 20289
rect 88431 20277 88432 20278
rect 89030 20277 89031 20278
rect 88430 20276 88431 20277
rect 89031 20276 89032 20277
rect 88430 19677 88431 19678
rect 89031 19677 89032 19678
rect 88431 19676 88432 19677
rect 89030 19676 89031 19677
rect 89043 19665 89077 20289
rect 89089 20277 89090 20278
rect 89688 20277 89689 20278
rect 89088 20276 89089 20277
rect 89689 20276 89690 20277
rect 89088 19677 89089 19678
rect 89689 19677 89690 19678
rect 89089 19676 89090 19677
rect 89688 19676 89689 19677
rect 89701 19665 89735 20289
rect 89747 20277 89748 20278
rect 90346 20277 90347 20278
rect 89746 20276 89747 20277
rect 90347 20276 90348 20277
rect 90359 19684 90393 20289
rect 90405 20277 90406 20278
rect 91004 20277 91005 20278
rect 90404 20276 90405 20277
rect 91005 20276 91006 20277
rect 90622 19684 90834 19814
rect 89746 19677 89747 19678
rect 89747 19676 89748 19677
rect 90178 19665 90834 19684
rect 91005 19677 91006 19678
rect 91004 19676 91005 19677
rect 91017 19665 91051 20289
rect 91063 20277 91064 20278
rect 91062 20276 91063 20277
rect 91560 20273 91641 20308
rect 91669 20299 91675 20301
rect 91560 20261 91647 20273
rect 91573 20200 91592 20261
rect 91601 20200 91647 20261
rect 91669 20228 91679 20299
rect 91607 19752 91654 20200
rect 91669 20160 91682 20228
rect 91709 20160 91721 21657
rect 91062 19677 91063 19678
rect 91063 19676 91064 19677
rect 91548 19665 91559 19676
rect 88271 19631 91559 19665
rect 91573 19653 91592 19752
rect 91601 19693 91647 19752
rect 91601 19681 91620 19693
rect 91641 19681 91647 19693
rect 91669 19653 91721 20160
rect 87166 19434 87556 19468
rect 86790 18967 87046 18970
rect 86818 18939 87018 18942
rect 87166 18936 87200 19434
rect 87380 19366 87427 19413
rect 87342 19332 87427 19366
rect 87269 19273 87314 19284
rect 87397 19273 87442 19284
rect 87280 19097 87314 19273
rect 87408 19097 87442 19273
rect 87380 19041 87427 19085
rect 87342 19019 87427 19041
rect 87326 19007 87427 19019
rect 87326 18988 87396 19007
rect 87522 18970 87556 19434
rect 87266 18967 87556 18970
rect 87300 18950 87420 18967
rect 87294 18939 87494 18942
rect 87294 18936 87448 18939
rect 87522 18936 87556 18967
rect 87166 18902 87556 18936
rect 87642 19434 88032 19468
rect 87642 18936 87676 19434
rect 87856 19366 87903 19413
rect 87818 19332 87903 19366
rect 87745 19273 87790 19284
rect 87873 19273 87918 19284
rect 87756 19097 87790 19273
rect 87884 19097 87918 19273
rect 87856 19041 87903 19085
rect 87818 19019 87903 19041
rect 87802 19007 87903 19019
rect 87802 18988 87872 19007
rect 87776 18950 87896 18952
rect 87998 18936 88032 19434
rect 87642 18902 88032 18936
rect 88271 19007 88305 19631
rect 88385 19007 88419 19631
rect 88431 19619 88432 19620
rect 89030 19619 89031 19620
rect 88430 19618 88431 19619
rect 89031 19618 89032 19619
rect 88430 19019 88431 19020
rect 89031 19019 89032 19020
rect 88431 19018 88432 19019
rect 89030 19018 89031 19019
rect 89043 19007 89077 19631
rect 89089 19619 89090 19620
rect 89688 19619 89689 19620
rect 89088 19618 89089 19619
rect 89689 19618 89690 19619
rect 89088 19019 89089 19020
rect 89689 19019 89690 19020
rect 89089 19018 89090 19019
rect 89688 19018 89689 19019
rect 89701 19007 89735 19631
rect 89747 19619 89748 19620
rect 89746 19618 89747 19619
rect 90178 19610 90834 19631
rect 91004 19619 91005 19620
rect 91005 19618 91006 19619
rect 89746 19019 89747 19020
rect 90347 19019 90348 19020
rect 89747 19018 89748 19019
rect 90346 19018 90347 19019
rect 90359 19007 90393 19610
rect 90622 19366 90834 19610
rect 90404 19019 90405 19020
rect 91005 19019 91006 19020
rect 90405 19018 90406 19019
rect 91004 19018 91005 19019
rect 91017 19007 91051 19631
rect 91063 19619 91064 19620
rect 91062 19618 91063 19619
rect 91560 19615 91641 19650
rect 91675 19643 91721 19653
rect 91560 19603 91647 19615
rect 91573 19538 91592 19603
rect 91601 19538 91647 19603
rect 91669 19538 91721 19643
rect 91607 19090 91641 19538
rect 91675 19090 91721 19538
rect 91062 19019 91063 19020
rect 91063 19018 91064 19019
rect 91548 19007 91559 19018
rect 88271 18973 91559 19007
rect 91573 18995 91592 19090
rect 91601 19035 91647 19090
rect 91601 19023 91620 19035
rect 91641 19023 91647 19035
rect 91669 18995 91721 19090
rect 87148 18746 87570 18852
rect 87624 18746 88046 18852
rect 87148 18534 88046 18746
rect 87148 18342 87570 18534
rect 87624 18342 88046 18534
rect 88271 18349 88305 18973
rect 88385 18349 88419 18973
rect 88431 18961 88432 18962
rect 89030 18961 89031 18962
rect 88430 18960 88431 18961
rect 89031 18960 89032 18961
rect 88430 18361 88431 18362
rect 89031 18361 89032 18362
rect 88431 18360 88432 18361
rect 89030 18360 89031 18361
rect 89043 18349 89077 18973
rect 89089 18961 89090 18962
rect 89688 18961 89689 18962
rect 89088 18960 89089 18961
rect 89689 18960 89690 18961
rect 89088 18361 89089 18362
rect 89689 18361 89690 18362
rect 89089 18360 89090 18361
rect 89688 18360 89689 18361
rect 89701 18349 89735 18973
rect 89747 18961 89748 18962
rect 90346 18961 90347 18962
rect 89746 18960 89747 18961
rect 90347 18960 90348 18961
rect 89746 18361 89747 18362
rect 90347 18361 90348 18362
rect 89747 18360 89748 18361
rect 90346 18360 90347 18361
rect 90359 18349 90393 18973
rect 90405 18961 90406 18962
rect 91004 18961 91005 18962
rect 90404 18960 90405 18961
rect 91005 18960 91006 18961
rect 90404 18361 90405 18362
rect 91005 18361 91006 18362
rect 90405 18360 90406 18361
rect 91004 18360 91005 18361
rect 91017 18349 91051 18973
rect 91063 18961 91064 18962
rect 91062 18960 91063 18961
rect 91560 18957 91641 18992
rect 91675 18985 91721 18995
rect 91560 18945 91647 18957
rect 91573 18880 91592 18945
rect 91601 18880 91647 18945
rect 91607 18432 91654 18880
rect 91062 18361 91063 18362
rect 91063 18360 91064 18361
rect 91548 18349 91559 18360
rect 83308 18315 88048 18342
rect 88271 18315 91559 18349
rect 91573 18337 91592 18432
rect 91601 18377 91647 18432
rect 91601 18365 91620 18377
rect 91641 18365 91647 18377
rect 91669 18337 91721 18985
rect 83308 18235 86782 18315
rect 87148 18308 87570 18315
rect 87624 18308 88046 18315
rect 86800 18281 88046 18308
rect 87148 18238 87570 18281
rect 87624 18238 88046 18281
rect 86876 18235 88046 18238
rect 88271 18235 88305 18315
rect 88385 18273 88419 18315
rect 89043 18286 89077 18315
rect 89701 18286 89735 18315
rect 90359 18286 90393 18315
rect 91017 18286 91051 18315
rect 91675 18286 91721 18337
rect 89015 18273 89077 18286
rect 89673 18273 89735 18286
rect 90331 18273 90393 18286
rect 90989 18273 91051 18286
rect 88385 18235 88425 18273
rect 89015 18245 89083 18273
rect 89673 18245 89741 18273
rect 90331 18245 90399 18273
rect 90989 18245 91057 18273
rect 91647 18245 91721 18286
rect 88435 18239 88453 18245
rect 89009 18239 89083 18245
rect 89093 18239 89111 18245
rect 89667 18239 89741 18245
rect 89751 18239 89769 18245
rect 90325 18239 90399 18245
rect 90409 18239 90427 18245
rect 90983 18239 91057 18245
rect 91067 18239 91085 18245
rect 91641 18239 91721 18245
rect 88431 18235 89083 18239
rect 89089 18235 89741 18239
rect 89747 18235 90399 18239
rect 90405 18235 91057 18239
rect 91063 18235 91721 18239
rect 83308 18201 91721 18235
rect 83308 18198 86782 18201
rect 83158 18196 86782 18198
rect 83194 18164 83228 18196
rect 83308 18165 86782 18196
rect 86876 18165 87846 18201
rect 83308 18164 83342 18165
rect 83192 18162 83448 18164
rect 83194 17339 83228 18162
rect 83308 18160 83342 18162
rect 83966 18160 84000 18165
rect 84624 18160 84658 18165
rect 85282 18160 85316 18165
rect 85940 18160 85974 18165
rect 86598 18160 86632 18165
rect 83290 18126 86666 18160
rect 83966 17339 84000 18126
rect 86748 17882 86760 18164
rect 86782 17916 86794 18138
rect 87130 17346 87592 17593
rect 83158 17303 86782 17339
rect 87148 17303 87570 17332
rect 88271 17303 88305 18201
rect 88407 18171 88425 18201
rect 88435 18199 88453 18201
rect 89009 18199 89027 18201
rect 89037 18171 89055 18201
rect 89065 18171 89083 18201
rect 89093 18199 89111 18201
rect 89667 18199 89685 18201
rect 89695 18171 89713 18201
rect 89723 18171 89741 18201
rect 89751 18199 89769 18201
rect 90325 18199 90343 18201
rect 90353 18171 90371 18201
rect 90381 18171 90399 18201
rect 90409 18199 90427 18201
rect 90983 18199 91001 18201
rect 91011 18171 91029 18201
rect 91039 18171 91057 18201
rect 91067 18199 91085 18201
rect 91641 18199 91659 18201
rect 91669 18171 91709 18201
rect 88385 18137 88419 18171
rect 89043 18137 89077 18171
rect 89701 18137 89735 18171
rect 90359 18137 90393 18171
rect 91017 18137 91051 18171
rect 91675 18137 91709 18171
rect 88367 18103 91721 18137
rect 91727 18103 91743 18137
rect 88385 17303 88419 17337
rect 89043 17303 89077 17337
rect 89701 17303 89735 17337
rect 90359 17303 90393 17337
rect 83158 17296 90851 17303
rect 82553 16519 82578 16570
rect 82581 16547 82606 16570
rect 83158 16537 86782 17296
rect 87148 17269 90851 17296
rect 86818 17222 87018 17223
rect 86790 17194 87046 17195
rect 87148 16712 87570 17269
rect 88118 17223 88174 17251
rect 87714 17218 88174 17223
rect 87974 17210 88174 17218
rect 87714 17190 88174 17195
rect 87946 17182 88174 17190
rect 88118 17154 88174 17182
rect 88271 17189 88305 17269
rect 88385 17189 88419 17269
rect 89043 17189 89077 17269
rect 89701 17189 89735 17269
rect 90359 17189 90393 17269
rect 90656 17189 90667 17200
rect 88271 17155 90667 17189
rect 87642 16780 88032 16814
rect 82668 16514 82944 16537
rect 83082 16514 86782 16537
rect 83158 16470 86782 16514
rect 87166 16531 87200 16712
rect 87342 16678 87427 16712
rect 87269 16619 87325 16630
rect 87397 16619 87453 16630
rect 87280 16570 87325 16619
rect 87408 16570 87453 16619
rect 87280 16531 87314 16570
rect 87325 16543 87326 16544
rect 87396 16543 87397 16544
rect 87326 16542 87327 16543
rect 87395 16542 87396 16543
rect 87408 16531 87442 16570
rect 87522 16531 87556 16712
rect 87166 16497 87556 16531
rect 87166 16470 87200 16497
rect 87280 16470 87314 16497
rect 87326 16485 87327 16486
rect 87395 16485 87396 16486
rect 87325 16484 87326 16485
rect 87396 16484 87397 16485
rect 87408 16470 87442 16497
rect 87522 16470 87556 16497
rect 87642 16531 87676 16780
rect 87856 16712 87903 16759
rect 87818 16678 87903 16712
rect 87998 16648 88032 16780
rect 87745 16619 87790 16630
rect 87873 16619 87918 16630
rect 87924 16624 88174 16648
rect 87998 16620 88032 16624
rect 87756 16531 87790 16619
rect 87801 16543 87802 16544
rect 87872 16543 87873 16544
rect 87802 16542 87803 16543
rect 87871 16542 87872 16543
rect 87884 16531 87918 16619
rect 87924 16596 88174 16620
rect 87998 16531 88032 16596
rect 88118 16568 88174 16596
rect 88271 16537 88305 17155
rect 87642 16497 88032 16531
rect 88190 16531 88352 16537
rect 88385 16531 88419 17155
rect 88431 17143 88432 17144
rect 89030 17143 89031 17144
rect 88430 17142 88431 17143
rect 89031 17142 89032 17143
rect 88430 16543 88431 16544
rect 89031 16543 89032 16544
rect 88431 16542 88432 16543
rect 89030 16542 89031 16543
rect 88460 16531 88502 16537
rect 88950 16531 89010 16537
rect 89043 16531 89077 17155
rect 89089 17143 89090 17144
rect 89688 17143 89689 17144
rect 89088 17142 89089 17143
rect 89689 17142 89690 17143
rect 89701 17014 89735 17155
rect 89747 17143 89748 17144
rect 90346 17143 90347 17144
rect 89746 17142 89747 17143
rect 90347 17142 90348 17143
rect 89680 16548 89754 17014
rect 89088 16543 89089 16544
rect 89089 16542 89090 16543
rect 89384 16531 89840 16548
rect 90347 16543 90348 16544
rect 90346 16542 90347 16543
rect 90359 16531 90393 17155
rect 90405 17143 90406 17144
rect 90404 17142 90405 17143
rect 90668 17127 90749 17174
rect 90715 16559 90749 17127
rect 90404 16543 90405 16544
rect 90405 16542 90406 16543
rect 90399 16531 90492 16537
rect 90656 16531 90667 16542
rect 88190 16514 90667 16531
rect 83158 16430 87616 16470
rect 83158 16414 86782 16430
rect 87166 16414 87200 16430
rect 87380 16414 87427 16430
rect 87522 16414 87556 16430
rect 83158 16374 87616 16414
rect 83158 15842 86782 16374
rect 87166 16282 87200 16374
rect 87342 16350 87427 16374
rect 87522 16282 87556 16374
rect 87166 16248 87556 16282
rect 87642 16282 87676 16497
rect 87756 16470 87790 16497
rect 87802 16485 87803 16486
rect 87871 16485 87872 16486
rect 87801 16484 87802 16485
rect 87872 16484 87873 16485
rect 87714 16431 87796 16470
rect 87884 16443 87918 16497
rect 87998 16442 88032 16497
rect 88271 16497 90667 16514
rect 87878 16440 88092 16442
rect 87878 16431 87924 16440
rect 87714 16430 87790 16431
rect 87856 16414 87903 16431
rect 87998 16414 88032 16440
rect 87714 16412 88092 16414
rect 87714 16403 87952 16412
rect 87714 16384 87852 16403
rect 87856 16384 87903 16403
rect 87714 16374 87903 16384
rect 87818 16350 87903 16374
rect 87998 16282 88032 16412
rect 87642 16248 88032 16282
rect 83158 15833 86798 15842
rect 83158 15814 86782 15833
rect 83158 15805 86798 15814
rect 74534 15472 77894 15506
rect 83158 15484 86782 15805
rect 87148 15752 87570 16198
rect 87624 15752 88046 16198
rect 87006 15734 88046 15752
rect 87148 15578 87570 15734
rect 87624 15578 88046 15734
rect 88271 15873 88305 16497
rect 88385 15873 88419 16497
rect 88431 16485 88432 16486
rect 89030 16485 89031 16486
rect 88430 16484 88431 16485
rect 89031 16484 89032 16485
rect 88954 16390 89037 16414
rect 88430 15885 88431 15886
rect 89031 15885 89032 15886
rect 88431 15884 88432 15885
rect 89030 15884 89031 15885
rect 89043 15873 89077 16497
rect 89089 16485 89090 16486
rect 89088 16484 89089 16485
rect 89384 16478 89840 16497
rect 90346 16485 90347 16486
rect 90347 16484 90348 16485
rect 89083 16390 89160 16414
rect 89608 16390 89660 16414
rect 89680 16360 89754 16478
rect 89768 16390 89822 16414
rect 90270 16390 90353 16414
rect 89088 15885 89089 15886
rect 89689 15885 89690 15886
rect 89089 15884 89090 15885
rect 89688 15884 89689 15885
rect 89701 15873 89735 16360
rect 89746 15885 89747 15886
rect 90347 15885 90348 15886
rect 89747 15884 89748 15885
rect 90346 15884 90347 15885
rect 90359 15873 90393 16497
rect 90405 16485 90406 16486
rect 90404 16484 90405 16485
rect 90668 16469 90749 16516
rect 90715 15901 90749 16469
rect 90404 15885 90405 15886
rect 90405 15884 90406 15885
rect 90656 15873 90667 15884
rect 88271 15839 90667 15873
rect 45630 14886 56014 14920
rect 45630 14850 50506 14886
rect 43952 14598 44054 14626
rect 43986 14564 44020 14592
rect 44068 14348 44468 14770
rect 44518 14718 45084 14752
rect 44518 14396 44552 14718
rect 44702 14638 44900 14649
rect 44586 14623 44688 14626
rect 44573 14598 44688 14623
rect 44713 14604 44900 14638
rect 44573 14576 44654 14598
rect 44901 14576 45029 14623
rect 44620 14538 44654 14576
rect 44948 14572 45029 14576
rect 44948 14538 44982 14572
rect 44889 14510 44900 14521
rect 44562 14474 44634 14480
rect 44713 14476 44900 14510
rect 44578 14418 44634 14424
rect 45050 14396 45084 14718
rect 44518 14362 45084 14396
rect 44104 13973 44138 14348
rect 44206 14340 44240 14348
rect 45116 14276 45750 14286
rect 50436 13973 50470 14850
rect 43715 13939 51889 13973
rect 44104 13920 44138 13939
rect 44144 13920 44200 13939
rect 44104 13916 44200 13920
rect 44104 13892 44138 13916
rect 44104 13871 44200 13892
rect 44104 13865 44287 13871
rect 43802 13860 44287 13865
rect 44104 13859 44138 13860
rect 44070 13825 44138 13859
rect 44159 13859 44287 13860
rect 50287 13859 50399 13871
rect 50436 13859 50470 13939
rect 44159 13856 50399 13859
rect 44159 13825 50384 13856
rect 50402 13825 50470 13859
rect 44104 13201 44138 13825
rect 44190 13813 44287 13825
rect 50287 13813 50384 13825
rect 44144 13784 44200 13798
rect 44144 13728 44200 13742
rect 44206 13698 44240 13813
rect 50334 13698 50368 13813
rect 50275 13670 50286 13681
rect 44159 13608 44240 13655
rect 44299 13636 50286 13670
rect 50287 13608 50368 13655
rect 44206 13214 44240 13608
rect 50334 13214 50368 13608
rect 50376 13294 50432 13300
rect 50376 13238 50430 13244
rect 44070 13167 44138 13201
rect 44159 13213 44240 13214
rect 50287 13213 50368 13214
rect 44159 13201 44287 13213
rect 50287 13201 50384 13213
rect 50436 13201 50470 13825
rect 44159 13167 50384 13201
rect 50402 13167 50470 13201
rect 44104 12898 44138 13167
rect 44190 13155 44287 13167
rect 50287 13155 50384 13167
rect 44206 13040 44240 13155
rect 50334 13040 50368 13155
rect 50436 13140 50470 13167
rect 50376 13116 51496 13140
rect 50376 13060 50432 13084
rect 50275 13012 50286 13023
rect 44299 12978 50286 13012
rect 50436 12898 50470 13116
rect 44104 12864 50470 12898
rect 44144 12580 45232 12584
rect 43814 12509 51790 12543
rect 45232 12444 45868 12450
rect 45176 12388 45924 12422
rect 54394 12156 54428 14886
rect 54434 12968 54454 14000
rect 54490 12968 54510 14056
rect 62994 12220 63028 13022
rect 63652 12220 63686 13022
rect 62544 11848 63724 12220
rect 49838 11724 51843 11752
rect 51889 11724 51902 11752
rect 32030 10772 41538 10842
rect 31970 10710 31980 10716
rect 32026 10710 41538 10772
rect 32030 10664 41538 10710
rect 19263 10470 27922 10504
rect 31348 10490 31368 10620
rect 31386 10548 31562 10600
rect 31382 10524 31864 10548
rect 31458 10486 31864 10524
rect 31970 10486 31980 10664
rect 32026 10486 41538 10664
rect 19263 10440 27232 10470
rect 27520 10440 27584 10470
rect 19263 10368 27784 10440
rect 19263 9278 27232 10368
rect 27420 10330 27478 10368
rect 27432 9278 27466 10330
rect 27520 9278 27584 10368
rect 27763 10318 27808 10329
rect 27774 9278 27808 10318
rect 27888 9278 27922 10470
rect 30288 10348 30648 10486
rect 31184 10374 41538 10486
rect 43583 10806 52021 10842
rect 56078 10806 56112 10932
rect 56192 10806 56226 10840
rect 56850 10806 56884 10840
rect 56964 10806 56998 10932
rect 57268 10806 57302 10932
rect 57382 10806 57416 10840
rect 43583 10772 58012 10806
rect 43583 10535 52021 10772
rect 43583 10385 53509 10535
rect 31184 10348 43178 10374
rect 30288 10314 43178 10348
rect 19263 9244 29092 9278
rect 19263 9176 27232 9244
rect 27432 9214 27466 9244
rect 27432 9192 27470 9214
rect 27420 9176 27478 9192
rect 27520 9176 27584 9244
rect 27774 9214 27808 9244
rect 27774 9176 27812 9214
rect 27888 9176 27922 9244
rect 28948 9214 28982 9244
rect 28190 9192 28228 9214
rect 28178 9176 28236 9192
rect 28544 9176 28982 9214
rect 19263 9142 28982 9176
rect 19263 8266 27232 9142
rect 27420 9104 27478 9142
rect 27432 8304 27466 9104
rect 27420 8266 27478 8304
rect 27520 8266 27584 9142
rect 27774 8304 27808 9142
rect 27774 8266 27812 8304
rect 27888 8266 27922 9142
rect 28178 9104 28236 9142
rect 28910 9108 28942 9132
rect 28190 8304 28224 9104
rect 28933 9092 28936 9103
rect 28938 9080 28942 9104
rect 28948 9092 28982 9142
rect 28944 8316 28982 9092
rect 28948 8304 28982 8316
rect 28178 8266 28236 8304
rect 28544 8266 28982 8304
rect 19263 8232 28982 8266
rect 19263 8164 27232 8232
rect 27420 8216 27478 8232
rect 27432 8188 27466 8216
rect 27432 8164 27477 8188
rect 27520 8164 27584 8232
rect 27774 8188 27808 8232
rect 27774 8164 27819 8188
rect 27888 8164 27922 8232
rect 28178 8216 28236 8232
rect 28914 8226 28928 8232
rect 28942 8198 28982 8232
rect 28948 8164 28982 8198
rect 29058 8164 29092 9244
rect 29916 8558 30238 8610
rect 29836 8188 30238 8558
rect 19263 8130 29092 8164
rect 19263 7820 27232 8130
rect 27432 7820 27477 8130
rect 27520 7820 27584 8130
rect 27774 7820 27819 8130
rect 27888 7820 27922 8130
rect 29916 8102 30238 8188
rect 30288 8048 30648 10314
rect 31184 8936 43178 10314
rect 31184 8668 41538 8936
rect 31184 8656 41880 8668
rect 31184 8048 32680 8656
rect 33920 8164 33954 8656
rect 34034 8316 34079 8656
rect 34366 8304 34411 8656
rect 35124 8304 35169 8656
rect 35882 8304 35927 8656
rect 36640 8304 36685 8656
rect 36994 8648 39302 8656
rect 36994 8490 39474 8648
rect 36806 8304 39474 8490
rect 34058 8266 39474 8304
rect 34096 8232 39474 8266
rect 34354 8216 34412 8232
rect 35112 8216 35170 8232
rect 35870 8216 35928 8232
rect 36628 8216 36686 8232
rect 36994 8164 39474 8232
rect 33920 8140 39474 8164
rect 33920 8130 39302 8140
rect 30578 7820 30612 8048
rect 30642 7958 30652 7966
rect 30670 7902 30708 7966
rect 31220 7820 31254 8048
rect 36994 7820 39302 8130
rect 39572 7820 41880 8656
rect 19263 7786 41880 7820
rect 19263 7726 27232 7786
rect 27432 7772 27477 7786
rect 19263 7706 22918 7726
rect 22930 7706 23306 7717
rect 23642 7706 23676 7726
rect 24370 7706 24434 7726
rect 24484 7712 24524 7726
rect 24542 7712 24552 7726
rect 24484 7706 24518 7712
rect 25142 7706 25192 7726
rect 25800 7706 25834 7726
rect 25916 7706 25950 7726
rect 26458 7706 26492 7726
rect 26534 7712 26562 7726
rect 26590 7712 26618 7726
rect 26674 7706 26708 7726
rect 27116 7706 27150 7726
rect 27432 7706 27466 7772
rect 27520 7706 27584 7786
rect 27774 7772 27819 7786
rect 27774 7766 27808 7772
rect 27888 7766 27922 7786
rect 28190 7766 28224 7786
rect 27716 7726 28352 7766
rect 27774 7710 27808 7726
rect 27888 7710 27922 7726
rect 28190 7710 28224 7726
rect 27660 7706 28352 7710
rect 28948 7706 28982 7786
rect 29706 7766 29740 7786
rect 29048 7726 30216 7766
rect 29706 7710 29740 7726
rect 29048 7706 30272 7710
rect 30300 7706 30334 7786
rect 19263 7684 30334 7706
rect 30466 7694 30500 7786
rect 30578 7706 30612 7786
rect 31220 7706 31254 7786
rect 31334 7706 31368 7786
rect 31380 7706 32080 7717
rect 32092 7706 32126 7786
rect 32138 7706 32838 7717
rect 32850 7706 32884 7786
rect 32896 7706 33498 7717
rect 33608 7706 33642 7786
rect 34366 7706 34400 7786
rect 35124 7706 35158 7786
rect 35882 7706 35916 7786
rect 36640 7706 36674 7786
rect 36700 7717 36708 7772
rect 36994 7717 39302 7786
rect 36700 7706 39494 7717
rect 39572 7706 41880 7786
rect 30464 7684 30500 7694
rect 19263 7682 30342 7684
rect 19263 7672 30436 7682
rect 19263 7660 22918 7672
rect 23574 7666 23636 7672
rect 22930 7660 22931 7661
rect 19263 7659 22930 7660
rect 19146 7512 19174 7568
rect 19263 7261 22929 7659
rect 23602 7638 23636 7664
rect 19263 7260 22930 7261
rect 23630 7260 23631 7261
rect 19263 7248 22918 7260
rect 22930 7259 22931 7260
rect 23629 7259 23630 7260
rect 22930 7248 23306 7259
rect 23642 7248 23676 7672
rect 23682 7666 23754 7672
rect 23682 7638 23726 7664
rect 23687 7260 23688 7261
rect 23688 7259 23689 7260
rect 24370 7248 24434 7672
rect 24484 7666 24518 7672
rect 25082 7666 25136 7672
rect 24446 7660 24447 7661
rect 24445 7659 24446 7660
rect 24484 7576 24524 7666
rect 24542 7576 24552 7666
rect 25110 7638 25136 7652
rect 24484 7332 24518 7576
rect 24445 7260 24446 7261
rect 24446 7259 24447 7260
rect 24484 7254 24524 7332
rect 24542 7254 24552 7332
rect 24484 7248 24518 7254
rect 25142 7248 25192 7672
rect 25198 7666 25262 7672
rect 25198 7638 25234 7652
rect 25800 7248 25834 7672
rect 25916 7248 25950 7672
rect 26458 7248 26492 7672
rect 26534 7576 26562 7666
rect 26590 7576 26618 7666
rect 26534 7254 26562 7332
rect 26590 7254 26618 7332
rect 26674 7248 26708 7672
rect 27116 7248 27150 7672
rect 27432 7248 27466 7672
rect 27660 7670 28352 7672
rect 27774 7248 27808 7670
rect 27888 7248 27922 7670
rect 28120 7666 28184 7670
rect 28148 7638 28184 7664
rect 28178 7260 28179 7261
rect 28177 7259 28178 7260
rect 28190 7248 28224 7670
rect 28230 7666 28300 7670
rect 28230 7638 28272 7664
rect 28935 7660 28936 7661
rect 28936 7659 28937 7660
rect 28235 7260 28236 7261
rect 28936 7260 28937 7261
rect 28236 7259 28237 7260
rect 28935 7259 28936 7260
rect 28948 7248 28982 7672
rect 29048 7670 30272 7672
rect 28994 7660 28995 7661
rect 29693 7660 29694 7661
rect 28993 7659 28994 7660
rect 29694 7659 29695 7660
rect 28993 7260 28994 7261
rect 29694 7260 29695 7261
rect 28994 7259 28995 7260
rect 29693 7259 29694 7260
rect 29706 7248 29740 7670
rect 29752 7660 29753 7661
rect 29751 7659 29752 7660
rect 30300 7656 30436 7672
rect 30458 7660 30500 7684
rect 30544 7672 30612 7706
rect 31186 7672 41880 7706
rect 30300 7644 30442 7656
rect 30300 7576 30342 7644
rect 30358 7576 30398 7644
rect 30300 7332 30334 7576
rect 30364 7332 30398 7576
rect 29751 7260 29752 7261
rect 29752 7259 29753 7260
rect 30300 7248 30342 7332
rect 30358 7264 30398 7332
rect 30364 7260 30398 7264
rect 30402 7576 30442 7644
rect 30402 7332 30436 7576
rect 30402 7264 30442 7332
rect 30402 7260 30436 7264
rect 30452 7260 30500 7660
rect 19263 7236 30342 7248
rect 30458 7236 30500 7260
rect 30578 7248 30612 7672
rect 31220 7248 31254 7672
rect 31268 7666 31328 7672
rect 31334 7660 31368 7672
rect 31374 7666 31448 7672
rect 31380 7660 31381 7661
rect 32079 7660 32080 7661
rect 32092 7660 32126 7672
rect 32138 7660 32139 7661
rect 32837 7660 32838 7661
rect 32850 7660 32884 7672
rect 32896 7660 32897 7661
rect 33595 7660 33596 7661
rect 31334 7659 31380 7660
rect 32080 7659 32081 7660
rect 32092 7659 32138 7660
rect 32838 7659 32839 7660
rect 32850 7659 32896 7660
rect 33596 7659 33597 7660
rect 31334 7656 31379 7659
rect 31296 7638 31328 7656
rect 31334 7638 31420 7656
rect 31334 7261 31379 7638
rect 32092 7261 32137 7659
rect 32850 7261 32895 7659
rect 31334 7260 31380 7261
rect 32080 7260 32081 7261
rect 32092 7260 32138 7261
rect 32838 7260 32839 7261
rect 32850 7260 32896 7261
rect 33596 7260 33597 7261
rect 31334 7248 31368 7260
rect 31380 7259 31381 7260
rect 32079 7259 32080 7260
rect 31380 7248 32080 7259
rect 32092 7248 32126 7260
rect 32138 7259 32139 7260
rect 32837 7259 32838 7260
rect 32138 7248 32838 7259
rect 32850 7248 32884 7260
rect 32896 7259 32897 7260
rect 33595 7259 33596 7260
rect 32896 7248 33498 7259
rect 33608 7248 33642 7672
rect 33654 7660 33655 7661
rect 34353 7660 34354 7661
rect 33653 7659 33654 7660
rect 34354 7659 34355 7660
rect 33653 7260 33654 7261
rect 34354 7260 34355 7261
rect 33654 7259 33655 7260
rect 34353 7259 34354 7260
rect 34366 7248 34400 7672
rect 34412 7660 34413 7661
rect 35111 7660 35112 7661
rect 34411 7659 34412 7660
rect 35112 7659 35113 7660
rect 34411 7260 34412 7261
rect 35112 7260 35113 7261
rect 34412 7259 34413 7260
rect 35111 7259 35112 7260
rect 35124 7248 35158 7672
rect 35810 7666 35876 7672
rect 35170 7660 35171 7661
rect 35869 7660 35870 7661
rect 35169 7659 35170 7660
rect 35870 7659 35871 7660
rect 35838 7638 35876 7648
rect 35169 7260 35170 7261
rect 35870 7260 35871 7261
rect 35170 7259 35171 7260
rect 35869 7259 35870 7260
rect 35882 7248 35916 7672
rect 35922 7666 35990 7672
rect 35928 7660 35929 7661
rect 36627 7660 36628 7661
rect 35927 7659 35928 7660
rect 36628 7659 36629 7660
rect 35922 7638 35962 7648
rect 35927 7260 35928 7261
rect 36628 7260 36629 7261
rect 35928 7259 35929 7260
rect 36627 7259 36628 7260
rect 36640 7248 36674 7672
rect 36686 7660 36687 7661
rect 36685 7659 36686 7660
rect 36685 7260 36686 7261
rect 36686 7259 36687 7260
rect 36700 7259 36708 7672
rect 36994 7259 39302 7672
rect 36700 7248 39494 7259
rect 39572 7248 41880 7672
rect 19263 7214 30334 7236
rect 30464 7226 30500 7236
rect 19263 7134 22918 7214
rect 23642 7134 23676 7214
rect 24370 7134 24434 7214
rect 24484 7208 24518 7214
rect 24484 7164 24524 7208
rect 24484 7134 24529 7164
rect 24542 7134 24552 7208
rect 25142 7164 25192 7214
rect 25800 7164 25834 7214
rect 25916 7164 25950 7214
rect 26458 7164 26492 7214
rect 25142 7134 25203 7164
rect 25800 7134 25845 7164
rect 25916 7134 25961 7164
rect 26458 7134 26503 7164
rect 26534 7134 26562 7208
rect 26590 7134 26618 7208
rect 26674 7164 26708 7214
rect 27116 7164 27150 7214
rect 27432 7164 27466 7214
rect 27774 7164 27808 7214
rect 26674 7134 26719 7164
rect 27116 7134 27161 7164
rect 27432 7134 27477 7164
rect 27774 7134 27819 7164
rect 27888 7134 27922 7214
rect 28190 7134 28224 7214
rect 28948 7134 28982 7214
rect 29706 7134 29740 7214
rect 30300 7192 30334 7214
rect 30246 7180 30334 7192
rect 30300 7134 30334 7180
rect 30466 7134 30500 7226
rect 30544 7214 30612 7248
rect 31186 7230 41880 7248
rect 31186 7214 40464 7230
rect 30578 7134 30612 7214
rect 31220 7134 31254 7214
rect 31334 7134 31368 7214
rect 32092 7134 32126 7214
rect 32850 7134 32884 7214
rect 33608 7134 33642 7214
rect 34366 7134 34400 7214
rect 35124 7134 35158 7214
rect 35882 7134 35916 7214
rect 36640 7134 36674 7214
rect 36700 7206 36708 7214
rect 37398 7134 37432 7214
rect 38156 7134 38190 7214
rect 38914 7134 38948 7214
rect 39672 7134 39706 7214
rect 40430 7134 40464 7214
rect 40614 7134 40648 7230
rect 19263 7100 40648 7134
rect 19088 6060 19134 6084
rect 7836 6028 7852 6032
rect 7864 6028 7908 6032
rect -2896 5990 5419 6026
rect 5438 6002 5454 6026
rect -2874 5792 -2847 5954
rect 3784 5920 5419 5990
rect 7852 5976 7864 6028
rect 14304 5920 14338 6039
rect 14406 6022 14464 6039
rect 14518 6022 14556 6039
rect 15064 6022 15122 6039
rect 15276 6022 15314 6039
rect 15722 6022 15780 6039
rect 16034 6022 16072 6039
rect 16380 6022 16438 6039
rect 16792 6022 16830 6039
rect 17038 6022 17096 6039
rect 17550 6022 17588 6039
rect 17678 6028 17754 6039
rect 17696 6022 17754 6028
rect 14406 5988 14556 6022
rect 14608 5988 15314 6022
rect 15366 5988 16072 6022
rect 16124 5988 16830 6022
rect 16882 5988 17588 6022
rect 17640 5988 17754 6022
rect 14406 5972 14464 5988
rect 15064 5972 15122 5988
rect 15722 5972 15780 5988
rect 16380 5972 16438 5988
rect 17038 5972 17096 5988
rect 17696 5972 17754 5988
rect 14406 5957 14421 5972
rect 14418 5920 14452 5954
rect 15076 5920 15110 5954
rect 15734 5920 15768 5954
rect 16392 5920 16426 5954
rect 17050 5920 17084 5972
rect 17739 5957 17754 5972
rect 17708 5920 17742 5954
rect 17822 5920 17856 6039
rect 19263 5920 22887 7100
rect 23492 6372 23954 7010
rect 23550 6288 23900 6322
rect 23550 5920 23584 6288
rect 23642 6258 23676 6288
rect 23682 6274 23726 6288
rect 23682 6258 23772 6272
rect 23642 6220 23780 6258
rect 23642 6182 23676 6220
rect 23708 6186 23780 6220
rect 23754 6182 23772 6186
rect 23642 6150 23682 6182
rect 23688 6178 23710 6182
rect 23754 6178 23764 6182
rect 23782 6154 23800 6288
rect 23782 6150 23792 6154
rect 23642 6136 23676 6150
rect 23688 6136 23698 6147
rect 23741 6136 23786 6147
rect 23642 6072 23698 6136
rect 23664 6060 23698 6072
rect 23752 6060 23786 6136
rect 23664 6022 23710 6060
rect 23740 6022 23798 6060
rect 23664 5988 23798 6022
rect 23664 5974 23710 5988
rect 23652 5972 23710 5974
rect 23740 5972 23798 5988
rect 23652 5960 23698 5972
rect 23652 5954 23692 5960
rect 23758 5954 23798 5972
rect 23652 5948 23698 5954
rect 23664 5944 23698 5948
rect 23752 5948 23798 5954
rect 23752 5944 23786 5948
rect 23674 5920 23776 5944
rect 23866 5920 23900 6288
rect 24370 6084 24404 7100
rect 24484 6142 24529 7100
rect 24370 6060 24440 6084
rect 24484 6060 24524 6142
rect 24370 5988 24388 6060
rect 24472 6022 24530 6060
rect 24542 6028 24552 7100
rect 25142 6142 25203 7100
rect 25800 6142 25845 7100
rect 25916 6142 25961 7100
rect 26458 6142 26503 7100
rect 25142 6084 25192 6142
rect 25142 6060 25198 6084
rect 25800 6060 25834 6142
rect 25916 6084 25950 6142
rect 25910 6072 25950 6084
rect 25910 6060 25956 6072
rect 26458 6060 26492 6142
rect 25130 6022 25182 6060
rect 25208 6022 25238 6028
rect 25788 6022 25846 6060
rect 25888 6028 25956 6060
rect 25854 6022 25956 6028
rect 26446 6022 26504 6060
rect 26534 6028 26562 7100
rect 26590 6028 26618 7100
rect 26674 6142 26719 7100
rect 27116 6142 27161 7100
rect 27432 6142 27477 7100
rect 27774 6142 27819 7100
rect 26674 6072 26708 6142
rect 27116 6060 27150 6142
rect 27432 6072 27466 6142
rect 27774 6060 27808 6142
rect 26646 6022 26684 6060
rect 27104 6022 27162 6060
rect 27404 6022 27442 6060
rect 27762 6022 27820 6060
rect 24472 6000 25182 6022
rect 25204 6000 25956 6022
rect 24472 5988 25176 6000
rect 25204 5988 25210 6000
rect 25220 5988 25926 6000
rect 25978 5988 26684 6022
rect 26736 5988 27442 6022
rect 27494 5988 27820 6022
rect 24370 5920 24404 5988
rect 24472 5972 24530 5988
rect 25130 5972 25176 5988
rect 25788 5972 25846 5988
rect 26446 5972 26504 5988
rect 27104 5972 27162 5988
rect 27762 5972 27820 5988
rect 24472 5957 24487 5972
rect 24484 5920 24518 5954
rect 25142 5920 25176 5972
rect 25800 5920 25834 5954
rect 26458 5920 26492 5972
rect 27805 5957 27820 5972
rect 27116 5920 27150 5954
rect 27774 5920 27808 5954
rect 27888 5920 27922 7100
rect 28184 6060 28230 6084
rect 28942 6060 28988 6084
rect 29700 6060 29746 6084
rect 30458 6072 30498 6084
rect 30458 6060 30504 6072
rect 30578 5982 30612 7100
rect -2836 5830 -2809 5916
rect 3784 5886 30516 5920
rect 3784 5850 5419 5886
rect -2874 5316 -2847 5478
rect -2836 5354 -2809 5440
rect -2754 5202 -2134 5624
rect -2084 5572 -1518 5606
rect -2084 5544 -2050 5572
rect -1552 5544 -1518 5572
rect -2118 5541 -2050 5544
rect -1586 5541 -1484 5544
rect -2084 5478 -2050 5541
rect -1713 5492 -1702 5503
rect -2084 5454 -2044 5478
rect -2029 5472 -1948 5477
rect -2036 5454 -1948 5472
rect -1889 5458 -1702 5492
rect -2084 5250 -2050 5454
rect -2029 5430 -1948 5454
rect -1701 5430 -1620 5477
rect -1982 5392 -1948 5430
rect -1654 5392 -1620 5430
rect -1713 5364 -1702 5375
rect -1889 5330 -1702 5364
rect -1552 5250 -1518 5541
rect -2084 5216 -1518 5250
rect -2754 4726 -2134 5148
rect -2084 5096 -1518 5130
rect -2084 5024 -2050 5096
rect -2084 5006 -1912 5024
rect -1713 5016 -1702 5027
rect -2084 4916 -2050 5006
rect -2029 4996 -1948 5001
rect -2036 4978 -1940 4996
rect -1889 4982 -1702 5016
rect -1690 5006 -1582 5008
rect -1701 4980 -1620 5001
rect -1701 4978 -1610 4980
rect -2036 4923 -2034 4978
rect -2029 4954 -1948 4978
rect -1701 4954 -1620 4978
rect -1982 4929 -1948 4954
rect -1654 4929 -1620 4954
rect -1998 4917 -1901 4929
rect -1701 4917 -1604 4929
rect -1998 4916 -1604 4917
rect -1552 4916 -1518 5096
rect -2084 4883 -1518 4916
rect -2084 4774 -2050 4883
rect -2036 4876 -2034 4877
rect -1889 4871 -1713 4883
rect -1889 4854 -1702 4871
rect -1552 4774 -1518 4883
rect -2084 4740 -1518 4774
rect 3236 4756 5241 4784
rect 5287 4756 5300 4784
rect -2908 4340 5308 4351
rect -2897 4328 5297 4340
rect -2908 4317 5308 4328
rect -2881 4271 -2847 4317
rect -2256 4308 -2248 4317
rect -2062 4308 -2056 4317
rect -2092 4259 -1438 4280
rect -2788 4213 5188 4259
rect -2788 4203 5199 4213
rect -2881 3607 -2847 4197
rect -2072 4182 -1418 4203
rect 942 4008 1390 4018
rect 934 3806 1390 4008
rect 934 3796 1382 3806
rect -1226 3612 -954 3639
rect 3878 3612 4334 3616
rect -2799 3601 5199 3612
rect 5247 3607 5281 4197
rect -2788 3591 5199 3601
rect -2788 3545 5188 3591
rect 3916 3531 4372 3545
rect 5213 3531 5315 3551
rect 5349 3531 5383 5850
rect -2881 3517 -2847 3521
rect 3319 3497 6775 3531
rect 3319 3487 3353 3497
rect 3542 3494 4894 3497
rect -2919 3467 5319 3487
rect 5349 3467 5383 3497
rect -2919 3453 5383 3467
rect -2890 3368 -2881 3402
rect -2908 3357 -1374 3368
rect -2897 3345 -1374 3357
rect -2908 3334 -1374 3345
rect -2983 3160 -2918 3272
rect -2881 3160 -2880 3334
rect -2800 3266 -2366 3313
rect -2208 3266 -2161 3313
rect -1550 3266 -1503 3313
rect -2776 3232 -2161 3266
rect -2118 3232 -1503 3266
rect -2876 3185 -2847 3211
rect -2838 3185 -2804 3194
rect -2876 3184 -2800 3185
rect -2876 3160 -2793 3184
rect -2191 3173 -2146 3184
rect -1533 3173 -1488 3184
rect -6114 3126 -2562 3160
rect -6114 2926 -6080 3126
rect -5804 3074 -5758 3105
rect -5816 3058 -5758 3074
rect -5938 3024 -5758 3058
rect -5816 2977 -5758 3024
rect -6011 2965 -5966 2976
rect -6000 2926 -5966 2965
rect -6256 2864 -5960 2926
rect -6114 2534 -6080 2864
rect -6000 2683 -5966 2864
rect -5804 2695 -5770 2977
rect -6012 2636 -5953 2683
rect -5832 2636 -5785 2683
rect -6012 2602 -5785 2636
rect -6012 2586 -5954 2602
rect -6012 2571 -5997 2586
rect -5690 2534 -5656 3126
rect -8586 2500 -5656 2534
rect -5306 2972 -5302 2977
rect -5306 2786 -5278 2972
rect -8586 2464 -6628 2500
rect -8566 2458 -8532 2464
rect -26468 2392 -8594 2426
rect -26468 2346 -12220 2392
rect -12182 2346 -12148 2392
rect -12120 2346 -8594 2392
rect -26468 2310 -8594 2346
rect -8592 2310 -8586 2458
rect -8566 2310 -8530 2458
rect -8254 2310 -6628 2464
rect -26468 2276 -6628 2310
rect -26468 2208 -8594 2276
rect -8592 2266 -8586 2276
rect -8566 2266 -8530 2276
rect -8566 2208 -8532 2266
rect -8254 2208 -6628 2276
rect -26468 2174 -6628 2208
rect -26468 2158 -8594 2174
rect -26470 1694 -8594 2158
rect -8566 1694 -8532 2174
rect -8254 1954 -6628 2174
rect -8254 1756 -6604 1954
rect -8128 1694 -8083 1756
rect -7510 1694 -7476 1756
rect -7470 1694 -7438 1756
rect -7396 1694 -7362 1756
rect -26470 918 -7300 1694
rect -28336 852 -7300 918
rect -7030 1664 -6628 1700
rect -6114 1664 -6080 2500
rect -5306 2100 -5302 2786
rect -5038 2038 -5004 3126
rect -4924 3089 -4877 3105
rect -4936 3058 -4877 3089
rect -4712 3058 -4665 3105
rect -4266 3074 -4219 3105
rect -4278 3058 -4219 3074
rect -4054 3058 -4007 3105
rect -3852 3058 -3460 3126
rect -4936 3024 -4665 3058
rect -4622 3024 -4007 3058
rect -3964 3024 -3460 3058
rect -4936 2977 -4878 3024
rect -4278 2977 -4220 3024
rect -4924 2199 -4890 2977
rect -4695 2965 -4650 2976
rect -4684 2187 -4650 2965
rect -4266 2199 -4232 2977
rect -4037 2966 -3992 2976
rect -4050 2830 -3972 2966
rect -3852 2830 -3460 3024
rect -3346 2990 -3328 3092
rect -3318 3018 -3272 3064
rect -2983 3058 -2918 3126
rect -2881 3105 -2793 3126
rect -2881 3058 -2791 3105
rect -2738 3058 -2691 3105
rect -2983 3024 -2691 3058
rect -4050 2778 -3460 2830
rect -4026 2684 -3460 2778
rect -4026 2187 -3992 2684
rect -4696 2140 -4637 2187
rect -4294 2140 -4247 2187
rect -4038 2140 -3979 2187
rect -3852 2182 -3460 2684
rect -3636 2140 -3589 2182
rect -4862 2106 -4247 2140
rect -4204 2106 -3589 2140
rect -4696 2090 -4638 2106
rect -4038 2090 -3980 2106
rect -4684 2038 -4644 2090
rect -3494 2038 -3460 2182
rect -5038 2004 -3460 2038
rect -2983 2906 -2918 3024
rect -2881 2977 -2792 3024
rect -2881 2949 -2847 2977
rect -2872 2933 -2847 2949
rect -2838 2921 -2804 2977
rect -2721 2965 -2676 2976
rect -2710 2921 -2676 2965
rect -2596 2921 -2562 3126
rect -2192 2933 -2191 2934
rect -2193 2932 -2192 2933
rect -2180 2921 -2146 3173
rect -2135 2933 -2134 2934
rect -1534 2933 -1533 2934
rect -2134 2932 -2133 2933
rect -1535 2932 -1534 2933
rect -1522 2921 -1488 3173
rect -1408 2921 -1374 3334
rect -848 3366 2704 3370
rect 3319 3366 3353 3453
rect 3448 3429 5200 3453
rect 5247 3429 5281 3453
rect 5349 3429 5383 3453
rect 6608 3435 6640 3448
rect 6664 3435 6668 3476
rect 3495 3395 4110 3429
rect 4153 3395 4768 3429
rect 4811 3402 5383 3429
rect 4811 3395 5391 3402
rect 5247 3370 5281 3395
rect 5318 3389 5391 3395
rect 5457 3389 5540 3402
rect 5988 3389 6049 3402
rect 6115 3389 6192 3402
rect 6640 3389 6664 3402
rect 5349 3370 5383 3389
rect 6608 3370 6640 3389
rect 6664 3370 6668 3389
rect -848 3336 4492 3366
rect 4738 3336 4794 3347
rect -848 2921 -814 3336
rect -104 3268 -57 3315
rect 554 3268 601 3315
rect 934 3268 1382 3336
rect 1598 3332 4492 3336
rect 1598 3268 1632 3332
rect 1870 3268 1917 3315
rect -672 3234 -57 3268
rect -14 3234 601 3268
rect 644 3264 1917 3268
rect 1944 3268 1960 3311
rect 2528 3268 2575 3315
rect 1944 3264 2575 3268
rect 2670 3311 2704 3332
rect 3319 3311 3353 3332
rect 3433 3314 3478 3332
rect 4091 3314 4136 3332
rect 3433 3311 3467 3314
rect 4091 3311 4125 3314
rect 2670 3264 2717 3311
rect 3000 3264 3047 3311
rect 3319 3264 3366 3311
rect 3433 3280 3480 3311
rect 3421 3264 3480 3280
rect 3658 3264 3705 3311
rect 4091 3280 4138 3311
rect 4079 3264 4138 3280
rect 4316 3264 4363 3311
rect 644 3234 3047 3264
rect -745 3175 -700 3186
rect -87 3175 -42 3186
rect 571 3175 616 3186
rect -734 2921 -700 3175
rect -689 2933 -688 2934
rect -88 2933 -87 2934
rect -688 2932 -687 2933
rect -89 2932 -88 2933
rect -76 2921 -42 3175
rect 582 3014 616 3175
rect 934 3130 1382 3234
rect 1216 3014 1294 3130
rect 1314 3014 1344 3066
rect -31 2933 -30 2934
rect 570 2933 571 2934
rect -30 2932 -29 2933
rect 569 2932 570 2933
rect 582 2927 622 3014
rect 1216 3010 1314 3014
rect 1344 3010 1370 3014
rect 1216 2996 1294 3010
rect 1314 2996 1344 3010
rect 627 2933 628 2934
rect 628 2932 629 2933
rect 582 2921 616 2927
rect 1214 2921 1382 2996
rect 1598 2984 1632 3234
rect 1774 3230 2389 3234
rect 2432 3230 3047 3234
rect 3090 3230 3705 3264
rect 3748 3230 4363 3264
rect 1886 3183 1944 3187
rect 2544 3183 2602 3187
rect 1701 3171 1746 3182
rect 1887 3175 1932 3183
rect 1598 2966 1668 2984
rect 1598 2928 1632 2966
rect 1598 2921 1668 2928
rect 1712 2921 1746 3171
rect 1898 2921 1932 3175
rect 2359 3171 2404 3182
rect 2545 3175 2590 3183
rect 2370 2921 2404 3171
rect 2556 2921 2590 3175
rect 2670 2921 2704 3230
rect 3017 3171 3062 3182
rect 3016 2933 3017 2934
rect 3015 2932 3016 2933
rect 3028 2921 3062 3171
rect 3064 2927 3068 3014
rect 3150 2966 3206 2984
rect 3073 2933 3074 2934
rect 3074 2932 3075 2933
rect 3150 2921 3206 2928
rect 3319 2921 3353 3230
rect 3421 3183 3479 3230
rect 4079 3183 4137 3230
rect 3433 2921 3467 3183
rect 3675 3171 3720 3182
rect 3686 2921 3720 3171
rect 4091 2926 4125 3183
rect 4333 3171 4378 3182
rect 3892 2921 4188 2926
rect 4344 2921 4378 3171
rect 4458 2921 4492 3332
rect 4749 3314 4794 3336
rect 5110 3336 6688 3370
rect 4737 2933 4738 2934
rect 4736 2932 4737 2933
rect 4749 2921 4783 3314
rect 4794 2933 4795 2934
rect 4795 2932 4796 2933
rect 5110 2921 5144 3336
rect 5247 3314 5328 3336
rect 5349 3315 5383 3336
rect 5407 3315 5417 3336
rect 6640 3333 6688 3336
rect 5247 3268 5281 3314
rect 5346 3268 6559 3315
rect 5247 3234 5901 3268
rect 5944 3234 6559 3268
rect 5247 3209 5281 3234
rect 5247 3186 5292 3209
rect 5213 3175 5292 3186
rect 5224 2949 5292 3175
rect 5224 2933 5269 2949
rect 5188 2921 5199 2932
rect -2983 2859 -2847 2906
rect -2983 2248 -2918 2859
rect -2881 2291 -2847 2859
rect -2872 2275 -2847 2291
rect -2838 2887 -2793 2921
rect -2788 2887 -1374 2921
rect -882 2887 5204 2921
rect 5224 2906 5258 2933
rect -2838 2263 -2804 2887
rect -2710 2263 -2676 2887
rect -2596 2263 -2562 2887
rect -2193 2875 -2192 2876
rect -2192 2874 -2191 2875
rect -2192 2275 -2191 2276
rect -2193 2274 -2192 2275
rect -2180 2263 -2146 2887
rect -2134 2875 -2133 2876
rect -1535 2875 -1534 2876
rect -2135 2874 -2134 2875
rect -1534 2874 -1533 2875
rect -1966 2684 -1716 2830
rect -1902 2570 -1748 2684
rect -2135 2275 -2134 2276
rect -1534 2275 -1533 2276
rect -2134 2274 -2133 2275
rect -1535 2274 -1534 2275
rect -1522 2263 -1488 2887
rect -1408 2263 -1374 2887
rect -848 2263 -814 2887
rect -734 2263 -700 2887
rect -688 2875 -687 2876
rect -89 2875 -88 2876
rect -689 2874 -688 2875
rect -88 2874 -87 2875
rect -689 2275 -688 2276
rect -88 2275 -87 2276
rect -688 2274 -687 2275
rect -89 2274 -88 2275
rect -76 2263 -42 2887
rect 582 2881 616 2887
rect -30 2875 -29 2876
rect 569 2875 570 2876
rect -31 2874 -30 2875
rect 570 2874 571 2875
rect 582 2836 622 2881
rect 628 2875 629 2876
rect 627 2874 628 2875
rect 582 2758 616 2836
rect 1214 2828 1382 2887
rect 1200 2826 1382 2828
rect 1598 2864 1668 2887
rect 1598 2836 1632 2864
rect 1200 2810 1234 2826
rect 1168 2790 1234 2800
rect 1240 2790 1274 2826
rect 1280 2810 1344 2826
rect 1598 2808 1668 2836
rect 622 2758 1274 2790
rect 1280 2782 1344 2800
rect 582 2696 1274 2758
rect 1288 2776 1344 2782
rect 1598 2776 1632 2808
rect 1712 2776 1746 2887
rect 1288 2754 1858 2776
rect 1292 2742 1858 2754
rect 1292 2696 1326 2742
rect 582 2647 1390 2696
rect 1598 2662 1632 2742
rect 1712 2679 1746 2742
rect 1824 2683 1858 2742
rect 1898 2774 1932 2887
rect 1898 2683 1943 2774
rect 2370 2695 2404 2887
rect 2556 2683 2590 2887
rect 2670 2683 2704 2887
rect 3015 2875 3016 2876
rect 3016 2874 3017 2875
rect 3010 2820 3020 2830
rect 3006 2800 3020 2820
rect 3028 2695 3062 2887
rect 3064 2830 3068 2881
rect 3074 2875 3075 2876
rect 3073 2874 3074 2875
rect 3150 2864 3206 2887
rect 3064 2820 3082 2830
rect 3064 2800 3086 2820
rect 3150 2808 3206 2836
rect 3319 2683 3353 2887
rect 3433 2692 3467 2887
rect 3686 2695 3720 2887
rect 3892 2864 4188 2887
rect 4091 2692 4125 2864
rect 4344 2820 4378 2887
rect 4334 2750 4386 2820
rect 4218 2694 4386 2750
rect 3433 2683 3478 2692
rect 4091 2683 4136 2692
rect 4218 2683 4354 2694
rect 1663 2662 1674 2673
rect 582 2562 1428 2647
rect 1487 2628 1674 2662
rect 582 2536 1418 2562
rect 582 2484 1390 2536
rect 1598 2534 1632 2628
rect 1675 2600 1756 2647
rect 1824 2636 2048 2683
rect 2342 2636 2389 2683
rect 2544 2636 2603 2683
rect 2670 2636 2717 2683
rect 3000 2636 3047 2683
rect 3306 2636 4363 2683
rect 1758 2602 2389 2636
rect 2432 2602 3047 2636
rect 3090 2602 3705 2636
rect 3748 2602 4363 2636
rect 1722 2546 1756 2600
rect 1663 2534 1674 2545
rect 1824 2534 1858 2602
rect 1886 2586 1944 2602
rect 2544 2586 2602 2602
rect 1898 2534 1943 2586
rect 2556 2534 2590 2586
rect 2670 2534 2704 2602
rect 3319 2534 3353 2602
rect 3421 2586 3479 2602
rect 4079 2586 4137 2602
rect 3433 2534 3478 2586
rect 4091 2534 4136 2586
rect 4458 2534 4492 2887
rect 4736 2875 4737 2876
rect 4737 2874 4738 2875
rect 1487 2500 4492 2534
rect 4749 2692 4783 2887
rect 4795 2875 4796 2876
rect 4794 2874 4795 2875
rect 582 2368 1274 2484
rect 1292 2420 1326 2484
rect 1824 2420 1858 2500
rect 1292 2386 1858 2420
rect 582 2276 627 2368
rect -31 2275 -30 2276
rect 570 2275 571 2276
rect 582 2275 628 2276
rect 1228 2275 1229 2276
rect -30 2274 -29 2275
rect 569 2274 570 2275
rect 480 2263 570 2274
rect 582 2263 616 2275
rect 628 2274 629 2275
rect 1227 2274 1228 2275
rect 628 2263 698 2274
rect 1240 2263 1274 2368
rect 1898 2276 1943 2500
rect 1285 2275 1286 2276
rect 1886 2275 1887 2276
rect 1898 2275 1944 2276
rect 2544 2275 2545 2276
rect 1286 2274 1287 2275
rect 1885 2274 1886 2275
rect 1826 2263 1886 2274
rect 1898 2263 1932 2275
rect 1944 2274 1945 2275
rect 2543 2274 2544 2275
rect 1944 2263 2048 2274
rect 2556 2263 2590 2500
rect 2670 2263 2704 2500
rect 3319 2263 3353 2500
rect 3433 2276 3478 2500
rect 4074 2284 4144 2500
rect 3433 2275 3479 2276
rect 3433 2263 3467 2275
rect 3479 2274 3480 2275
rect 3900 2274 4356 2284
rect 4749 2276 4794 2692
rect 4737 2275 4738 2276
rect 4749 2275 4795 2276
rect 4736 2274 4737 2275
rect 3479 2263 4737 2274
rect 4749 2263 4783 2275
rect 4795 2274 4796 2275
rect 5110 2274 5144 2887
rect 5211 2859 5281 2906
rect 5224 2692 5292 2859
rect 5224 2291 5328 2692
rect 4795 2263 5199 2274
rect -2983 2201 -2847 2248
rect -2983 2036 -2918 2201
rect -2881 2070 -2847 2201
rect -2838 2229 -2793 2263
rect -2788 2240 -1374 2263
rect -882 2242 2704 2263
rect 3285 2242 5199 2263
rect 5224 2248 5269 2291
rect 5211 2246 5328 2248
rect -882 2240 5199 2242
rect -2788 2229 5199 2240
rect -2838 2197 -2804 2229
rect -2776 2223 -2740 2229
rect -2838 2181 -2813 2197
rect -2776 2190 -2772 2223
rect -2710 2185 -2676 2229
rect -2596 2185 -2562 2229
rect -2242 2223 -2086 2229
rect -1588 2223 -740 2229
rect -2193 2217 -2192 2218
rect -2192 2216 -2191 2217
rect -2186 2185 -2140 2223
rect -2134 2217 -2133 2218
rect -2135 2216 -2134 2217
rect -1550 2196 -1456 2223
rect -1548 2188 -1458 2196
rect -1528 2185 -1482 2188
rect -2776 2162 -2744 2184
rect -2722 2138 -2663 2185
rect -2596 2138 -2549 2185
rect -2208 2184 -2161 2185
rect -1550 2184 -1503 2185
rect -2214 2157 -2112 2184
rect -1578 2168 -1428 2184
rect -1576 2160 -1430 2168
rect -1556 2157 -1454 2160
rect -2208 2138 -2161 2157
rect -1550 2138 -1503 2157
rect -2776 2104 -2161 2138
rect -2118 2104 -1503 2138
rect -2722 2088 -2664 2104
rect -2890 2036 -2847 2070
rect -2710 2036 -2676 2088
rect -2596 2036 -2562 2104
rect -1408 2036 -1374 2223
rect -7030 1630 -4758 1664
rect -7030 888 -6628 1630
rect -6178 1266 -6156 1476
rect -6114 888 -6080 1630
rect -6012 1562 -5932 1609
rect -5592 1562 -5545 1609
rect -5342 1578 -5295 1609
rect -5354 1562 -5295 1578
rect -4934 1562 -4887 1609
rect -6012 1528 -5545 1562
rect -5502 1528 -4887 1562
rect -6012 1481 -5954 1528
rect -5354 1481 -5296 1528
rect -6000 888 -5955 1481
rect -5575 1469 -5530 1480
rect -5564 1192 -5530 1469
rect -5342 1192 -5308 1481
rect -4917 1469 -4872 1480
rect -4906 1192 -4872 1469
rect -7030 852 -5918 888
rect -28336 818 -5918 852
rect -28336 749 -7300 818
rect -7030 749 -5918 818
rect -28336 712 -5918 749
rect -28336 678 -5656 712
rect -28336 610 -5918 678
rect -5832 610 -5785 657
rect -28336 576 -5785 610
rect -28336 434 -5918 576
rect -5815 517 -5770 528
rect -5804 481 -5770 517
rect -5804 434 -5757 481
rect -5690 434 -5656 678
rect -5564 660 -5519 1192
rect -5342 660 -5297 1192
rect -4906 716 -4861 1192
rect -4792 716 -4758 1630
rect -4684 1550 -4644 2004
rect -2983 2002 -1374 2036
rect -2983 1970 -2949 2002
rect -2881 1970 -2847 2002
rect -2710 1970 -2676 2002
rect -2596 1970 -2562 2002
rect -848 1970 -814 2223
rect -734 1970 -700 2229
rect -694 2223 -634 2229
rect -138 2223 -82 2229
rect -688 2217 -687 2218
rect -89 2217 -88 2218
rect -689 2216 -688 2217
rect -88 2216 -87 2217
rect -76 1970 -42 2229
rect -36 2223 16 2229
rect -40 2184 -36 2223
rect -30 2217 -29 2218
rect 569 2217 570 2218
rect 582 2217 616 2229
rect 628 2217 629 2218
rect 1227 2217 1228 2218
rect -31 2216 -30 2217
rect 570 2216 571 2217
rect 582 2216 628 2217
rect 1228 2216 1229 2217
rect 582 2020 627 2216
rect 582 1970 616 2020
rect 1240 2000 1274 2229
rect 1840 2223 1892 2229
rect 1286 2217 1287 2218
rect 1285 2216 1286 2217
rect 1316 2188 1332 2223
rect 1288 2130 1332 2188
rect 1344 2130 1388 2223
rect 1885 2217 1886 2218
rect 1898 2217 1932 2229
rect 1938 2223 1994 2229
rect 2490 2223 2550 2229
rect 1944 2217 1945 2218
rect 2543 2217 2544 2218
rect 1886 2216 1887 2217
rect 1898 2216 1944 2217
rect 2544 2216 2545 2217
rect 1898 2002 1943 2216
rect 934 1970 1382 2000
rect 1898 1970 1932 2002
rect 2556 1970 2590 2229
rect 2596 2223 3292 2229
rect 2670 1970 2704 2223
rect 3236 2167 3292 2186
rect 3319 1970 3353 2229
rect 3433 2217 3467 2229
rect 3479 2217 3480 2218
rect 3433 2216 3479 2217
rect 3433 1970 3478 2216
rect 3900 2214 4356 2229
rect 4736 2217 4737 2218
rect 4749 2217 4783 2229
rect 4795 2217 4796 2218
rect 4737 2216 4738 2217
rect 4749 2216 4795 2217
rect 4074 2064 4144 2214
rect 4091 1970 4136 2064
rect 4749 1970 4794 2216
rect 5110 2038 5144 2229
rect 5200 2199 5328 2246
rect 5247 2187 5328 2199
rect 5349 2187 5383 3234
rect 5395 3187 5453 3234
rect 6053 3187 6111 3234
rect 5407 2187 5452 3187
rect 5871 3175 5927 3186
rect 5882 2199 5927 3175
rect 6065 2187 6110 3187
rect 6529 3175 6585 3186
rect 6540 2199 6585 3175
rect 5239 2140 6559 2187
rect 5247 2106 5901 2140
rect 5944 2106 6559 2140
rect 5247 2051 5328 2106
rect 5200 2038 5328 2051
rect 5349 2038 5383 2106
rect 5395 2090 5453 2106
rect 6053 2090 6111 2106
rect 5407 2038 5417 2090
rect 6608 2038 6640 2048
rect 6654 2038 6688 3333
rect 5110 2004 6688 2038
rect 5247 1970 5328 2004
rect 5349 1970 5383 2004
rect 5407 1970 5417 2004
rect -2996 1576 5424 1970
rect -4706 1538 -4698 1550
rect -4710 1286 -4698 1538
rect -4706 1274 -4698 1286
rect -4704 1264 -4698 1274
rect -4684 1264 -4650 1550
rect -4684 716 -4644 1264
rect -2996 1248 5441 1576
rect 5448 1286 5479 1538
rect -2996 877 5424 1248
rect 6608 877 6640 2004
rect 6664 877 6668 2004
rect 6723 1876 6757 3336
rect 6837 1876 6871 3435
rect 6906 3404 6907 3567
rect 9476 3536 9510 3964
rect 9590 3536 9624 3570
rect 10248 3536 10282 3570
rect 10362 3536 10396 3964
rect 10666 3536 10700 3964
rect 10780 3536 10814 3570
rect 11438 3536 11472 3570
rect 11552 3536 11586 3964
rect 8486 3502 11846 3536
rect 9476 3406 9510 3502
rect 10242 3472 10244 3476
rect 9578 3406 9830 3472
rect 9844 3434 10294 3472
rect 9882 3406 10294 3434
rect 10362 3406 10396 3502
rect 10666 3406 10700 3502
rect 10768 3406 11146 3472
rect 11160 3434 11484 3472
rect 11198 3406 11484 3434
rect 11552 3406 11586 3502
rect 11976 3406 11996 3590
rect 14304 3585 14338 5886
rect 16392 5490 16426 5886
rect 15950 5252 16664 5490
rect 17050 5252 17084 5886
rect 15942 4880 17122 5252
rect 16392 3586 16426 4880
rect 17050 3586 17084 4880
rect 17674 4054 17698 4344
rect 17708 4054 17732 4344
rect 14406 3585 17754 3586
rect 14304 3567 17754 3585
rect 12862 3406 12896 3424
rect 7160 1966 7161 3404
rect 7906 2172 7908 2200
rect 7906 2158 7980 2172
rect 7990 2158 8062 2172
rect 7906 2102 7952 2144
rect 8018 2102 8062 2144
rect 8354 1966 8810 3404
rect 9264 3402 12896 3406
rect 9084 3394 9146 3402
rect 9212 3394 12896 3402
rect 6723 1172 7104 1876
rect 6723 877 6757 1172
rect -2996 843 6769 877
rect -2996 822 5424 843
rect 6608 822 6640 843
rect 6664 822 6668 843
rect 6723 822 6757 843
rect -2996 775 6757 822
rect -2996 763 5424 775
rect -2996 750 -2526 763
rect -5038 682 -3460 716
rect -5564 493 -5530 660
rect -5342 481 -5308 660
rect -5592 434 -5545 481
rect -5354 434 -5295 481
rect -5038 434 -5004 682
rect -4906 660 -4861 682
rect -4792 661 -4758 682
rect -4684 661 -4644 682
rect -4906 614 -4872 660
rect -4805 614 -4430 661
rect -4294 614 -4247 661
rect -4039 614 -3589 661
rect -4906 580 -4247 614
rect -4204 584 -3589 614
rect -3494 584 -3460 682
rect -4204 580 -3460 584
rect -4906 532 -4872 580
rect -4935 521 -4872 532
rect -4924 493 -4872 521
rect -4924 481 -4879 493
rect -4934 477 -4879 481
rect -4934 434 -4887 477
rect -28336 400 -5545 434
rect -5502 400 -4887 434
rect -28336 332 -5918 400
rect -5804 332 -5770 400
rect -5690 332 -5656 400
rect -5354 384 -5296 400
rect -5306 332 -5302 384
rect -5038 332 -5004 400
rect -4924 332 -4890 400
rect -4792 332 -4758 580
rect -4696 533 -4638 580
rect -4038 533 -3980 580
rect -28336 298 -4758 332
rect -28336 246 -5918 298
rect -28336 216 -8594 246
rect -8586 216 -5918 246
rect -28336 210 -5918 216
rect -28336 188 -8594 210
rect -8586 188 -5918 210
rect -28336 182 -5918 188
rect -28336 166 -8594 182
rect -8586 166 -5918 182
rect -28336 132 -5918 166
rect -28336 88 -8594 132
rect -28336 -94 -12220 88
rect -12182 -94 -12148 88
rect -12120 -30 -8594 88
rect -8586 96 -5918 132
rect -5804 124 -5770 298
rect -5690 124 -5656 298
rect -5306 124 -5302 298
rect -5038 124 -5004 298
rect -4924 124 -4890 298
rect -4684 236 -4639 533
rect -4277 521 -4232 532
rect -4684 128 -4650 236
rect -4266 128 -4232 521
rect -4026 176 -3981 533
rect -3852 176 -3460 580
rect -4026 128 -3460 176
rect -2996 546 -1338 750
rect -884 748 2848 763
rect 3118 748 5424 763
rect -884 716 5424 748
rect 5429 716 5447 775
rect 5457 741 6084 775
rect 5457 735 5475 741
rect 6031 735 6049 741
rect 6059 716 6077 741
rect 6087 716 6105 775
rect 6115 741 6757 775
rect 6115 735 6133 741
rect 6608 716 6640 735
rect 6664 716 6668 735
rect -884 682 6688 716
rect -884 661 5424 682
rect -884 614 6452 661
rect 6512 614 6559 661
rect -884 580 5901 614
rect 5944 580 6559 614
rect -2996 532 -1082 546
rect -884 533 5453 580
rect 6053 533 6111 580
rect -2996 128 -1338 532
rect -12120 -80 -8592 -30
rect -12120 -94 -8594 -80
rect -28336 -118 -8594 -94
rect -8586 -118 -6080 96
rect -6034 -18 -6014 96
rect -6000 29 -5966 96
rect -6012 0 -5954 29
rect -6012 -18 -5953 0
rect -5916 -18 -4890 124
rect -6012 -52 -4890 -18
rect -28336 -120 -6080 -118
rect -6034 -120 -6014 -52
rect -6012 -68 -5954 -52
rect -6012 -83 -5980 -68
rect -6000 -120 -5980 -83
rect -5916 -120 -4890 -52
rect -28336 -152 -4890 -120
rect -28336 -182 -8594 -152
rect -8586 -154 -4890 -152
rect -8586 -182 -6080 -154
rect -28336 -190 -6080 -182
rect -28336 -220 -7888 -190
rect -7874 -220 -7230 -190
rect -7216 -220 -6572 -190
rect -28336 -254 -8532 -220
rect -8494 -254 -7888 -220
rect -7836 -254 -7230 -220
rect -7178 -254 -6572 -220
rect -28336 -344 -8594 -254
rect -8566 -293 -8532 -254
rect -8566 -344 -8511 -293
rect -8358 -344 -8324 -254
rect -8256 -292 -8198 -254
rect -8244 -344 -8199 -292
rect -8128 -344 -8083 -254
rect -7598 -292 -7540 -254
rect -7482 -292 -7404 -254
rect -7909 -304 -7853 -293
rect -7898 -344 -7853 -304
rect -7586 -344 -7541 -292
rect -7472 -344 -7404 -292
rect -7251 -304 -7195 -293
rect -28336 -378 -7362 -344
rect -28336 -408 -8594 -378
rect -8566 -408 -8511 -378
rect -8358 -408 -8324 -378
rect -8244 -408 -8199 -378
rect -8128 -408 -8083 -378
rect -7898 -408 -7853 -378
rect -7586 -408 -7541 -378
rect -28336 -480 -7500 -408
rect -28336 -960 -8594 -480
rect -8568 -518 -8510 -480
rect -8566 -826 -8511 -518
rect -8486 -722 -8428 -588
rect -8426 -722 -8368 -588
rect -8566 -960 -8522 -826
rect -8358 -960 -8324 -480
rect -8244 -826 -8199 -480
rect -8128 -826 -8083 -480
rect -8244 -960 -8210 -826
rect -8128 -960 -8094 -826
rect -7898 -960 -7853 -480
rect -7586 -960 -7541 -480
rect -7472 -519 -7404 -378
rect -7521 -530 -7404 -519
rect -7510 -960 -7404 -530
rect -7396 -960 -7362 -378
rect -28336 -1324 -7300 -960
rect -28676 -1634 -7300 -1324
rect -7240 -1634 -7195 -304
rect -28676 -1772 -7195 -1634
rect -28336 -1802 -7195 -1772
rect -7048 -954 -7014 -254
rect -6946 -292 -6888 -254
rect -6934 -826 -6889 -292
rect -6812 -826 -6767 -254
rect -6934 -954 -6900 -826
rect -6812 -954 -6778 -826
rect -6698 -954 -6664 -254
rect -6593 -304 -6537 -293
rect -6582 -826 -6537 -304
rect -6582 -954 -6548 -826
rect -6468 -954 -6434 -190
rect -6282 -954 -6280 -190
rect -6150 -954 -6080 -190
rect -6034 -826 -6014 -154
rect -6000 -860 -5980 -154
rect -5916 -455 -4890 -154
rect -4756 92 -1338 128
rect -884 236 5452 533
rect 5871 521 5916 532
rect -884 128 5441 236
rect 5882 128 5916 521
rect 6065 128 6099 533
rect 6529 521 6574 532
rect 6540 128 6574 521
rect 6608 128 6640 682
rect 6654 620 6688 682
rect 6654 128 6696 620
rect 6723 128 6757 741
rect 6837 336 6871 1172
rect 6906 750 6907 1004
rect 8390 750 8424 1966
rect 9162 1530 9196 3350
rect 9264 2738 12896 3394
rect 13288 3090 13298 3448
rect 13431 3429 14100 3567
rect 14268 3552 17754 3567
rect 14268 3518 17531 3552
rect 17674 3522 17698 3542
rect 17708 3522 17742 3552
rect 17674 3518 17742 3522
rect 14268 3494 17742 3518
rect 14268 3484 17531 3494
rect 17680 3490 17742 3494
rect 17674 3484 17742 3490
rect 14268 3450 17742 3484
rect 14118 3435 14146 3448
rect 14174 3435 14202 3448
rect 14268 3429 17531 3450
rect 17674 3444 17692 3450
rect 13431 3395 17531 3429
rect 17702 3416 17742 3450
rect 17702 3404 17704 3416
rect 13431 3347 14100 3395
rect 14146 3389 14174 3395
rect 13288 2876 13316 3090
rect 13288 2870 13298 2876
rect 9264 2668 12888 2738
rect 9232 1682 9254 2158
rect 9264 2034 11978 2668
rect 12040 2486 12044 2668
rect 12818 2486 12852 2668
rect 13431 2660 14102 3347
rect 14118 3346 14146 3389
rect 14174 3346 14202 3389
rect 14268 3347 17531 3395
rect 14228 3336 17531 3347
rect 17678 3346 17704 3404
rect 13467 2486 13501 2660
rect 13581 2486 13615 2520
rect 13943 2486 13977 2660
rect 14057 2486 14102 2660
rect 14239 2828 17531 3336
rect 17708 2866 17742 3416
rect 17680 2828 17742 2866
rect 14239 2794 17742 2828
rect 14239 2726 17531 2794
rect 17708 2726 17742 2794
rect 14239 2692 17754 2726
rect 17760 2692 17776 2726
rect 14239 2486 17531 2692
rect 12030 2452 17531 2486
rect 12030 2352 12064 2452
rect 12159 2384 12750 2431
rect 12082 2352 12086 2359
rect 12030 2296 12086 2352
rect 12206 2350 12750 2384
rect 12692 2303 12750 2350
rect 12818 2325 12852 2452
rect 12030 2034 12064 2296
rect 12080 2034 12086 2296
rect 12108 2034 12114 2296
rect 12133 2291 12189 2302
rect 12144 2034 12189 2291
rect 12704 2034 12749 2303
rect 12796 2034 12800 2303
rect 12818 2034 12870 2325
rect 13384 2302 13398 2344
rect 13426 2288 13440 2302
rect 13467 2291 13501 2452
rect 13943 2431 13977 2452
rect 14057 2431 14102 2452
rect 13569 2418 14104 2431
rect 13522 2350 13539 2384
rect 13569 2350 14124 2418
rect 13569 2303 13627 2350
rect 9162 1500 9202 1530
rect 9264 1518 12932 2034
rect 13396 2026 13398 2272
rect 13424 2026 13426 2244
rect 13460 2218 13501 2291
rect 13581 2218 13626 2303
rect 13432 2040 13776 2218
rect 13460 2026 13501 2040
rect 13581 2026 13626 2040
rect 13943 2026 13977 2350
rect 14045 2303 14103 2350
rect 14057 2026 14102 2303
rect 14107 2291 14163 2302
rect 9228 1502 12932 1518
rect 9222 1500 12932 1502
rect 9162 882 9196 1500
rect 9228 1392 12932 1500
rect 9228 1262 9234 1392
rect 9264 1084 12932 1392
rect 13108 1303 14102 2026
rect 14118 1315 14163 2291
rect 14174 1962 14214 2158
rect 14174 1512 14186 1962
rect 14118 1303 14158 1308
rect 14174 1303 14186 1308
rect 13108 1290 14103 1303
rect 14118 1290 14146 1303
rect 13108 1222 14146 1290
rect 13108 1206 14103 1222
rect 13108 1154 14102 1206
rect 14118 1154 14146 1222
rect 14174 1154 14202 1303
rect 14232 1227 17531 2452
rect 14228 1216 17531 1227
rect 14232 1154 17531 1216
rect 13108 1120 17531 1154
rect 13108 1084 14102 1120
rect 9264 882 12896 1084
rect 8492 848 12896 882
rect 9162 818 9196 848
rect 9264 818 12896 848
rect 8528 814 12896 818
rect 8526 780 12896 814
rect 8526 750 8544 780
rect 8554 750 9202 780
rect 7160 336 7161 750
rect 8354 746 9202 750
rect 7944 350 7962 526
rect 8354 336 8810 746
rect 9128 740 9146 746
rect 9156 712 9202 746
rect 9212 746 12896 780
rect 9212 740 9230 746
rect 6814 312 8810 336
rect 6837 280 6871 312
rect 7160 280 7161 312
rect 8354 280 8810 312
rect 6814 256 8810 280
rect 6837 128 6871 256
rect 7160 128 7161 256
rect 8354 128 8810 256
rect -4756 58 -1168 92
rect -4756 28 -1338 58
rect -4756 -44 -1306 28
rect -4756 -54 -1338 -44
rect -4756 -70 -1248 -54
rect -4756 -154 -1338 -70
rect -1322 -83 -1276 -82
rect -1327 -94 -1276 -83
rect -1322 -98 -1276 -94
rect -1328 -142 -1327 -141
rect -1329 -143 -1328 -142
rect -1322 -148 -1320 -98
rect -1316 -154 -1282 -98
rect -1202 -154 -1168 58
rect -4756 -188 -1168 -154
rect -5916 -616 -4924 -455
rect -4756 -514 -1338 -188
rect -1329 -200 -1328 -199
rect -1328 -201 -1327 -200
rect -1322 -286 -1320 -194
rect -4862 -548 -1338 -514
rect -4756 -616 -1338 -548
rect -7048 -990 -6080 -954
rect -5956 -990 -5936 -618
rect -5916 -650 -1338 -616
rect -5916 -990 -4924 -650
rect -4756 -688 -1338 -650
rect -4756 -720 -2526 -688
rect -1974 -720 -1940 -688
rect -1316 -720 -1282 -188
rect -1202 -720 -1168 -188
rect -884 -190 6907 128
rect -884 -720 2740 -190
rect 3100 -720 3134 -190
rect 3214 -720 3248 -190
rect 3252 -286 3270 -194
rect 3283 -720 6907 -190
rect 7160 92 8810 128
rect 7160 58 8980 92
rect 7160 28 8810 58
rect 7160 -44 8842 28
rect 7160 -688 8810 -44
rect 8821 -94 8866 -83
rect -4756 -754 6907 -720
rect -4756 -812 -2526 -754
rect -2040 -790 -1980 -776
rect -1974 -794 -1940 -754
rect -1934 -790 -1874 -776
rect -1376 -790 -1322 -776
rect -2092 -812 -1438 -794
rect -1328 -800 -1327 -799
rect -1329 -801 -1328 -800
rect -1316 -812 -1282 -754
rect -1202 -812 -1168 -754
rect -884 -812 2740 -754
rect 3100 -812 3134 -754
rect 3214 -812 3248 -754
rect 3252 -806 3254 -754
rect 3259 -800 3260 -799
rect 3260 -801 3261 -800
rect 3283 -812 6907 -754
rect -4756 -868 6907 -812
rect -7048 -1024 -4758 -990
rect -7048 -1092 -6080 -1024
rect -6006 -1026 -5936 -1024
rect -5916 -1070 -4924 -1024
rect -4792 -1070 -4758 -1024
rect -5938 -1092 -4758 -1070
rect -7048 -1104 -4758 -1092
rect -7048 -1126 -4924 -1104
rect -7048 -1172 -6080 -1126
rect -5916 -1151 -4924 -1126
rect -5916 -1172 -4838 -1151
rect -4792 -1172 -4758 -1104
rect -4756 -1172 -2526 -868
rect -2056 -892 -1402 -868
rect -7048 -1206 -2526 -1172
rect -7048 -1670 -6092 -1206
rect -5916 -1382 -4908 -1206
rect -5916 -1670 -4924 -1382
rect -7048 -1704 -4924 -1670
rect -7048 -1725 -6092 -1704
rect -7048 -1766 -6032 -1725
rect -6030 -1766 -5983 -1725
rect -7048 -1802 -5918 -1766
rect -28336 -1812 -5918 -1802
rect -5916 -1812 -4924 -1704
rect -4912 -1764 -4908 -1382
rect -4792 -1562 -4758 -1206
rect -4756 -1242 -2526 -1206
rect -4756 -1562 -4722 -1242
rect -4720 -1562 -4686 -1242
rect -4606 -1390 -4572 -1242
rect -4606 -1506 -4566 -1390
rect -4606 -1526 -4544 -1506
rect -4606 -1562 -4572 -1526
rect -4812 -1582 -4544 -1562
rect -4906 -1812 -4880 -1786
rect -28336 -1816 -4868 -1812
rect -28336 -1836 -5918 -1816
rect -28336 -1905 -7195 -1836
rect -7132 -1905 -7108 -1850
rect -28336 -1916 -7108 -1905
rect -7098 -1905 -7074 -1850
rect -7048 -1868 -5918 -1836
rect -7030 -1905 -5918 -1868
rect -5916 -1820 -4924 -1816
rect -5916 -1896 -4914 -1820
rect -7098 -1916 -5918 -1905
rect -28336 -1950 -5918 -1916
rect -28336 -2272 -7195 -1950
rect -28336 -2322 -7300 -2272
rect -28336 -2363 -7268 -2322
rect -7240 -2363 -7195 -2272
rect -7132 -2363 -7108 -1950
rect -28336 -2374 -7108 -2363
rect -7098 -2363 -7074 -1950
rect -7030 -2202 -5918 -1950
rect -5888 -2202 -5854 -1896
rect -7030 -2236 -5854 -2202
rect -5768 -2202 -5734 -1896
rect -5654 -2041 -5609 -1896
rect -5600 -1910 -5586 -1896
rect -5564 -1910 -5530 -1896
rect -5526 -1910 -5481 -1896
rect -5412 -1910 -5378 -1896
rect -5628 -2053 -5614 -2041
rect -5600 -2053 -5248 -1910
rect -5639 -2088 -5248 -2053
rect -5639 -2100 -5502 -2088
rect -5592 -2110 -5502 -2100
rect -5618 -2166 -5502 -2110
rect -5618 -2173 -5518 -2166
rect -5618 -2174 -5528 -2173
rect -5626 -2188 -5514 -2186
rect -5412 -2202 -5378 -2088
rect -5768 -2213 -5565 -2202
rect -5529 -2213 -5378 -2202
rect -5768 -2214 -5576 -2213
rect -5518 -2214 -5378 -2213
rect -4988 -2214 -4964 -2180
rect -4940 -2208 -4914 -1896
rect -4906 -2177 -4880 -1816
rect -4960 -2211 -4914 -2208
rect -4960 -2214 -4936 -2211
rect -5768 -2216 -5378 -2214
rect -5768 -2225 -5576 -2216
rect -5518 -2225 -5378 -2216
rect -5768 -2236 -5565 -2225
rect -5529 -2236 -5378 -2225
rect -7030 -2286 -5918 -2236
rect -4792 -2260 -4758 -1582
rect -7030 -2363 -5840 -2286
rect -7098 -2374 -5840 -2363
rect -28336 -2392 -5840 -2374
rect -5786 -2392 -5364 -2286
rect -4756 -2392 -4722 -1582
rect -28336 -2408 -6400 -2392
rect -6392 -2396 -6334 -2392
rect -6260 -2408 -6158 -2392
rect -28757 -2648 -28712 -2458
rect -29142 -2680 -28712 -2648
rect -28336 -2488 -17288 -2408
rect -17191 -2458 -8590 -2408
rect -8566 -2458 -8522 -2408
rect -17191 -2488 -8594 -2458
rect -8566 -2488 -8511 -2458
rect -8128 -2488 -8060 -2408
rect -7974 -2422 -7584 -2408
rect -7974 -2424 -7853 -2422
rect -7942 -2444 -7853 -2424
rect -7936 -2458 -7853 -2444
rect -7898 -2474 -7853 -2458
rect -8014 -2488 -7912 -2474
rect -7898 -2488 -7824 -2474
rect -7778 -2488 -7744 -2422
rect -7618 -2488 -7584 -2422
rect -7494 -2424 -7388 -2408
rect -7470 -2458 -7388 -2424
rect -7470 -2474 -7425 -2458
rect -7538 -2488 -7348 -2474
rect -7302 -2488 -7268 -2408
rect -7240 -2488 -7195 -2408
rect -7132 -2458 -7108 -2408
rect -7098 -2458 -7074 -2408
rect -6812 -2488 -6767 -2408
rect -6698 -2488 -6664 -2408
rect -6656 -2484 -6642 -2414
rect -6628 -2470 -6586 -2414
rect -6588 -2484 -6586 -2470
rect -6656 -2488 -6588 -2484
rect -6582 -2488 -6548 -2408
rect -6468 -2428 -6434 -2408
rect -6542 -2470 -6428 -2428
rect -6468 -2484 -6434 -2470
rect -6542 -2488 -6400 -2484
rect -6226 -2488 -6192 -2408
rect -6144 -2414 -6128 -2392
rect -6118 -2458 -6086 -2392
rect -6084 -2458 -6052 -2424
rect -6022 -2426 -6018 -2424
rect -5988 -2426 -5954 -2392
rect -6036 -2458 -6034 -2441
rect -5988 -2458 -5987 -2426
rect -6146 -2488 -6044 -2474
rect -28336 -2496 -6025 -2488
rect -28336 -2522 -5978 -2496
rect -5960 -2522 -5954 -2426
rect -29142 -2682 -28723 -2680
rect -29142 -3180 -29108 -2682
rect -28939 -2703 -28905 -2682
rect -28939 -2750 -28892 -2703
rect -28966 -2784 -28892 -2750
rect -28939 -2832 -28905 -2784
rect -28900 -2832 -28871 -2827
rect -29039 -2843 -28994 -2832
rect -29028 -3019 -28994 -2843
rect -28939 -2843 -28866 -2832
rect -28862 -2836 -28834 -2682
rect -28806 -2836 -28723 -2682
rect -28939 -3031 -28905 -2843
rect -28900 -3019 -28866 -2843
rect -28900 -3031 -28871 -3019
rect -28939 -3035 -28871 -3031
rect -28786 -3032 -28723 -2836
rect -28939 -3078 -28892 -3035
rect -28966 -3112 -28892 -3078
rect -28939 -3180 -28905 -3112
rect -28862 -3180 -28834 -3032
rect -28806 -3180 -28723 -3032
rect -29142 -3214 -28723 -3180
rect -28939 -3264 -28905 -3214
rect -28862 -3264 -28834 -3214
rect -28806 -3264 -28778 -3214
rect -28757 -3264 -28723 -3214
rect -29156 -3808 -28723 -3264
rect -28336 -2838 -17288 -2522
rect -17191 -2558 -8594 -2522
rect -17191 -2566 -12220 -2558
rect -17214 -2838 -12220 -2566
rect -28336 -2910 -12220 -2838
rect -28336 -2978 -17288 -2910
rect -17214 -2978 -12220 -2910
rect -28336 -3001 -12220 -2978
rect -12182 -3001 -12148 -2558
rect -12120 -2610 -8594 -2558
rect -8566 -2610 -8511 -2522
rect -8128 -2582 -8060 -2522
rect -7980 -2582 -7935 -2522
rect -7898 -2582 -7847 -2522
rect -7778 -2582 -7744 -2522
rect -7618 -2582 -7584 -2522
rect -7504 -2582 -7425 -2522
rect -8358 -2610 -7425 -2582
rect -7416 -2610 -7371 -2522
rect -7302 -2610 -7268 -2522
rect -7240 -2610 -7195 -2522
rect -6812 -2574 -6767 -2522
rect -6698 -2574 -6664 -2522
rect -6582 -2574 -6548 -2522
rect -6468 -2574 -6434 -2522
rect -6226 -2574 -6192 -2522
rect -7048 -2608 -6192 -2574
rect -6149 -2608 -6128 -2574
rect -7048 -2610 -7014 -2608
rect -6812 -2610 -6767 -2608
rect -6698 -2610 -6664 -2608
rect -6582 -2610 -6548 -2608
rect -12120 -2676 -6514 -2610
rect -6468 -2676 -6434 -2608
rect -12120 -2710 -6304 -2676
rect -12120 -2902 -6514 -2710
rect -6468 -2902 -6434 -2710
rect -12120 -2988 -6434 -2902
rect -12120 -3001 -6514 -2988
rect -28336 -3012 -6514 -3001
rect -28336 -3048 -17291 -3012
rect -28336 -3071 -18484 -3048
rect -28336 -3380 -23708 -3071
rect -29156 -3884 -28712 -3808
rect -28939 -4026 -28894 -3884
rect -28939 -5494 -28905 -4026
rect -28862 -5547 -28834 -3884
rect -28806 -5547 -28778 -3884
rect -28757 -4026 -28712 -3884
rect -28757 -5494 -28723 -4026
rect -28336 -4568 -23715 -3380
rect -28336 -4871 -23708 -4568
rect -28336 -5553 -27439 -4871
rect -29853 -5587 -27439 -5553
rect -30625 -5655 -30591 -5621
rect -29967 -5655 -29933 -5621
rect -29853 -5655 -29819 -5587
rect -29532 -5600 -29504 -5593
rect -29476 -5600 -29448 -5593
rect -28862 -5600 -28834 -5593
rect -28806 -5600 -28778 -5593
rect -28336 -5655 -27439 -5587
rect -31503 -5689 -27439 -5655
rect -31941 -5844 -31907 -5810
rect -32608 -5878 -32218 -5844
rect -32608 -5906 -32574 -5878
rect -32608 -6314 -32540 -5906
rect -32394 -5946 -32347 -5899
rect -32432 -5980 -32347 -5946
rect -32505 -6039 -32460 -6028
rect -32377 -6039 -32332 -6028
rect -32494 -6215 -32460 -6039
rect -32366 -6215 -32332 -6039
rect -32394 -6274 -32347 -6227
rect -32432 -6308 -32347 -6274
rect -32608 -6376 -32574 -6314
rect -32252 -6376 -32218 -5878
rect -32608 -6410 -32218 -6376
rect -32132 -5878 -31742 -5844
rect -32132 -6376 -32098 -5878
rect -31941 -5912 -31894 -5899
rect -31941 -5924 -31884 -5912
rect -31962 -5980 -31884 -5924
rect -32052 -6032 -32034 -5999
rect -31962 -6023 -31888 -5980
rect -31962 -6027 -31873 -6023
rect -32024 -6028 -32006 -6027
rect -31962 -6028 -31860 -6027
rect -32029 -6039 -31984 -6028
rect -32018 -6215 -31984 -6039
rect -31962 -6034 -31856 -6028
rect -31962 -6038 -31850 -6034
rect -31962 -6215 -31856 -6038
rect -31962 -6218 -31860 -6215
rect -31962 -6227 -31850 -6218
rect -32010 -6228 -31984 -6227
rect -31982 -6231 -31873 -6227
rect -31982 -6240 -31888 -6231
rect -31982 -6256 -31884 -6240
rect -31962 -6284 -31884 -6256
rect -31982 -6308 -31884 -6284
rect -31982 -6348 -31888 -6308
rect -31998 -6362 -31982 -6360
rect -31962 -6376 -31888 -6348
rect -31876 -6376 -31874 -6231
rect -31776 -6376 -31742 -5878
rect -32132 -6410 -31742 -6376
rect -31962 -6460 -31888 -6410
rect -33291 -7044 -33268 -6970
rect -33263 -7072 -33240 -6970
rect -32626 -7080 -32204 -6460
rect -32150 -7080 -31728 -6460
rect -33291 -7334 -33268 -7212
rect -33263 -7306 -33240 -7184
rect -29853 -7393 -29819 -5689
rect -28336 -5725 -27439 -5689
rect -27339 -5180 -23708 -4871
rect -23686 -4968 -23641 -3071
rect -23210 -4968 -23165 -3071
rect -23140 -3380 -23112 -3071
rect -23110 -3112 -18484 -3071
rect -23110 -3250 -18534 -3112
rect -18518 -3180 -18484 -3112
rect -18418 -3180 -17291 -3048
rect -18518 -3214 -17291 -3180
rect -23084 -3380 -23056 -3250
rect -23028 -3300 -22983 -3250
rect -22914 -3300 -22880 -3250
rect -22783 -3300 -18534 -3250
rect -18418 -3264 -17291 -3214
rect -23052 -3334 -18534 -3300
rect -23052 -3814 -22983 -3334
rect -22914 -3364 -22880 -3334
rect -22914 -3436 -22822 -3364
rect -22914 -3475 -22880 -3436
rect -22783 -3464 -18534 -3334
rect -18532 -3464 -17291 -3264
rect -22949 -3486 -22880 -3475
rect -22861 -3486 -22805 -3475
rect -22938 -3662 -22880 -3486
rect -22850 -3662 -22805 -3486
rect -22783 -3514 -17291 -3464
rect -17214 -3035 -6514 -3012
rect -17214 -3071 -12220 -3035
rect -17214 -3492 -13567 -3071
rect -17224 -3500 -13567 -3492
rect -22783 -3524 -18534 -3514
rect -18532 -3524 -17291 -3514
rect -22783 -3606 -17291 -3524
rect -22914 -3674 -22880 -3662
rect -22914 -3746 -22822 -3674
rect -22914 -3814 -22880 -3746
rect -22783 -3814 -18534 -3606
rect -23052 -3848 -18534 -3814
rect -27339 -5530 -23715 -5180
rect -23686 -5480 -23652 -4968
rect -23210 -5480 -23176 -4968
rect -23140 -5180 -23112 -4568
rect -23084 -5180 -23056 -4568
rect -23028 -4968 -22983 -3848
rect -23028 -5480 -22994 -4968
rect -22914 -5530 -22880 -3848
rect -22783 -3853 -18534 -3848
rect -18532 -3853 -17291 -3606
rect -22783 -3884 -17291 -3853
rect -22783 -3934 -18472 -3884
rect -22783 -4002 -18516 -3934
rect -18500 -3968 -18472 -3934
rect -18500 -4002 -18482 -3968
rect -18418 -4002 -17291 -3884
rect -22783 -4036 -17291 -4002
rect -22783 -4086 -18534 -4036
rect -18418 -4086 -17291 -4036
rect -22783 -4558 -17291 -4086
rect -17214 -4288 -13567 -3500
rect -13308 -4288 -13263 -3071
rect -13062 -4032 -13017 -3071
rect -12650 -3480 -12605 -3071
rect -12684 -3622 -12658 -3480
rect -12650 -3622 -12616 -3480
rect -13100 -4146 -12908 -4032
rect -12650 -4134 -12605 -3622
rect -13080 -4288 -13006 -4146
rect -17214 -4356 -12802 -4288
rect -17214 -4514 -13274 -4356
rect -22783 -4706 -18332 -4558
rect -18278 -4706 -17856 -4558
rect -17802 -4706 -17291 -4558
rect -22783 -4848 -18644 -4706
rect -22783 -4856 -22368 -4848
rect -22268 -4856 -18644 -4848
rect -22783 -4890 -18644 -4856
rect -22783 -4940 -22368 -4890
rect -22268 -4940 -18644 -4890
rect -18226 -4904 -18210 -4706
rect -18154 -4724 -18008 -4706
rect -18154 -4788 -18061 -4724
rect -18154 -4798 -18080 -4788
rect -18132 -4826 -18099 -4798
rect -22783 -5530 -18644 -4940
rect -27339 -5564 -18644 -5530
rect -27339 -5632 -23715 -5564
rect -22914 -5580 -22880 -5564
rect -22914 -5591 -22903 -5580
rect -22891 -5591 -22880 -5580
rect -22783 -5570 -18644 -5564
rect -17712 -5530 -17291 -4706
rect -17191 -4871 -13274 -4514
rect -16904 -5492 -16870 -4871
rect -16280 -5492 -16248 -4871
rect -16246 -5492 -16212 -4871
rect -17260 -5530 -16212 -5492
rect -16054 -5492 -16020 -4871
rect -15940 -5492 -15906 -4871
rect -15808 -5492 -15774 -4871
rect -15694 -5480 -15660 -4871
rect -15588 -5492 -15554 -4871
rect -16054 -5530 -16016 -5492
rect -15940 -5530 -15902 -5492
rect -15808 -5530 -15770 -5492
rect -15588 -5530 -15550 -5492
rect -15282 -5530 -15248 -4871
rect -15036 -5480 -15002 -4871
rect -14930 -5492 -14896 -4871
rect -14930 -5530 -14892 -5492
rect -14624 -5530 -14590 -4871
rect -14378 -5480 -14344 -4871
rect -14272 -5492 -14238 -4871
rect -14272 -5530 -14234 -5492
rect -14158 -5530 -14124 -4871
rect -13966 -5484 -13932 -4871
rect -13740 -4926 -13274 -4871
rect -13264 -4926 -12802 -4356
rect -13720 -4976 -13686 -4926
rect -13720 -5010 -13336 -4976
rect -13720 -5480 -13652 -5010
rect -13494 -5078 -13456 -5040
rect -13528 -5112 -13456 -5078
rect -13583 -5162 -13538 -5151
rect -13495 -5162 -13450 -5151
rect -13572 -5338 -13538 -5162
rect -13484 -5338 -13450 -5162
rect -13494 -5388 -13456 -5350
rect -13528 -5422 -13456 -5388
rect -13966 -5492 -13921 -5484
rect -13686 -5490 -13652 -5480
rect -13370 -5490 -13336 -5010
rect -13686 -5492 -13336 -5490
rect -13308 -5484 -13274 -4926
rect -13062 -4976 -13028 -4926
rect -13210 -5010 -12860 -4976
rect -13308 -5492 -13263 -5484
rect -13210 -5490 -13176 -5010
rect -13062 -5044 -13028 -5010
rect -13086 -5078 -13028 -5044
rect -13018 -5078 -12980 -5040
rect -13062 -5112 -12980 -5078
rect -13062 -5151 -13028 -5112
rect -13008 -5151 -12994 -5146
rect -13107 -5162 -13028 -5151
rect -13019 -5162 -12974 -5151
rect -13096 -5338 -13028 -5162
rect -13062 -5354 -13028 -5338
rect -13008 -5338 -12974 -5162
rect -13008 -5350 -12994 -5338
rect -13086 -5388 -13028 -5354
rect -13018 -5388 -12980 -5350
rect -13062 -5422 -12980 -5388
rect -13062 -5480 -13028 -5422
rect -12894 -5490 -12860 -5010
rect -13210 -5492 -12860 -5490
rect -12650 -5492 -12616 -4134
rect -14070 -5530 -13710 -5492
rect -13696 -5524 -12856 -5492
rect -13696 -5530 -13052 -5524
rect -13038 -5530 -12856 -5524
rect -12662 -5530 -12604 -5492
rect -17712 -5564 -16870 -5530
rect -16842 -5564 -16212 -5530
rect -16200 -5564 -13710 -5530
rect -13658 -5564 -13052 -5530
rect -13000 -5564 -12604 -5530
rect -22783 -5587 -18618 -5570
rect -22783 -5632 -22368 -5587
rect -27339 -5655 -22368 -5632
rect -22268 -5655 -18644 -5587
rect -27339 -5666 -18644 -5655
rect -27339 -5702 -23715 -5666
rect -22783 -5689 -18644 -5666
rect -22783 -5702 -22368 -5689
rect -27339 -7353 -24712 -5702
rect -24595 -6114 -24574 -6032
rect -24557 -6152 -24536 -5994
rect -23906 -6124 -23853 -6070
rect -23785 -6124 -23751 -5702
rect -22268 -5725 -18644 -5689
rect -17712 -5632 -17291 -5564
rect -16904 -5632 -16870 -5564
rect -16280 -5628 -16248 -5564
rect -16246 -5632 -16212 -5564
rect -16054 -5632 -16020 -5564
rect -15940 -5628 -15906 -5564
rect -15940 -5632 -15895 -5628
rect -15808 -5632 -15774 -5564
rect -15588 -5628 -15554 -5564
rect -15282 -5628 -15248 -5564
rect -14930 -5628 -14896 -5564
rect -14624 -5628 -14590 -5564
rect -14272 -5628 -14238 -5564
rect -15588 -5632 -15543 -5628
rect -15282 -5632 -15237 -5628
rect -14930 -5632 -14885 -5628
rect -14624 -5632 -14579 -5628
rect -14272 -5632 -14227 -5628
rect -14158 -5632 -14124 -5564
rect -13978 -5580 -13920 -5564
rect -13320 -5580 -13262 -5564
rect -12662 -5580 -12604 -5564
rect -12619 -5595 -12604 -5580
rect -12536 -5632 -12502 -3071
rect -12398 -3622 -12370 -3480
rect -12364 -3622 -12336 -3480
rect -12182 -3554 -12148 -3035
rect -12120 -3306 -6514 -3035
rect -12120 -3632 -8594 -3306
rect -8566 -3480 -8522 -3306
rect -8566 -3632 -8532 -3480
rect -8494 -3564 -8485 -3530
rect -8358 -3632 -8324 -3306
rect -8244 -3492 -8199 -3306
rect -7898 -3378 -7853 -3306
rect -7924 -3434 -7853 -3378
rect -7586 -3434 -7541 -3306
rect -7472 -3434 -7438 -3306
rect -7240 -3434 -7206 -3306
rect -8148 -3492 -7686 -3434
rect -7672 -3480 -7206 -3434
rect -7672 -3492 -7210 -3480
rect -8256 -3564 -7210 -3492
rect -8256 -3580 -8198 -3564
rect -8256 -3595 -8210 -3580
rect -8244 -3632 -8210 -3595
rect -8148 -3632 -7686 -3564
rect -7672 -3632 -7210 -3564
rect -7048 -3632 -7014 -3306
rect -6934 -3492 -6889 -3306
rect -6602 -3410 -6514 -3306
rect -6654 -3486 -6504 -3410
rect -6946 -3552 -6572 -3492
rect -6996 -3564 -6572 -3552
rect -6996 -3570 -6888 -3564
rect -6946 -3580 -6888 -3570
rect -6946 -3595 -6931 -3580
rect -6996 -3626 -6940 -3608
rect -6934 -3632 -6900 -3598
rect -6894 -3626 -6840 -3608
rect -6468 -3632 -6434 -2988
rect -6282 -3544 -6272 -2748
rect -6251 -2870 -6230 -2748
rect -6226 -2836 -6192 -2608
rect -6162 -2836 -6128 -2608
rect -6124 -2696 -6074 -2522
rect -5926 -2556 -5920 -2392
rect -5910 -2418 -5900 -2392
rect -5910 -2662 -5876 -2418
rect -5750 -2566 -5716 -2418
rect -5636 -2566 -5602 -2532
rect -5548 -2566 -5514 -2532
rect -5434 -2566 -5400 -2418
rect -5784 -2600 -5056 -2566
rect -5910 -2774 -5846 -2662
rect -6226 -2870 -6176 -2836
rect -6162 -2870 -5972 -2836
rect -6282 -3570 -6280 -3544
rect -12120 -3666 -6434 -3632
rect -12120 -3686 -8594 -3666
rect -11312 -4288 -11278 -3686
rect -9548 -3896 -9514 -3686
rect -9434 -3744 -9389 -3686
rect -9356 -3756 -9282 -3686
rect -8776 -3744 -8731 -3686
rect -9410 -3794 -8766 -3756
rect -9372 -3828 -8766 -3794
rect -9356 -3896 -9282 -3828
rect -8662 -3834 -8612 -3686
rect -8662 -3896 -8634 -3834
rect -9548 -3930 -8634 -3896
rect -9356 -3944 -9282 -3930
rect -12390 -4708 -12364 -4568
rect -11872 -4716 -11410 -4288
rect -11396 -4716 -10934 -4288
rect -9316 -4436 -9304 -4088
rect -9278 -4398 -9266 -4126
rect -11872 -4722 -10934 -4716
rect -12212 -4924 -12196 -4822
rect -11872 -4848 -11410 -4722
rect -11396 -4848 -10934 -4722
rect -8600 -4774 -8590 -4134
rect -8566 -4716 -8532 -3666
rect -8358 -3834 -8324 -3666
rect -8244 -3744 -8210 -3666
rect -8148 -3794 -7686 -3666
rect -7672 -3702 -7210 -3666
rect -7672 -3794 -7402 -3702
rect -8148 -3828 -7402 -3794
rect -8148 -3966 -7686 -3828
rect -7672 -3966 -7402 -3828
rect -7672 -4072 -7432 -3966
rect -8094 -4368 -7712 -4130
rect -7980 -4484 -7946 -4368
rect -7892 -4484 -7858 -4368
rect -7048 -4426 -7014 -3666
rect -6940 -3926 -6930 -3818
rect -6162 -4426 -6128 -2870
rect -5880 -4418 -5846 -2774
rect -5750 -2836 -5716 -2600
rect -5648 -2696 -5502 -2630
rect -5630 -2702 -5520 -2696
rect -5592 -2740 -5558 -2734
rect -5592 -2768 -5520 -2740
rect -5434 -2794 -5400 -2600
rect -5434 -2814 -5178 -2794
rect -5434 -2836 -5400 -2814
rect -5750 -2870 -5400 -2836
rect -5382 -2999 -5381 -2814
rect -5198 -2999 -5178 -2814
rect -5382 -3000 -5178 -2999
rect -8566 -4774 -8556 -4716
rect -12184 -4924 -12168 -4850
rect -11708 -4870 -11554 -4850
rect -11396 -4868 -11156 -4848
rect -11396 -4870 -11078 -4868
rect -11396 -4926 -11156 -4870
rect -12196 -5124 -12020 -5098
rect -11664 -5120 -11622 -5098
rect -7132 -5138 -7108 -4444
rect -7098 -5138 -7074 -4478
rect -12390 -5180 -12364 -5154
rect -11146 -5162 -11132 -5154
rect -11228 -5338 -11194 -5162
rect -11146 -5180 -11106 -5162
rect -11140 -5338 -11106 -5180
rect -17712 -5666 -12352 -5632
rect -17712 -5725 -17291 -5666
rect -24328 -6158 -23938 -6124
rect -24328 -6656 -24294 -6158
rect -24199 -6226 -24067 -6179
rect -24152 -6260 -24067 -6226
rect -24225 -6319 -24169 -6308
rect -24097 -6319 -24041 -6308
rect -24214 -6495 -24169 -6319
rect -24086 -6495 -24041 -6319
rect -24199 -6520 -24067 -6507
rect -24199 -6540 -24064 -6520
rect -24199 -6554 -24067 -6540
rect -24152 -6588 -24067 -6554
rect -23972 -6656 -23938 -6158
rect -23877 -6186 -23853 -6124
rect -23886 -6220 -23853 -6186
rect -23877 -6540 -23853 -6220
rect -24328 -6690 -23938 -6656
rect -23886 -6690 -23853 -6540
rect -23852 -6158 -23799 -6124
rect -23785 -6158 -23558 -6124
rect -23852 -6656 -23818 -6158
rect -23785 -6656 -23751 -6158
rect -23750 -6507 -23697 -6307
rect -23726 -6540 -23588 -6520
rect -23692 -6574 -23622 -6554
rect -23852 -6690 -23799 -6656
rect -23785 -6690 -23558 -6656
rect -23886 -6722 -23865 -6690
rect -23888 -6740 -23853 -6722
rect -23785 -6740 -23751 -6690
rect -24346 -7353 -23924 -6740
rect -23888 -6776 -23715 -6740
rect -27466 -7356 -24585 -7353
rect -27466 -7364 -24552 -7356
rect -27339 -7387 -24552 -7364
rect -24495 -7360 -23924 -7353
rect -23870 -6950 -23715 -6776
rect -23870 -7150 -23697 -6950
rect -23870 -7360 -23715 -7150
rect -24495 -7387 -23927 -7360
rect -27339 -7502 -24712 -7387
rect -23785 -7393 -23751 -7360
rect -22268 -7502 -19159 -5725
rect -18748 -6066 -18726 -5725
rect -18714 -6066 -18692 -5725
rect -17820 -6726 -17358 -6088
rect -17676 -6776 -17642 -6726
rect -17562 -6776 -17528 -6742
rect -17676 -6810 -17416 -6776
rect -17676 -6962 -17642 -6810
rect -17562 -6840 -17528 -6810
rect -17574 -6878 -17528 -6840
rect -17624 -6912 -17528 -6878
rect -17574 -6950 -17528 -6912
rect -17562 -6962 -17528 -6950
rect -17664 -7138 -17642 -6962
rect -17564 -7138 -17528 -6962
rect -17954 -7502 -17944 -7222
rect -17926 -7530 -17916 -7222
rect -17676 -7290 -17642 -7138
rect -17562 -7150 -17528 -7138
rect -17574 -7188 -17528 -7150
rect -17624 -7222 -17528 -7188
rect -17574 -7253 -17528 -7222
rect -17562 -7280 -17528 -7253
rect -17450 -7290 -17416 -6810
rect -16904 -7280 -16870 -5666
rect -16054 -6076 -16020 -5666
rect -15940 -5924 -15895 -5666
rect -15588 -5936 -15543 -5666
rect -15282 -5924 -15237 -5666
rect -14930 -5936 -14885 -5666
rect -14624 -5924 -14579 -5666
rect -14272 -5936 -14227 -5666
rect -15916 -5974 -15272 -5936
rect -15258 -5974 -14614 -5936
rect -14600 -5974 -14226 -5936
rect -15878 -6008 -15272 -5974
rect -15220 -6008 -14614 -5974
rect -14562 -6008 -14226 -5974
rect -15600 -6024 -15542 -6008
rect -14942 -6024 -14884 -6008
rect -14284 -6024 -14226 -6008
rect -15588 -6076 -15554 -6042
rect -14930 -6076 -14896 -6024
rect -14272 -6039 -14226 -6024
rect -14272 -6076 -14238 -6039
rect -14158 -6076 -14124 -5666
rect -13966 -5696 -13932 -5666
rect -14074 -6008 -13994 -5994
rect -13598 -6008 -13436 -5994
rect -12536 -6014 -12502 -5666
rect -4720 -6014 -4686 -1582
rect -4606 -1708 -4572 -1582
rect -4606 -2562 -4566 -1708
rect -3296 -2562 -3272 -1242
rect -2960 -1584 -2926 -1242
rect -2858 -1464 -2824 -1242
rect -2632 -1470 -2598 -1242
rect -1974 -1470 -1940 -892
rect -1316 -1470 -1282 -868
rect -1202 -1470 -1168 -868
rect -884 -960 2740 -868
rect 3100 -954 3134 -868
rect 3214 -954 3248 -868
rect 3252 -938 3254 -874
rect 3283 -954 6907 -868
rect -884 -1470 2848 -960
rect 3100 -1470 6907 -954
rect -2896 -1554 -2824 -1516
rect -2774 -1526 6907 -1470
rect -2645 -1538 -2644 -1537
rect -2644 -1539 -2643 -1538
rect -2858 -1580 -2824 -1554
rect -2896 -1584 -2824 -1580
rect -2632 -1584 -2598 -1526
rect -2586 -1538 -2585 -1537
rect -1987 -1538 -1986 -1537
rect -2587 -1539 -2586 -1538
rect -1986 -1539 -1985 -1538
rect -1974 -1584 -1940 -1526
rect -1928 -1538 -1927 -1537
rect -1329 -1538 -1328 -1537
rect -1929 -1539 -1928 -1538
rect -1328 -1539 -1327 -1538
rect -1316 -1584 -1282 -1526
rect -1202 -1584 -1168 -1526
rect -884 -1584 2848 -1526
rect 3100 -1584 6907 -1526
rect -2960 -1618 6907 -1584
rect -2960 -1728 -2926 -1618
rect -2858 -1672 -2824 -1618
rect -2858 -1728 -2786 -1672
rect -2960 -1814 -2786 -1728
rect -2960 -2212 -2926 -1814
rect -2858 -2056 -2786 -1814
rect -2632 -2056 -2598 -1618
rect -1974 -2002 -1940 -1618
rect -2858 -2090 -2270 -2056
rect -2858 -2122 -2784 -2090
rect -2818 -2174 -2784 -2122
rect -2644 -2138 -2643 -2137
rect -2645 -2139 -2644 -2138
rect -2632 -2150 -2598 -2090
rect -2304 -2118 -2270 -2090
rect -2587 -2138 -2586 -2137
rect -2586 -2139 -2585 -2138
rect -2338 -2150 -2236 -2118
rect -2220 -2132 -1582 -2002
rect -1376 -2066 -1322 -2052
rect -1322 -2108 -1320 -2066
rect -2220 -2139 -1430 -2132
rect -1328 -2138 -1327 -2137
rect -1329 -2139 -1328 -2138
rect -2220 -2150 -1428 -2139
rect -1316 -2150 -1282 -1618
rect -1202 -2150 -1168 -1618
rect -2896 -2212 -2784 -2174
rect -2774 -2184 -1168 -2150
rect -2960 -2290 -2784 -2212
rect -2754 -2214 -2682 -2184
rect -2645 -2196 -2644 -2195
rect -2644 -2197 -2643 -2196
rect -2716 -2248 -2682 -2214
rect -2632 -2204 -2445 -2184
rect -2960 -2562 -2926 -2290
rect -2858 -2372 -2784 -2290
rect -2632 -2258 -2598 -2204
rect -2444 -2214 -2372 -2184
rect -2456 -2258 -2445 -2247
rect -2406 -2248 -2372 -2214
rect -2632 -2292 -2445 -2258
rect -2632 -2372 -2598 -2292
rect -2304 -2372 -2270 -2184
rect -2858 -2406 -2270 -2372
rect -2220 -2206 -1430 -2184
rect -1329 -2196 -1328 -2195
rect -1328 -2197 -1327 -2196
rect -2858 -2532 -2786 -2406
rect -2632 -2532 -2598 -2406
rect -2220 -2464 -1582 -2206
rect -1322 -2276 -1320 -2216
rect -1974 -2478 -1940 -2464
rect -2858 -2558 -2270 -2532
rect -2896 -2562 -2270 -2558
rect -2220 -2562 -1582 -2478
rect -1316 -2562 -1282 -2184
rect -1202 -2562 -1168 -2184
rect -4618 -2596 -1168 -2562
rect -4606 -2602 -4566 -2596
rect -4612 -2658 -4566 -2602
rect -3948 -2626 -3914 -2596
rect -3296 -2602 -3256 -2596
rect -3296 -2626 -3250 -2602
rect -2960 -2626 -2926 -2596
rect -2858 -2626 -2784 -2596
rect -2632 -2626 -2598 -2596
rect -2304 -2626 -2270 -2596
rect -2220 -2626 -1582 -2596
rect -1316 -2626 -1282 -2596
rect -4606 -2704 -4566 -2658
rect -4556 -2664 -4538 -2658
rect -3976 -2664 -3914 -2626
rect -3834 -2664 -2778 -2626
rect -2660 -2630 -2598 -2626
rect -2494 -2630 -2440 -2626
rect -2660 -2646 -2440 -2630
rect -2678 -2664 -2440 -2646
rect -2304 -2664 -2266 -2626
rect -2220 -2664 -1428 -2626
rect -1344 -2664 -1282 -2626
rect -4560 -2698 -3914 -2664
rect -3902 -2698 -3250 -2664
rect -4556 -2704 -4538 -2698
rect -4612 -2742 -4566 -2704
rect -4606 -2802 -4540 -2742
rect -4516 -2802 -4512 -2714
rect -4606 -3002 -4572 -2802
rect -4606 -3148 -4540 -3002
rect -4606 -3258 -4566 -3148
rect -4516 -3176 -4512 -3002
rect -4612 -3314 -4566 -3258
rect -3948 -3282 -3914 -2698
rect -3324 -2704 -3306 -2698
rect -3296 -2760 -3250 -2698
rect -3240 -2680 -1282 -2664
rect -3240 -2698 -2598 -2680
rect -2586 -2698 -1282 -2680
rect -3240 -2704 -3222 -2698
rect -3290 -3088 -3256 -2760
rect -3296 -3258 -3256 -3088
rect -3296 -3282 -3250 -3258
rect -2960 -3282 -2926 -2698
rect -2858 -2780 -2784 -2698
rect -2716 -2724 -2682 -2698
rect -2672 -2724 -2638 -2700
rect -2644 -2774 -2638 -2728
rect -2632 -2734 -2598 -2698
rect -2592 -2724 -2538 -2700
rect -2592 -2734 -2538 -2728
rect -2456 -2734 -2445 -2723
rect -2406 -2724 -2372 -2698
rect -2632 -2768 -2445 -2734
rect -2818 -2832 -2784 -2780
rect -2644 -2796 -2643 -2795
rect -2645 -2797 -2644 -2796
rect -2632 -2808 -2598 -2768
rect -2592 -2780 -2538 -2768
rect -2587 -2796 -2586 -2795
rect -2586 -2797 -2585 -2796
rect -2304 -2808 -2270 -2698
rect -2220 -2797 -1582 -2698
rect -1328 -2796 -1327 -2795
rect -1329 -2797 -1328 -2796
rect -2220 -2808 -1428 -2797
rect -1322 -2802 -1320 -2750
rect -1316 -2808 -1282 -2698
rect -1202 -2808 -1168 -2596
rect -2774 -2814 -1168 -2808
rect -2896 -2848 -2784 -2832
rect -2778 -2842 -1168 -2814
rect -2632 -2848 -2598 -2842
rect -2304 -2848 -2270 -2842
rect -2896 -2870 -2270 -2848
rect -2858 -2882 -2270 -2870
rect -2858 -2886 -2786 -2882
rect -4606 -3360 -4566 -3314
rect -4556 -3320 -4538 -3314
rect -3976 -3320 -3914 -3282
rect -3834 -3320 -2922 -3282
rect -2858 -3320 -2824 -2886
rect -2632 -3282 -2598 -2882
rect -2220 -2940 -1582 -2842
rect -1329 -2854 -1328 -2853
rect -1328 -2855 -1327 -2854
rect -1322 -2940 -1320 -2848
rect -1974 -3282 -1940 -2940
rect -1316 -3282 -1282 -2842
rect -2660 -3320 -2598 -3282
rect -2002 -3320 -1940 -3282
rect -1344 -3320 -1282 -3282
rect -4560 -3354 -3914 -3320
rect -3902 -3354 -3250 -3320
rect -4556 -3360 -4538 -3354
rect -4612 -3416 -4566 -3360
rect -4606 -3422 -4566 -3416
rect -3948 -3422 -3914 -3354
rect -3324 -3360 -3306 -3354
rect -3296 -3416 -3250 -3354
rect -3240 -3354 -2598 -3320
rect -2586 -3354 -1940 -3320
rect -1928 -3354 -1282 -3320
rect -3240 -3360 -3222 -3354
rect -3296 -3422 -3256 -3416
rect -2960 -3422 -2926 -3354
rect -2858 -3412 -2824 -3354
rect -2632 -3412 -2598 -3354
rect -1974 -3412 -1940 -3354
rect -1316 -3412 -1282 -3354
rect -2858 -3422 -2786 -3412
rect -2632 -3422 -2587 -3412
rect -1974 -3422 -1929 -3412
rect -1316 -3422 -1271 -3412
rect -1202 -3422 -1168 -2842
rect -4624 -3456 -1168 -3422
rect -4572 -4252 -4566 -3456
rect -3894 -3924 -3850 -3908
rect -3860 -3950 -3850 -3942
rect -3888 -4196 -3874 -3950
rect -3860 -4252 -3818 -3950
rect -3296 -3996 -3272 -3456
rect -2960 -4238 -2926 -3456
rect -2785 -3466 -2644 -3456
rect -2632 -3466 -2598 -3456
rect -2586 -3466 -1986 -3456
rect -1974 -3466 -1940 -3456
rect -1928 -3466 -1328 -3456
rect -1316 -3466 -1282 -3456
rect -1202 -3466 -1168 -3456
rect -884 -2398 2848 -1618
rect 3100 -1756 6907 -1618
rect 3064 -1766 6907 -1756
rect 3100 -1868 6907 -1766
rect 3118 -2392 6907 -1868
rect -884 -2808 2740 -2398
rect 3283 -2562 6907 -2392
rect 7516 -2562 7550 -688
rect 7570 -1154 7604 -688
rect 7690 -748 7800 -710
rect 7728 -782 7800 -748
rect 7673 -832 7729 -821
rect 7761 -832 7817 -821
rect 7684 -1008 7729 -832
rect 7772 -1008 7817 -832
rect 7690 -1058 7800 -1020
rect 7728 -1092 7800 -1058
rect 7566 -1160 7604 -1154
rect 7886 -1160 7920 -688
rect 8082 -824 8108 -720
rect 8138 -824 8164 -720
rect 7566 -1194 7920 -1160
rect 7566 -1372 7584 -1194
rect 8082 -2176 8108 -1372
rect 8138 -2176 8164 -1372
rect 8174 -2176 8208 -688
rect 8390 -2176 8424 -688
rect 8504 -2176 8549 -688
rect 8832 -1312 8866 -94
rect 8946 -1312 8980 58
rect 9118 -822 9140 52
rect 9162 -1124 9196 712
rect 9264 646 12896 746
rect 9264 600 12988 646
rect 13288 610 13298 1084
rect 13431 877 14102 1084
rect 14118 877 14146 1120
rect 14174 877 14202 1120
rect 14239 877 17531 1120
rect 13431 843 17531 877
rect 13431 822 14102 843
rect 14118 822 14146 843
rect 13431 809 14146 822
rect 14174 822 14202 843
rect 14239 822 17531 843
rect 17674 840 17698 1946
rect 14174 818 17531 822
rect 14174 809 17686 818
rect 13431 741 17686 809
rect 13431 740 14102 741
rect 13431 735 14174 740
rect 13431 725 14146 735
rect 14174 725 14202 735
rect 14239 725 17686 741
rect 13431 678 17686 725
rect 13431 610 14146 678
rect 14150 644 17686 678
rect 14150 638 14202 644
rect 13080 600 14146 610
rect 9264 590 12896 600
rect 9264 572 12932 590
rect 13288 582 13298 600
rect 13431 594 14146 600
rect 14174 594 14202 638
rect 13431 582 14164 594
rect 13108 572 14164 582
rect 9264 320 12896 572
rect 13288 436 13298 572
rect 13288 320 13316 436
rect 13431 354 14164 572
rect 14174 354 14192 594
rect 9232 -972 9254 132
rect 9264 14 12932 320
rect 9264 -440 11988 14
rect 11996 -168 12044 14
rect 12046 -168 12080 14
rect 12562 -168 12596 14
rect 12624 -168 12638 14
rect 12652 -168 12694 14
rect 12704 -168 12738 14
rect 12818 -80 12852 14
rect 13108 6 13404 320
rect 13431 6 14146 354
rect 14174 298 14220 354
rect 14174 82 14202 298
rect 14239 174 17686 644
rect 17702 212 17704 2158
rect 17708 806 17732 1980
rect 17708 208 17742 230
rect 17698 174 17776 196
rect 14239 140 17696 174
rect 12768 -108 12988 -80
rect 12768 -126 12888 -108
rect 12768 -142 12944 -126
rect 12818 -168 12852 -142
rect 12888 -144 12944 -142
rect 13334 -168 13368 0
rect 13431 -132 13658 6
rect 13467 -168 13501 -132
rect 13943 -168 13977 6
rect 13986 -168 14020 6
rect 14057 -168 14091 6
rect 14100 -168 14146 6
rect 14239 60 17686 140
rect 17698 106 17730 174
rect 17822 134 17856 5886
rect 19263 5850 22887 5886
rect 23550 5870 23584 5886
rect 23866 5870 23900 5886
rect 19299 3780 19333 5850
rect 18272 3746 21728 3780
rect 18176 296 18210 3684
rect 18256 3542 18276 3635
rect 18290 3508 18310 3601
rect 18948 3597 18982 3601
rect 18942 3572 18982 3597
rect 18984 3572 18988 3597
rect 19299 3572 19333 3746
rect 19413 3709 19460 3725
rect 19401 3678 19460 3709
rect 19578 3678 19625 3725
rect 20071 3694 20118 3725
rect 20059 3678 20118 3694
rect 20236 3678 20283 3725
rect 20729 3694 20776 3725
rect 20717 3678 20776 3694
rect 20894 3678 20941 3725
rect 21387 3694 21434 3725
rect 21375 3678 21434 3694
rect 21552 3678 21599 3725
rect 19401 3644 19625 3678
rect 19668 3644 20283 3678
rect 20326 3644 20941 3678
rect 20984 3644 21599 3678
rect 19401 3597 19459 3644
rect 19413 3572 19447 3597
rect 19606 3596 19640 3601
rect 20059 3597 20117 3644
rect 19595 3585 19640 3596
rect 19606 3572 19640 3585
rect 20071 3572 20105 3597
rect 20264 3596 20298 3601
rect 20717 3597 20775 3644
rect 20253 3585 20298 3596
rect 20264 3572 20298 3585
rect 20729 3572 20763 3597
rect 20922 3596 20956 3601
rect 21375 3597 21433 3644
rect 20911 3585 20956 3596
rect 20922 3572 20956 3585
rect 21387 3572 21421 3597
rect 21492 3572 21514 3638
rect 21520 3596 21570 3638
rect 21580 3596 21614 3601
rect 21520 3585 21614 3596
rect 21520 3572 21570 3585
rect 21580 3572 21614 3585
rect 21694 3572 21728 3746
rect 18502 2097 22602 3572
rect 24370 3567 24404 5886
rect 26458 3567 26492 5886
rect 27888 3567 27922 5886
rect 31220 4242 31254 7100
rect 41946 7062 41980 8936
rect 42734 8826 42738 8936
rect 43614 8934 45264 10372
rect 45718 10370 49342 10374
rect 49885 10370 53509 10385
rect 54712 10372 54738 10664
rect 54740 10372 54794 10664
rect 54854 10636 54878 10738
rect 54882 10704 54906 10710
rect 56078 10704 56112 10772
rect 56180 10704 56358 10742
rect 56372 10704 56896 10742
rect 54882 10670 55562 10704
rect 55652 10670 56358 10704
rect 56410 10670 56896 10704
rect 54882 10664 54906 10670
rect 55590 10504 55624 10620
rect 56078 10504 56112 10670
rect 56180 10632 56238 10670
rect 56838 10632 56896 10670
rect 56192 10504 56237 10632
rect 56337 10620 56393 10631
rect 56348 10504 56393 10620
rect 56850 10504 56895 10632
rect 56964 10504 56998 10772
rect 57268 10504 57302 10772
rect 57370 10670 57874 10742
rect 57978 10710 58012 10772
rect 57370 10632 57428 10670
rect 57382 10504 57427 10632
rect 57853 10620 57909 10631
rect 57864 10504 57909 10620
rect 57978 10520 58030 10710
rect 58040 10538 58046 10744
rect 57978 10504 58012 10520
rect 58040 10504 58074 10538
rect 58154 10504 58188 10932
rect 54992 10470 58448 10504
rect 54992 10372 55026 10470
rect 55590 10440 55624 10470
rect 55722 10440 55742 10470
rect 56078 10440 56112 10470
rect 56192 10440 56237 10470
rect 56348 10440 56393 10470
rect 56850 10440 56895 10470
rect 56964 10440 56998 10470
rect 57268 10440 57302 10470
rect 57382 10440 57427 10470
rect 57864 10440 57909 10470
rect 57978 10440 58012 10470
rect 58040 10440 58046 10470
rect 55130 10402 55774 10440
rect 55788 10402 56432 10440
rect 56446 10402 57090 10440
rect 57104 10402 57748 10440
rect 57762 10402 58086 10440
rect 55168 10372 55774 10402
rect 45718 9432 53509 10370
rect 42768 8826 42772 8904
rect 45718 8902 49342 9432
rect 49885 8902 53509 9432
rect 53762 10368 55774 10372
rect 55826 10374 56432 10402
rect 56484 10374 57090 10402
rect 57106 10374 57748 10402
rect 57800 10374 58086 10402
rect 58154 10374 58188 10470
rect 58578 10374 58598 10558
rect 62994 10535 63028 11848
rect 63652 10535 63686 11848
rect 75116 11780 75150 15472
rect 75116 11692 75174 11780
rect 59464 10374 59498 10392
rect 55826 10368 59498 10374
rect 53762 8934 55412 10368
rect 55578 10330 55636 10368
rect 55590 10282 55635 10330
rect 43642 8868 53509 8902
rect 43642 7062 43676 8868
rect 44084 8794 44110 8852
rect 44112 8794 44138 8824
rect 44220 8788 44254 8868
rect 44978 8788 45012 8868
rect 45718 8788 49342 8868
rect 49526 8788 49560 8868
rect 49885 8788 53509 8868
rect 43706 8726 43778 8764
rect 43828 8754 53509 8788
rect 43744 8158 43778 8726
rect 44084 8688 44110 8748
rect 44112 8716 44138 8748
rect 44207 8742 44208 8743
rect 44208 8741 44209 8742
rect 44208 8142 44209 8143
rect 44207 8141 44208 8142
rect 44220 8130 44254 8754
rect 44266 8742 44267 8743
rect 44965 8742 44966 8743
rect 44265 8741 44266 8742
rect 44966 8741 44967 8742
rect 44265 8142 44266 8143
rect 44966 8142 44967 8143
rect 44266 8141 44267 8142
rect 44965 8141 44966 8142
rect 44978 8130 45012 8754
rect 45024 8742 45025 8743
rect 45023 8741 45024 8742
rect 45718 8662 49342 8754
rect 49513 8742 49514 8743
rect 49514 8741 49515 8742
rect 45023 8142 45024 8143
rect 45024 8141 45025 8142
rect 45718 8130 49450 8662
rect 49514 8142 49515 8143
rect 49513 8141 49514 8142
rect 49526 8130 49560 8754
rect 49572 8742 49573 8743
rect 49571 8741 49572 8742
rect 49885 8668 53509 8754
rect 49571 8142 49572 8143
rect 49572 8141 49573 8142
rect 49720 8130 53509 8668
rect 43706 8068 43778 8106
rect 43828 8096 53509 8130
rect 44207 8084 44208 8085
rect 44208 8083 44209 8084
rect 43744 7500 43778 8068
rect 44090 7478 44110 7542
rect 44118 7478 44138 7514
rect 44208 7484 44209 7485
rect 44207 7483 44208 7484
rect 44220 7472 44254 8096
rect 44266 8084 44267 8085
rect 44965 8084 44966 8085
rect 44265 8083 44266 8084
rect 44966 8083 44967 8084
rect 44265 7484 44266 7485
rect 44966 7484 44967 7485
rect 44266 7483 44267 7484
rect 44965 7483 44966 7484
rect 44978 7472 45012 8096
rect 45024 8084 45025 8085
rect 45023 8083 45024 8084
rect 45023 7484 45024 7485
rect 45024 7483 45025 7484
rect 45718 7472 49450 8096
rect 49513 8084 49514 8085
rect 49514 8083 49515 8084
rect 49476 7478 49484 7556
rect 49514 7484 49515 7485
rect 49513 7483 49514 7484
rect 49526 7472 49560 8096
rect 49572 8084 49573 8085
rect 49571 8083 49572 8084
rect 49571 7484 49572 7485
rect 49572 7483 49573 7484
rect 49720 7472 53509 8096
rect 43706 7410 43778 7448
rect 43828 7438 53509 7472
rect 43744 7064 43778 7410
rect 44090 7378 44110 7432
rect 44118 7406 44138 7432
rect 44207 7426 44208 7427
rect 44208 7425 44209 7426
rect 43706 7062 43778 7064
rect 44220 7062 44254 7438
rect 44266 7426 44267 7427
rect 44965 7426 44966 7427
rect 44265 7425 44266 7426
rect 44966 7425 44967 7426
rect 44978 7062 45012 7438
rect 45024 7426 45025 7427
rect 45023 7425 45024 7426
rect 45718 7224 49450 7438
rect 49476 7346 49484 7432
rect 49513 7426 49514 7427
rect 49514 7425 49515 7426
rect 45718 7062 49342 7224
rect 49526 7062 49560 7438
rect 49572 7426 49573 7427
rect 49571 7425 49572 7426
rect 49720 7230 53509 7438
rect 49885 7062 53509 7230
rect 54712 7164 54738 8934
rect 54740 7164 54794 8934
rect 54832 7062 54866 8934
rect 54914 7062 54924 7164
rect 54992 7062 55026 8934
rect 55106 7062 55151 8934
rect 55590 7062 55624 10282
rect 55666 9810 55686 10362
rect 55664 8800 55686 9810
rect 55722 9754 55742 10362
rect 55753 10318 55809 10329
rect 55720 8800 55742 9754
rect 55764 10282 55809 10318
rect 55764 9514 55798 10282
rect 55866 9706 59498 10368
rect 59890 10058 59900 10416
rect 60033 10397 60702 10535
rect 60720 10403 60748 10416
rect 60776 10403 60804 10416
rect 60870 10397 64133 10535
rect 64276 10462 64300 11568
rect 64310 10428 64334 11602
rect 60033 10363 64133 10397
rect 60033 10315 60702 10363
rect 59890 9844 59918 10058
rect 59890 9838 59900 9844
rect 55866 9636 59490 9706
rect 55764 8666 55809 9514
rect 55764 8654 55812 8666
rect 55666 7062 55686 8600
rect 55722 7062 55742 8600
rect 55764 8006 55809 8654
rect 55816 8616 55824 8654
rect 55866 8486 58580 9636
rect 58642 9454 58646 9636
rect 59420 9454 59454 9636
rect 60033 9628 60704 10315
rect 60069 9454 60103 9628
rect 60183 9454 60217 9488
rect 60545 9454 60579 9628
rect 60659 9454 60704 9628
rect 60720 9454 60748 10357
rect 60776 9704 60804 10357
rect 60870 10315 64133 10363
rect 60830 10304 64133 10315
rect 60841 9624 64133 10304
rect 64304 9834 64306 10416
rect 60841 9454 60886 9624
rect 55830 8360 58580 8486
rect 55830 8230 55836 8360
rect 55764 7062 55798 8006
rect 55866 7252 58580 8360
rect 58632 9420 60886 9454
rect 58632 9320 58666 9420
rect 58761 9352 59352 9399
rect 58684 9320 58688 9327
rect 58632 9264 58688 9320
rect 58808 9318 59352 9352
rect 59294 9271 59352 9318
rect 59420 9293 59454 9420
rect 58632 8122 58666 9264
rect 58682 8940 58688 9264
rect 58710 8968 58716 9264
rect 58735 9259 58791 9270
rect 58684 8215 58688 8940
rect 58746 8283 58791 9259
rect 58886 8734 59078 8786
rect 59306 8734 59351 9271
rect 58862 8666 59351 8734
rect 59306 8271 59351 8666
rect 59398 8486 59402 9271
rect 59372 8276 59402 8486
rect 59420 8317 59472 9293
rect 59404 8283 59472 8317
rect 59398 8271 59402 8276
rect 58761 8224 59352 8271
rect 58808 8190 59352 8224
rect 59294 8174 59352 8190
rect 59337 8159 59352 8174
rect 59420 8122 59454 8283
rect 60069 8122 60103 9420
rect 60545 9399 60579 9420
rect 60659 9399 60704 9420
rect 60171 9386 60706 9399
rect 60720 9386 60748 9420
rect 60124 9318 60141 9352
rect 60171 9318 60748 9386
rect 60171 9271 60229 9318
rect 60183 8271 60228 9271
rect 60545 8271 60579 9318
rect 60647 9271 60705 9318
rect 60720 9271 60748 9318
rect 60834 9392 60886 9420
rect 60659 8271 60704 9271
rect 60720 9270 60760 9271
rect 60709 9259 60765 9270
rect 60720 8283 60765 9259
rect 60776 8480 60788 9299
rect 60720 8271 60760 8276
rect 60171 8258 60706 8271
rect 60720 8258 60748 8271
rect 60124 8190 60141 8224
rect 60171 8190 60748 8258
rect 60776 8243 60788 8276
rect 60834 8195 60902 9392
rect 60171 8174 60229 8190
rect 60171 8159 60186 8174
rect 60183 8122 60217 8156
rect 60545 8122 60579 8190
rect 60647 8174 60705 8190
rect 60659 8122 60704 8174
rect 60720 8122 60748 8190
rect 60830 8184 60902 8195
rect 61317 8850 61351 9624
rect 60834 8122 60886 8184
rect 58632 8088 60886 8122
rect 58642 7252 58646 8088
rect 59420 7252 59454 8088
rect 60069 7542 60103 8088
rect 60183 7542 60217 8088
rect 55866 7218 59874 7252
rect 55866 7197 58580 7218
rect 58642 7197 58646 7218
rect 55866 7150 59352 7197
rect 55866 7116 59183 7150
rect 59226 7116 59352 7150
rect 55866 7110 58580 7116
rect 58636 7110 58694 7116
rect 59294 7110 59352 7116
rect 55866 7062 58590 7110
rect 31322 7028 58590 7062
rect 31334 6998 31368 7028
rect 32092 6998 32126 7028
rect 32850 6998 32884 7028
rect 33608 6998 33642 7028
rect 34366 6998 34400 7028
rect 35124 6998 35158 7028
rect 35882 6998 35916 7028
rect 36640 6998 36674 7028
rect 37054 7006 37974 7028
rect 37054 6998 37088 7006
rect 37940 6998 37974 7006
rect 38156 6998 38190 7028
rect 38244 7006 39164 7028
rect 38244 6998 38278 7006
rect 39130 6998 39164 7006
rect 39554 7014 40474 7028
rect 39554 6998 39588 7014
rect 39672 6998 39706 7014
rect 40430 6998 40474 7014
rect 40722 7022 41642 7028
rect 31334 6976 37408 6998
rect 37422 6976 38924 6998
rect 38938 6976 40588 6998
rect 31334 6960 40588 6976
rect 40722 6960 40756 7022
rect 41182 6998 41228 7022
rect 41160 6970 41228 6998
rect 41234 6970 41250 6992
rect 41160 6966 41250 6970
rect 41154 6960 41256 6966
rect 41608 6960 41642 7022
rect 41882 7026 45434 7028
rect 41882 6960 41916 7026
rect 41946 6998 41980 7026
rect 42734 6998 42738 7026
rect 41918 6960 41980 6998
rect 42676 6994 42714 6998
rect 42728 6994 42738 6998
rect 42768 6998 42772 7026
rect 43642 6998 43676 7026
rect 42768 6996 43472 6998
rect 43486 6996 43680 6998
rect 42676 6974 42738 6994
rect 42750 6974 42766 6996
rect 42676 6960 42766 6974
rect 42768 6960 43680 6996
rect 43744 6960 43778 7026
rect 44220 6998 44254 7026
rect 44978 6998 45012 7026
rect 44192 6996 44254 6998
rect 44950 6996 45012 6998
rect 44192 6974 44258 6996
rect 44266 6974 44282 6996
rect 44192 6960 44282 6974
rect 44950 6974 45016 6996
rect 45024 6974 45040 6996
rect 44950 6960 45040 6974
rect 45400 6960 45434 7026
rect 45718 6998 49342 7028
rect 49526 6998 49560 7028
rect 45708 6960 49342 6998
rect 49498 6960 49560 6998
rect 49702 7026 55582 7028
rect 49702 7014 53509 7026
rect 49702 6960 49736 7014
rect 49885 6960 53509 7014
rect 54114 6998 54576 7010
rect 54832 6998 54866 7026
rect 54914 6998 54924 7026
rect 54992 6998 55026 7026
rect 55106 6998 55151 7026
rect 54046 6996 54084 6998
rect 54098 6996 54108 6998
rect 54046 6992 54112 6996
rect 54114 6992 55330 6998
rect 54046 6960 55330 6992
rect 55548 6960 55582 7026
rect 31334 6084 31368 6960
rect 31396 6926 32132 6960
rect 32058 6920 32076 6926
rect 32086 6892 32132 6926
rect 32142 6926 32884 6960
rect 32912 6926 33648 6960
rect 32142 6920 32160 6926
rect 31328 6060 31374 6084
rect 32092 6060 32126 6892
rect 32850 6084 32884 6926
rect 33574 6920 33592 6926
rect 33602 6892 33648 6926
rect 33658 6926 34400 6960
rect 34428 6926 35164 6960
rect 33658 6920 33676 6926
rect 32844 6060 32890 6084
rect 33608 6060 33642 6892
rect 34366 6084 34400 6926
rect 35090 6920 35108 6926
rect 35118 6892 35164 6926
rect 35174 6926 35916 6960
rect 35944 6926 36680 6960
rect 35174 6920 35192 6926
rect 34360 6060 34406 6084
rect 35124 6060 35158 6892
rect 35882 6084 35916 6926
rect 36606 6920 36624 6926
rect 36634 6892 36680 6926
rect 36690 6926 38196 6960
rect 36690 6920 36708 6926
rect 35876 6060 35922 6084
rect 36640 6060 36674 6892
rect 31328 6022 33498 6060
rect 33580 6022 33642 6060
rect 34338 6028 34406 6060
rect 34332 6022 34406 6028
rect 34416 6022 34434 6028
rect 35096 6022 35158 6060
rect 35854 6028 35922 6060
rect 35848 6022 35922 6028
rect 35932 6022 35950 6028
rect 36612 6022 36674 6060
rect 36760 6028 36776 6082
rect 37054 6022 37088 6926
rect 37230 6904 37836 6926
rect 37157 6854 37213 6865
rect 37168 6142 37213 6854
rect 37168 6060 37202 6142
rect 37168 6022 37206 6060
rect 37214 6028 37264 6898
rect 37270 6028 37292 6898
rect 37386 6866 37444 6904
rect 37398 6142 37443 6866
rect 37815 6854 37871 6865
rect 37826 6142 37871 6854
rect 37398 6060 37432 6142
rect 37370 6022 37432 6060
rect 37826 6060 37860 6142
rect 37826 6022 37864 6060
rect 37940 6022 37974 6926
rect 38122 6920 38140 6926
rect 38150 6892 38196 6926
rect 38206 6946 40474 6960
rect 38206 6926 39712 6946
rect 38206 6920 38224 6926
rect 38100 6028 38102 6730
rect 38156 6060 38190 6892
rect 38128 6022 38190 6060
rect 38244 6022 38278 6926
rect 38420 6904 39026 6926
rect 38902 6866 38960 6904
rect 38347 6854 38403 6865
rect 38358 6142 38403 6854
rect 38358 6060 38392 6142
rect 38914 6084 38959 6866
rect 38982 6268 39000 6894
rect 39010 6865 39056 6866
rect 39058 6865 39084 6894
rect 39005 6854 39084 6865
rect 39010 6212 39084 6854
rect 39016 6200 39084 6212
rect 38908 6060 38959 6084
rect 38980 6060 39010 6200
rect 39016 6060 39061 6200
rect 39130 6060 39164 6926
rect 38358 6022 38396 6060
rect 38580 6022 39494 6060
rect 39554 6022 39588 6926
rect 39638 6920 39656 6926
rect 39666 6892 39712 6926
rect 39672 6878 39712 6892
rect 39714 6926 40474 6946
rect 40492 6926 41980 6960
rect 41992 6926 49560 6960
rect 49572 6926 55582 6960
rect 39714 6920 40422 6926
rect 39714 6912 40336 6920
rect 39714 6906 39740 6912
rect 39672 6874 39706 6878
rect 39714 6874 39718 6906
rect 39657 6862 39660 6873
rect 39672 6870 39712 6874
rect 39714 6870 39717 6874
rect 40362 6873 40366 6874
rect 39672 6862 39724 6870
rect 40315 6862 40371 6873
rect 39668 6772 39724 6862
rect 39668 6060 39752 6772
rect 39644 6028 39752 6060
rect 39762 6028 39780 6800
rect 40326 6142 40371 6862
rect 40390 6284 40422 6920
rect 40326 6060 40360 6142
rect 40430 6084 40474 6926
rect 40424 6060 40474 6084
rect 39644 6022 39706 6028
rect 31328 6000 31374 6022
rect 31384 6000 32126 6022
rect 31334 5920 31368 6000
rect 31396 5988 32126 6000
rect 32154 6000 32890 6022
rect 32900 6000 33642 6022
rect 32154 5988 32884 6000
rect 32912 5988 33642 6000
rect 33654 6000 34406 6022
rect 33654 5988 34400 6000
rect 34412 5988 35158 6022
rect 35170 6000 35922 6022
rect 35170 5988 35916 6000
rect 35928 5988 36674 6022
rect 36686 5988 37432 6022
rect 37444 5988 38190 6022
rect 38202 5988 38959 6022
rect 38964 6000 39706 6022
rect 38976 5988 39706 6000
rect 32092 5920 32126 5988
rect 32850 5920 32884 5988
rect 33608 5920 33642 5988
rect 34366 5920 34400 5988
rect 35044 5920 35052 5982
rect 35072 5920 35108 5982
rect 35124 5920 35158 5988
rect 35882 5920 35916 5988
rect 36640 5920 36674 5988
rect 37054 5920 37088 5988
rect 37168 5920 37202 5988
rect 37398 5920 37432 5988
rect 37826 5920 37860 5988
rect 37940 5920 37974 5988
rect 38156 5920 38190 5988
rect 38244 5920 38278 5988
rect 38358 5920 38392 5988
rect 38914 5920 38959 5988
rect 39016 5920 39061 5988
rect 39130 5920 39164 5988
rect 39554 5920 39588 5988
rect 39668 5920 39706 5988
rect 39714 5920 39717 6028
rect 40326 6022 40364 6060
rect 40402 6028 40474 6060
rect 40396 6022 40474 6028
rect 40480 6022 40498 6028
rect 40722 6022 40756 6926
rect 40898 6920 41504 6926
rect 41176 6882 41234 6920
rect 40825 6870 40870 6881
rect 40836 6060 40870 6870
rect 41188 6060 41222 6882
rect 41483 6870 41528 6881
rect 40836 6022 40874 6060
rect 41160 6022 41222 6060
rect 41494 6060 41528 6870
rect 41494 6022 41532 6060
rect 41608 6022 41642 6926
rect 41882 6028 41916 6926
rect 41946 6272 41980 6926
rect 42058 6924 42664 6926
rect 42700 6924 43322 6926
rect 43346 6924 43980 6926
rect 44032 6924 44638 6926
rect 44690 6924 45296 6926
rect 42018 6918 42020 6920
rect 42046 6918 42048 6920
rect 41990 6886 42020 6918
rect 41990 6880 42036 6886
rect 41990 6874 42062 6880
rect 41996 6474 42062 6874
rect 41996 6272 42036 6474
rect 42080 6446 42090 6908
rect 42670 6885 42688 6890
rect 42643 6874 42688 6885
rect 41946 6084 41986 6272
rect 41940 6060 41986 6084
rect 41918 6056 41986 6060
rect 41990 6056 42036 6272
rect 41918 6028 42036 6056
rect 42654 6060 42688 6874
rect 42700 6886 42750 6924
rect 42654 6056 42692 6060
rect 42700 6056 42738 6886
rect 41882 6022 42030 6028
rect 42654 6022 42738 6056
rect 42768 6060 42772 6924
rect 43346 6920 43408 6924
rect 43334 6890 43346 6920
rect 43362 6918 43408 6920
rect 43346 6885 43352 6886
rect 43301 6874 43357 6885
rect 43312 6862 43357 6874
rect 43406 6862 43432 6918
rect 43450 6886 43508 6924
rect 43312 6534 43376 6862
rect 43312 6060 43357 6534
rect 43406 6060 43408 6534
rect 43462 6060 43507 6886
rect 43642 6060 43676 6924
rect 43744 6842 43778 6924
rect 44208 6886 44266 6924
rect 44966 6886 45024 6924
rect 43959 6874 44004 6885
rect 43970 6814 44004 6874
rect 44220 6814 44254 6886
rect 44617 6874 44662 6885
rect 44628 6814 44662 6874
rect 44978 6814 45012 6886
rect 45275 6874 45320 6885
rect 45286 6814 45320 6874
rect 45400 6814 45434 6926
rect 45718 6814 49342 6926
rect 49476 6820 49484 6898
rect 49514 6826 49515 6827
rect 49513 6825 49514 6826
rect 49526 6814 49560 6926
rect 49571 6826 49572 6827
rect 49572 6825 49573 6826
rect 49702 6814 49736 6926
rect 49878 6912 53509 6926
rect 53522 6924 54786 6926
rect 54822 6924 55444 6926
rect 49805 6862 49850 6873
rect 49816 6814 49850 6862
rect 49885 6814 53509 6912
rect 54062 6886 54108 6924
rect 43706 6752 43778 6790
rect 43828 6780 53509 6814
rect 43744 6184 43778 6752
rect 43970 6156 44004 6780
rect 44220 6156 44254 6780
rect 44628 6156 44662 6780
rect 44978 6156 45012 6780
rect 45286 6156 45320 6780
rect 45400 6156 45434 6780
rect 45662 6774 49342 6780
rect 45718 6772 49342 6774
rect 45690 6746 49342 6772
rect 45718 6156 49342 6746
rect 49476 6682 49484 6774
rect 49513 6768 49514 6769
rect 49514 6767 49515 6768
rect 49514 6168 49515 6169
rect 49513 6167 49514 6168
rect 49526 6156 49560 6780
rect 49572 6768 49573 6769
rect 49571 6767 49572 6768
rect 49571 6168 49572 6169
rect 49572 6167 49573 6168
rect 49702 6156 49736 6780
rect 49816 6156 49850 6780
rect 49885 6156 53509 6780
rect 43706 6094 43778 6132
rect 43828 6122 53509 6156
rect 42768 6022 43680 6060
rect 43744 6022 43778 6094
rect 43970 6060 44004 6122
rect 44220 6060 44254 6122
rect 43970 6022 44008 6060
rect 44192 6022 44254 6060
rect 44628 6060 44662 6122
rect 44978 6060 45012 6122
rect 44628 6022 44666 6060
rect 44950 6022 45012 6060
rect 45286 6060 45320 6122
rect 45286 6022 45324 6060
rect 45400 6022 45434 6122
rect 45718 6060 49342 6122
rect 49513 6110 49514 6111
rect 49514 6109 49515 6110
rect 49526 6060 49560 6122
rect 49572 6110 49573 6111
rect 49571 6109 49572 6110
rect 45708 6022 49342 6060
rect 49498 6022 49560 6060
rect 49702 6022 49736 6122
rect 49816 6060 49850 6122
rect 49816 6022 49854 6060
rect 49885 6022 53509 6122
rect 54074 6060 54108 6886
rect 54114 6372 54576 6924
rect 54822 6886 54878 6924
rect 54765 6874 54820 6885
rect 54776 6590 54820 6874
rect 54712 6554 54738 6590
rect 54740 6582 54820 6590
rect 54714 6448 54738 6554
rect 54770 6448 54820 6582
rect 54046 6056 54108 6060
rect 54118 6056 54152 6372
rect 54046 6022 54152 6056
rect 54172 6288 54522 6322
rect 54172 6022 54206 6288
rect 54292 6220 54402 6258
rect 54330 6186 54402 6220
rect 54275 6136 54331 6147
rect 54363 6136 54419 6147
rect 54286 6060 54331 6136
rect 54374 6060 54419 6136
rect 54488 6060 54522 6288
rect 54776 6248 54820 6448
rect 54714 6144 54738 6248
rect 54770 6144 54820 6248
rect 54776 6060 54820 6144
rect 54250 6056 54820 6060
rect 54822 6060 54877 6886
rect 54992 6060 55026 6924
rect 55106 6060 55151 6924
rect 55423 6874 55468 6885
rect 55434 6060 55468 6874
rect 54822 6056 55330 6060
rect 54250 6022 55330 6056
rect 55434 6022 55472 6060
rect 55548 6022 55582 6926
rect 39718 5988 40474 6022
rect 40476 5988 41222 6022
rect 41234 6000 41986 6022
rect 41990 6000 42738 6022
rect 41234 5988 41980 6000
rect 41992 5988 42738 6000
rect 42750 5988 43507 6022
rect 43524 5988 44254 6022
rect 44266 5988 45012 6022
rect 45024 5988 49560 6022
rect 49572 5988 54108 6022
rect 40326 5920 40360 5988
rect 40430 5920 40474 5988
rect 40722 5920 40756 5988
rect 40836 5920 40870 5988
rect 41188 5920 41222 5988
rect 41494 5920 41528 5988
rect 41608 5920 41642 5988
rect 41882 5920 41916 5988
rect 41946 5920 41980 5988
rect 41996 5920 42030 5988
rect 42654 5920 42688 5988
rect 42700 5920 42738 5988
rect 42768 5920 42772 5988
rect 43312 5920 43357 5988
rect 43462 5920 43507 5988
rect 43642 5920 43676 5988
rect 43744 5924 43778 5988
rect 43706 5920 43816 5924
rect 43970 5920 44004 5988
rect 44220 5920 44254 5988
rect 44628 5920 44662 5988
rect 44978 5920 45012 5988
rect 45286 5920 45320 5988
rect 45400 5920 45434 5988
rect 45718 5936 49342 5988
rect 45736 5920 45770 5936
rect 46494 5920 46528 5936
rect 47202 5920 47236 5936
rect 47252 5920 47286 5936
rect 47316 5920 47350 5936
rect 47974 5920 48008 5936
rect 48010 5920 48044 5936
rect 48088 5920 48122 5936
rect 48392 5920 48426 5936
rect 48506 5920 48540 5936
rect 48768 5920 48802 5936
rect 49164 5920 49198 5936
rect 49278 5920 49312 5936
rect 49526 5920 49560 5988
rect 49702 5920 49736 5988
rect 49816 5920 49850 5988
rect 49885 5920 53509 5988
rect 54074 5920 54108 5988
rect 54118 5988 54877 6022
rect 54894 5988 55582 6022
rect 54118 5920 54152 5988
rect 54172 5920 54206 5988
rect 54286 5960 54331 5988
rect 54374 5960 54419 5988
rect 54296 5924 54398 5944
rect 54292 5920 54402 5924
rect 54488 5920 54522 5988
rect 54776 5920 54820 5988
rect 54822 5920 54877 5988
rect 54992 5920 55026 5988
rect 55106 5920 55151 5988
rect 55434 5920 55468 5988
rect 55548 5920 55582 5988
rect 55590 5920 55624 7028
rect 55666 6966 55686 7028
rect 55722 6966 55742 7028
rect 55764 6998 55798 7028
rect 55764 6960 55802 6998
rect 55866 6960 58590 7028
rect 55636 6926 58590 6960
rect 55666 6028 55686 6920
rect 55722 6028 55742 6920
rect 55764 6060 55798 6926
rect 55866 6569 58590 6926
rect 58598 7069 58694 7110
rect 58598 6569 58646 7069
rect 58648 6569 58693 7069
rect 59153 7057 59209 7068
rect 59164 6581 59209 7057
rect 59226 6569 59240 7110
rect 59254 7069 59352 7110
rect 59254 6569 59296 7069
rect 59306 6569 59351 7069
rect 59420 6888 59454 7218
rect 59370 6860 59546 6888
rect 59370 6842 59490 6860
rect 59370 6826 59546 6842
rect 55866 6522 59352 6569
rect 55866 6488 59183 6522
rect 59226 6488 59352 6522
rect 55866 6420 58580 6488
rect 58636 6472 58694 6488
rect 59294 6472 59352 6488
rect 58642 6420 58646 6472
rect 59337 6457 59352 6472
rect 59420 6420 59454 6826
rect 59490 6824 59546 6826
rect 55866 6386 59874 6420
rect 55764 6022 55802 6060
rect 55866 6022 58580 6386
rect 58642 6368 58646 6386
rect 58620 6160 58646 6368
rect 58642 6155 58646 6160
rect 59420 6068 59454 6386
rect 60033 6350 60260 7542
rect 55636 5988 58580 6022
rect 55666 5920 55686 5982
rect 55722 5920 55742 5982
rect 55764 5920 55798 5988
rect 55866 5936 58580 5988
rect 56348 5920 56382 5936
rect 56422 5920 56462 5936
rect 56482 5920 56518 5936
rect 57080 5920 57151 5936
rect 57738 5920 57783 5936
rect 57864 5920 57909 5936
rect 57978 5920 58012 5936
rect 31316 5886 58012 5920
rect 32092 4242 32126 5886
rect 32850 4242 32884 5886
rect 35044 5354 35052 5886
rect 35072 5382 35108 5886
rect 37054 5726 37088 5886
rect 37168 5878 37213 5886
rect 37398 5866 37443 5886
rect 37826 5878 37871 5886
rect 37192 5828 37836 5866
rect 37230 5794 37836 5828
rect 37386 5778 37444 5794
rect 37398 5726 37432 5778
rect 37940 5726 37974 5886
rect 37054 5692 37974 5726
rect 30216 4224 33784 4242
rect 30216 4222 30760 4224
rect 31098 4214 33784 4224
rect 31220 4186 31254 4214
rect 32092 4186 32126 4214
rect 32850 4186 32884 4214
rect 30216 4168 33784 4186
rect 30216 4166 30816 4168
rect 31042 4158 33784 4168
rect 24334 3531 27958 3567
rect 28650 3536 30023 3567
rect 31220 3536 31254 4158
rect 31334 3536 31368 3596
rect 32092 3558 32126 4158
rect 32850 3558 32884 4158
rect 37398 3567 37432 5692
rect 38156 3567 38190 5886
rect 38244 5726 38278 5886
rect 38358 5878 38403 5886
rect 38914 5866 38959 5886
rect 39016 5878 39061 5886
rect 38382 5828 39026 5866
rect 38420 5794 39026 5828
rect 38902 5778 38960 5794
rect 38914 5726 38948 5778
rect 39130 5726 39164 5886
rect 38244 5692 39164 5726
rect 38508 5254 38848 5290
rect 38876 5254 38890 5492
rect 38470 5216 38810 5252
rect 38914 3567 38948 5692
rect 39554 5134 39588 5886
rect 39668 5286 39706 5886
rect 39672 5274 39706 5286
rect 39714 5274 39717 5886
rect 40326 5286 40371 5886
rect 39672 5236 40336 5274
rect 39672 5134 39706 5236
rect 39714 5186 39718 5236
rect 39730 5202 40336 5236
rect 40440 5134 40474 5886
rect 39554 5100 40474 5134
rect 40722 5142 40756 5886
rect 40836 5294 40881 5886
rect 41188 5282 41233 5886
rect 41494 5294 41539 5886
rect 40860 5244 41504 5282
rect 40898 5210 41504 5244
rect 41176 5194 41234 5210
rect 41188 5142 41222 5194
rect 41608 5142 41642 5886
rect 40722 5108 41642 5142
rect 31372 3536 32884 3558
rect 28650 3531 35058 3536
rect 24334 3502 35058 3531
rect 24334 3497 30023 3502
rect 18502 1126 21794 2097
rect 18278 1092 21794 1126
rect 18290 296 18324 1092
rect 18502 1024 21794 1092
rect 18336 990 21794 1024
rect 18502 882 21794 990
rect 21806 882 21828 2097
rect 21886 1788 21914 2097
rect 21942 882 21987 2097
rect 22056 882 22090 2097
rect 18502 848 22464 882
rect 18502 818 21794 848
rect 21806 818 21828 848
rect 21942 818 21987 848
rect 22056 818 22090 848
rect 22418 818 22452 848
rect 18502 780 21798 818
rect 21806 780 22452 818
rect 18502 746 22452 780
rect 14239 42 17856 60
rect 18140 42 18376 296
rect 14239 2 17892 42
rect 18136 6 18376 42
rect 18502 6 21794 746
rect 14239 -106 14273 2
rect 14239 -134 14284 -106
rect 14715 -134 14749 2
rect 14758 -130 14804 2
rect 14832 -74 14860 2
rect 14832 -130 14876 -74
rect 14758 -134 14820 -130
rect 14222 -168 14292 -134
rect 11996 -202 14292 -168
rect 11996 -399 12080 -202
rect 12562 -223 12596 -202
rect 12562 -270 12609 -223
rect 12624 -264 12638 -202
rect 12652 -264 12694 -202
rect 12704 -223 12738 -202
rect 12818 -223 12852 -202
rect 12704 -270 12751 -223
rect 12774 -270 12852 -223
rect 13220 -254 13266 -223
rect 13208 -270 13266 -254
rect 12206 -304 12852 -270
rect 12864 -304 13266 -270
rect 12133 -363 12178 -352
rect 12144 -399 12178 -363
rect 12562 -387 12596 -304
rect 12704 -399 12738 -304
rect 12818 -329 12852 -304
rect 12818 -352 12870 -329
rect 13208 -351 13266 -304
rect 12791 -363 12870 -352
rect 12802 -399 12870 -363
rect 13220 -387 13254 -351
rect 11996 -440 12092 -399
rect 9264 -446 11978 -440
rect 12030 -446 12092 -440
rect 12144 -446 12191 -399
rect 12534 -446 12581 -399
rect 12692 -446 12750 -399
rect 12790 -446 12870 -399
rect 13192 -446 13239 -399
rect 9264 -480 12581 -446
rect 12624 -480 13239 -446
rect 9264 -548 11978 -480
rect 12030 -496 12092 -480
rect 12030 -548 12086 -496
rect 12108 -548 12114 -486
rect 12144 -530 12178 -480
rect 12692 -496 12750 -480
rect 12790 -496 12870 -480
rect 12704 -530 12738 -496
rect 12144 -548 12189 -530
rect 12704 -548 12749 -530
rect 12796 -548 12800 -496
rect 12818 -514 12870 -496
rect 12802 -548 12870 -514
rect 13334 -548 13368 -202
rect 13433 -304 13448 -270
rect 9264 -582 13368 -548
rect 9264 -813 11978 -582
rect 12030 -600 12086 -582
rect 12108 -600 12114 -582
rect 12018 -808 12080 -600
rect 12082 -808 12114 -654
rect 12030 -813 12086 -808
rect 12138 -813 12142 -654
rect 12144 -813 12189 -582
rect 12704 -813 12749 -582
rect 9264 -860 12749 -813
rect 9264 -894 12086 -860
rect 9264 -962 11978 -894
rect 12012 -900 12086 -894
rect 12096 -894 12749 -860
rect 12096 -900 12114 -894
rect 12030 -956 12086 -900
rect 12030 -962 12080 -956
rect 12082 -962 12086 -956
rect 12144 -962 12189 -894
rect 12260 -956 12749 -894
rect 12704 -962 12749 -956
rect 12796 -962 12800 -582
rect 12818 -962 12870 -582
rect 9264 -996 12870 -962
rect 9162 -1154 9202 -1124
rect 9264 -1136 11978 -996
rect 9228 -1152 11978 -1136
rect 9222 -1154 11978 -1152
rect 8692 -1334 9014 -1312
rect 7554 -2198 8646 -2176
rect 7554 -2202 8606 -2198
rect 8082 -2396 8108 -2202
rect 8138 -2396 8164 -2202
rect 8174 -2556 8208 -2202
rect 8174 -2562 8270 -2556
rect 8390 -2562 8424 -2202
rect 8504 -2562 8549 -2202
rect 8832 -2396 8866 -1334
rect 8832 -2562 8877 -2396
rect 8946 -2562 8980 -1334
rect 3283 -2574 8980 -2562
rect 9162 -2574 9196 -1154
rect 9228 -1262 11978 -1154
rect 9228 -1392 9234 -1262
rect 9264 -2370 11978 -1262
rect 12030 -1500 12064 -996
rect 12082 -1407 12086 -996
rect 12144 -1062 12189 -996
rect 12704 -1062 12749 -996
rect 12144 -1339 12178 -1062
rect 12704 -1351 12738 -1062
rect 12740 -1136 12772 -1062
rect 12796 -1136 12800 -996
rect 12740 -1346 12800 -1136
rect 12818 -1305 12870 -996
rect 12802 -1339 12870 -1305
rect 12740 -1351 12772 -1346
rect 12796 -1351 12800 -1346
rect 12692 -1398 12772 -1351
rect 12206 -1432 12750 -1398
rect 12692 -1448 12772 -1432
rect 12706 -1463 12772 -1448
rect 12706 -1500 12738 -1463
rect 12740 -1500 12772 -1463
rect 12818 -1500 12852 -1339
rect 13467 -1500 13501 -202
rect 13581 -239 13615 -202
rect 13569 -254 13615 -239
rect 13569 -270 13627 -254
rect 13943 -270 13977 -202
rect 13986 -223 14020 -202
rect 13986 -270 14033 -223
rect 14057 -270 14091 -202
rect 14100 -270 14146 -202
rect 13506 -304 13539 -270
rect 13569 -304 14146 -270
rect 13569 -351 13627 -304
rect 13581 -530 13615 -351
rect 13943 -462 13977 -304
rect 13986 -462 14020 -304
rect 13581 -1351 13626 -530
rect 13800 -552 14020 -462
rect 14057 -530 14091 -304
rect 14100 -351 14146 -304
rect 14100 -407 14158 -351
rect 14118 -444 14158 -407
rect 14174 -444 14186 -323
rect 14222 -403 14292 -202
rect 14698 -398 14820 -134
rect 14832 -398 14848 -130
rect 14118 -450 14152 -444
rect 14222 -450 14594 -403
rect 14698 -444 14804 -398
rect 14832 -444 14876 -398
rect 14698 -450 14768 -444
rect 14118 -484 14768 -450
rect 14118 -490 14152 -484
rect 14118 -530 14158 -490
rect 14057 -552 14102 -530
rect 14118 -552 14163 -530
rect 14174 -552 14186 -490
rect 14222 -552 14688 -484
rect 14698 -490 14768 -484
rect 14780 -490 14804 -444
rect 14808 -450 14876 -444
rect 14897 -450 14931 2
rect 15373 -403 15407 2
rect 15361 -450 15407 -403
rect 15416 -407 15466 2
rect 14808 -484 15407 -450
rect 14808 -490 14860 -484
rect 14698 -546 14804 -490
rect 14698 -552 14768 -546
rect 14776 -552 14804 -546
rect 14832 -552 14860 -490
rect 14897 -530 14931 -484
rect 14897 -552 14942 -530
rect 14952 -552 15334 -484
rect 15361 -500 15407 -484
rect 15373 -530 15407 -500
rect 15373 -552 15418 -530
rect 15438 -552 15466 -407
rect 15494 -552 15522 2
rect 15530 -150 15589 2
rect 16031 -150 16065 2
rect 16072 -150 16106 2
rect 15530 -462 15604 -150
rect 15530 -552 15810 -462
rect 16010 -470 16106 -150
rect 13800 -586 15810 -552
rect 13800 -894 14012 -586
rect 13666 -910 14012 -894
rect 13666 -956 13977 -910
rect 13943 -1351 13977 -956
rect 14057 -1351 14102 -586
rect 14118 -1339 14163 -586
rect 14174 -1142 14186 -586
rect 14222 -590 14688 -586
rect 14698 -590 14768 -586
rect 14232 -910 14688 -590
rect 13522 -1432 13539 -1398
rect 13569 -1432 14102 -1351
rect 13569 -1448 13627 -1432
rect 13569 -1463 13615 -1448
rect 13581 -1500 13615 -1463
rect 13943 -1500 13977 -1432
rect 14057 -1500 14102 -1432
rect 14118 -1351 14158 -1346
rect 14118 -1500 14146 -1351
rect 14174 -1379 14186 -1346
rect 14232 -1500 14284 -910
rect 14476 -918 14688 -910
rect 14504 -998 14672 -918
rect 12030 -1534 14284 -1500
rect 12040 -2370 12044 -1534
rect 12706 -1982 12738 -1534
rect 12740 -1948 12772 -1534
rect 12818 -2370 12852 -1534
rect 13467 -2080 13501 -1534
rect 13581 -2080 13615 -1534
rect 9264 -2404 13272 -2370
rect 9264 -2472 11978 -2404
rect 12040 -2456 12044 -2404
rect 12046 -2456 12093 -2425
rect 12034 -2472 12093 -2456
rect 12534 -2472 12581 -2425
rect 12704 -2456 12750 -2425
rect 12692 -2472 12750 -2456
rect 9264 -2506 12581 -2472
rect 12624 -2506 12750 -2472
rect 9264 -2512 11978 -2506
rect 12034 -2512 12092 -2506
rect 12692 -2512 12750 -2506
rect 9264 -2574 11988 -2512
rect 3100 -2608 11988 -2574
rect 3100 -2808 3134 -2608
rect 3283 -2638 11988 -2608
rect 3238 -2676 11988 -2638
rect 3276 -2710 11988 -2676
rect 3180 -2724 3282 -2720
rect 3208 -2749 3254 -2748
rect 3203 -2752 3259 -2749
rect 3203 -2760 3270 -2752
rect 3214 -2796 3270 -2760
rect 3214 -2808 3248 -2796
rect 3252 -2797 3270 -2796
rect 3283 -2797 11988 -2710
rect 3252 -2802 11988 -2797
rect 3260 -2808 11988 -2802
rect -884 -2842 2744 -2808
rect 3066 -2842 11988 -2808
rect -884 -3466 2740 -2842
rect 3100 -3466 3134 -2842
rect 3214 -2854 3248 -2842
rect 3252 -2854 3270 -2848
rect 3214 -2940 3270 -2854
rect 3214 -3453 3259 -2940
rect 3283 -3094 11988 -2842
rect 11996 -2553 12092 -2512
rect 11996 -3053 12044 -2553
rect 12046 -3053 12080 -2553
rect 12551 -2565 12596 -2554
rect 12562 -3041 12596 -2565
rect 11996 -3094 12093 -3053
rect 3283 -3100 11978 -3094
rect 12034 -3100 12093 -3094
rect 12534 -3100 12581 -3053
rect 12624 -3094 12638 -2512
rect 12652 -2553 12750 -2512
rect 12652 -3053 12694 -2553
rect 12704 -3053 12738 -2553
rect 12818 -2734 12852 -2404
rect 12768 -2796 13064 -2734
rect 12652 -3094 12750 -3053
rect 12692 -3100 12750 -3094
rect 3283 -3134 12581 -3100
rect 12624 -3134 12750 -3100
rect 3283 -3202 11978 -3134
rect 12034 -3150 12092 -3134
rect 12692 -3150 12750 -3134
rect 12040 -3202 12044 -3150
rect 12735 -3165 12750 -3150
rect 12818 -3202 12852 -2796
rect 12888 -3202 13404 -3180
rect 3283 -3236 13404 -3202
rect 3214 -3454 3260 -3453
rect 3214 -3466 3248 -3454
rect 3252 -3460 3254 -3454
rect 3260 -3455 3261 -3454
rect 3283 -3455 11978 -3236
rect 12040 -3254 12044 -3236
rect 12018 -3280 12044 -3254
rect 12046 -3455 12080 -3236
rect 3260 -3466 11978 -3455
rect -2896 -3524 -2786 -3490
rect -2774 -3500 -1134 -3466
rect -884 -3500 2744 -3466
rect 3066 -3468 11978 -3466
rect 12692 -3467 12750 -3416
rect 3066 -3500 6907 -3468
rect -2645 -3512 -2644 -3511
rect -2632 -3512 -2598 -3500
rect -2586 -3512 -2585 -3511
rect -1987 -3512 -1986 -3511
rect -1974 -3512 -1940 -3500
rect -1928 -3512 -1927 -3511
rect -1329 -3512 -1328 -3511
rect -1316 -3512 -1282 -3500
rect -2644 -3513 -2643 -3512
rect -2632 -3513 -2586 -3512
rect -1986 -3513 -1985 -3512
rect -1974 -3513 -1928 -3512
rect -1328 -3513 -1327 -3512
rect -2896 -3528 -2764 -3524
rect -2858 -3538 -2764 -3528
rect -2858 -3924 -2786 -3538
rect -2632 -3924 -2587 -3513
rect -1974 -3924 -1929 -3513
rect -1316 -3924 -1271 -3512
rect -2858 -4096 -2824 -3924
rect -2644 -4112 -2643 -4111
rect -2645 -4113 -2644 -4112
rect -2632 -4124 -2598 -3924
rect -2587 -4112 -2586 -4111
rect -1986 -4112 -1985 -4111
rect -2586 -4113 -2585 -4112
rect -1987 -4113 -1986 -4112
rect -1974 -4124 -1940 -3924
rect -1929 -4112 -1928 -4111
rect -1328 -4112 -1327 -4111
rect -1928 -4113 -1927 -4112
rect -1329 -4113 -1328 -4112
rect -1316 -4124 -1282 -3924
rect -1202 -4124 -1168 -3500
rect -884 -3686 2740 -3500
rect 600 -3896 634 -3686
rect 714 -3744 759 -3686
rect 1372 -3744 1417 -3686
rect 738 -3794 1382 -3756
rect 776 -3828 1382 -3794
rect 1486 -3896 1520 -3686
rect 600 -3930 1520 -3896
rect 1790 -3896 1824 -3686
rect 1904 -3744 1949 -3686
rect 2562 -3744 2607 -3686
rect 1928 -3794 2572 -3756
rect 1966 -3828 2572 -3794
rect 2676 -3896 2710 -3686
rect 1790 -3930 2710 -3896
rect 1962 -4040 2512 -4038
rect 1990 -4068 2484 -4066
rect 3100 -4124 3134 -3500
rect 3214 -3512 3248 -3500
rect 3252 -3512 3254 -3506
rect 3260 -3512 3261 -3511
rect 3214 -3513 3260 -3512
rect 3214 -3924 3259 -3513
rect 3214 -4124 3248 -3924
rect 3252 -4118 3254 -4040
rect 3259 -4112 3260 -4111
rect 3260 -4113 3261 -4112
rect 3283 -4124 6907 -3500
rect -2774 -4158 -1168 -4124
rect 0 -4158 6907 -4124
rect -2632 -4238 -2598 -4158
rect -1974 -4238 -1940 -4158
rect -1316 -4238 -1282 -4158
rect -1202 -4238 -1168 -4158
rect 3100 -4238 3134 -4158
rect 3214 -4238 3248 -4158
rect 3252 -4238 3254 -4164
rect 3283 -4238 6907 -4158
rect -2960 -4272 6907 -4238
rect -2058 -4656 -2040 -4272
rect -2002 -4656 -1984 -4324
rect -2818 -4744 -2270 -4710
rect -2818 -5026 -2784 -4744
rect -2632 -4824 -2598 -4744
rect -2456 -4824 -2445 -4813
rect -2754 -4868 -2682 -4830
rect -2716 -4902 -2682 -4868
rect -2632 -4858 -2445 -4824
rect -2645 -4870 -2644 -4869
rect -2644 -4871 -2643 -4870
rect -2644 -4900 -2643 -4899
rect -2645 -4901 -2644 -4900
rect -2632 -4912 -2598 -4858
rect -2444 -4868 -2372 -4830
rect -2586 -4870 -2585 -4869
rect -2587 -4871 -2586 -4870
rect -2587 -4900 -2586 -4899
rect -2586 -4901 -2585 -4900
rect -2456 -4912 -2445 -4901
rect -2406 -4902 -2372 -4868
rect -2632 -4946 -2445 -4912
rect -2632 -5026 -2598 -4946
rect -2304 -5026 -2270 -4744
rect -2818 -5060 -2270 -5026
rect -2220 -5118 -1582 -4656
rect -2058 -5132 -2040 -5118
rect -2002 -5132 -1984 -5118
rect -2818 -5220 -2270 -5186
rect -2818 -5502 -2784 -5220
rect -2632 -5300 -2598 -5220
rect -2456 -5300 -2445 -5289
rect -2754 -5340 -2682 -5306
rect -2632 -5334 -2445 -5300
rect -2754 -5344 -2674 -5340
rect -2716 -5378 -2674 -5344
rect -2645 -5346 -2644 -5345
rect -2644 -5347 -2643 -5346
rect -2644 -5376 -2643 -5375
rect -2645 -5377 -2644 -5376
rect -2700 -5394 -2674 -5378
rect -2644 -5396 -2638 -5382
rect -2632 -5388 -2598 -5334
rect -2444 -5344 -2372 -5306
rect -2586 -5346 -2585 -5345
rect -2587 -5347 -2586 -5346
rect -2587 -5376 -2586 -5375
rect -2586 -5377 -2585 -5376
rect -2592 -5388 -2538 -5382
rect -2456 -5388 -2445 -5377
rect -2406 -5378 -2372 -5344
rect -2632 -5422 -2445 -5388
rect -2632 -5502 -2598 -5422
rect -2304 -5502 -2270 -5220
rect -2818 -5536 -2270 -5502
rect -2220 -5594 -1582 -5132
rect -1322 -5322 -1320 -4308
rect -1202 -6014 -1168 -4272
rect 3100 -4426 3134 -4272
rect 3252 -4348 3254 -4272
rect 3283 -4308 6907 -4272
rect 3283 -4558 4056 -4308
rect -14036 -6046 -13956 -6032
rect -13560 -6046 -13474 -6032
rect -16054 -6110 -12598 -6076
rect -14930 -7280 -14896 -6110
rect -14272 -7280 -14238 -6110
rect -17676 -7324 -17416 -7290
rect -17676 -7370 -17642 -7324
rect -14158 -7370 -14124 -6110
rect -13740 -6146 -13278 -6110
rect -13264 -6146 -12802 -6110
rect -13264 -6726 -13024 -6146
rect 3319 -7393 3353 -4558
rect 3433 -4652 3467 -4558
rect 4057 -4652 4062 -4478
rect 4091 -4652 4125 -4308
rect 4232 -4550 5224 -4308
rect 4749 -4652 4783 -4550
rect 5392 -4652 6907 -4308
rect 3433 -4693 4062 -4652
rect 4063 -4665 4125 -4652
rect 4063 -4693 4131 -4665
rect 3433 -4699 4131 -4693
rect 4141 -4699 4159 -4693
rect 4222 -4699 5234 -4652
rect 5379 -4693 6907 -4652
rect 5373 -4699 6907 -4693
rect 3433 -4700 3467 -4699
rect 3495 -4700 4131 -4699
rect 3433 -4767 3473 -4700
rect 3483 -4733 4131 -4700
rect 4137 -4733 4783 -4699
rect 4811 -4733 6907 -4699
rect 3483 -4739 3501 -4733
rect 4057 -4739 4075 -4733
rect 3433 -4801 3467 -4767
rect 4057 -4801 4062 -4739
rect 4085 -4767 4131 -4733
rect 4141 -4739 4159 -4733
rect 4091 -4801 4125 -4767
rect 4749 -4801 4783 -4733
rect 5373 -4739 5391 -4733
rect 5392 -4801 6907 -4733
rect 3415 -4835 6907 -4801
rect 3433 -5924 3467 -4835
rect 4057 -6066 4062 -4835
rect 4091 -6066 4096 -4835
rect 4749 -5924 4783 -4835
rect 5392 -5228 6907 -4835
rect 7516 -4600 7550 -3468
rect 7570 -3814 7604 -3468
rect 7673 -3486 7729 -3475
rect 7761 -3486 7817 -3475
rect 7684 -3662 7729 -3486
rect 7772 -3662 7817 -3486
rect 7690 -3712 7800 -3674
rect 7728 -3746 7800 -3712
rect 7886 -3814 7920 -3468
rect 7570 -3848 7920 -3814
rect 7566 -4026 7584 -3924
rect 7516 -4856 7556 -4600
rect 7564 -4828 7584 -4628
rect 7516 -5228 7550 -4856
rect 8084 -5050 8108 -4026
rect 8140 -4266 8164 -4026
rect 8174 -5228 8208 -3468
rect 8390 -4778 8424 -3468
rect 8504 -4638 8549 -3468
rect 8832 -3924 8877 -3468
rect 8832 -4638 8866 -3924
rect 8504 -4676 8728 -4638
rect 8832 -4676 8870 -4638
rect 8946 -4676 8980 -3468
rect 9162 -4638 9196 -3468
rect 9264 -3616 11978 -3468
rect 12362 -3492 12750 -3470
rect 12362 -3504 12714 -3492
rect 12362 -3564 12396 -3504
rect 12500 -3548 12614 -3534
rect 12818 -3554 12852 -3236
rect 12888 -3272 13404 -3236
rect 13431 -3272 13658 -2080
rect 12362 -3566 12373 -3564
rect 12385 -3566 12396 -3564
rect 12362 -3616 12396 -3566
rect 12538 -3586 12576 -3572
rect 12718 -3616 12752 -3566
rect 9264 -3650 12756 -3616
rect 9264 -3686 11978 -3650
rect 9820 -4638 9854 -3686
rect 10478 -4638 10512 -3686
rect 11136 -4638 11170 -3686
rect 11794 -4638 11828 -3686
rect 9134 -4642 9196 -4638
rect 9792 -4642 9854 -4638
rect 10450 -4642 10512 -4638
rect 11108 -4642 11170 -4638
rect 9134 -4670 9202 -4642
rect 9792 -4670 9860 -4642
rect 10450 -4670 10518 -4642
rect 11108 -4670 11176 -4642
rect 11766 -4670 11828 -4638
rect 9128 -4676 9202 -4670
rect 9212 -4676 9230 -4670
rect 9786 -4676 9860 -4670
rect 9870 -4676 9888 -4670
rect 10444 -4676 10518 -4670
rect 10528 -4676 10546 -4670
rect 11102 -4676 11176 -4670
rect 11186 -4676 11204 -4670
rect 11760 -4676 11828 -4670
rect 8504 -4778 8549 -4676
rect 8566 -4710 9202 -4676
rect 9208 -4710 9860 -4676
rect 9866 -4710 10518 -4676
rect 10524 -4710 11176 -4676
rect 11182 -4710 11828 -4676
rect 8832 -4774 8866 -4710
rect 8832 -4778 8877 -4774
rect 8946 -4778 8980 -4710
rect 9128 -4716 9146 -4710
rect 9156 -4744 9202 -4710
rect 9212 -4716 9230 -4710
rect 9786 -4716 9804 -4710
rect 9814 -4744 9860 -4710
rect 9870 -4716 9888 -4710
rect 10444 -4716 10462 -4710
rect 10472 -4744 10518 -4710
rect 10528 -4716 10546 -4710
rect 11102 -4716 11120 -4710
rect 11130 -4744 11176 -4710
rect 11186 -4716 11204 -4710
rect 11760 -4716 11778 -4710
rect 11788 -4744 11828 -4710
rect 9162 -4778 9196 -4744
rect 9820 -4778 9854 -4744
rect 10478 -4778 10512 -4744
rect 11136 -4778 11170 -4744
rect 11794 -4778 11828 -4744
rect 8390 -4812 11862 -4778
rect 8390 -5228 8424 -4812
rect 8504 -5228 8549 -4812
rect 8832 -5228 8877 -4812
rect 8946 -5228 8980 -4812
rect 9162 -5228 9196 -4812
rect 5392 -5302 9452 -5228
rect 5392 -5622 9536 -5302
rect 5392 -6122 9452 -5622
rect 5392 -6146 6907 -6122
rect 8390 -7370 8424 -6122
rect 8504 -7280 8538 -6122
rect 9162 -7280 9196 -6122
rect 11908 -7370 11942 -3686
rect 12362 -3940 12396 -3650
rect 12464 -3675 12522 -3653
rect 12592 -3675 12650 -3653
rect 12718 -3940 12752 -3650
rect 12496 -3988 12616 -3968
rect 12802 -3986 13042 -3686
rect 12802 -3988 13092 -3986
rect 12490 -4016 12644 -3996
rect 12802 -4014 13042 -3988
rect 12802 -4016 13120 -4014
rect 12802 -4072 13042 -4016
rect 13431 -4072 13518 -3272
rect 13467 -5834 13501 -4072
rect 13581 -4665 13615 -3272
rect 13581 -4767 13621 -4665
rect 13631 -4699 13649 -4693
rect 13943 -4699 13977 -1534
rect 14057 -1874 14102 -1534
rect 14118 -1874 14146 -1534
rect 14239 -1874 14284 -1534
rect 14715 -1874 14760 -590
rect 14776 -1874 14804 -586
rect 14832 -1874 14860 -586
rect 14897 -1874 14942 -586
rect 14952 -910 15334 -586
rect 14952 -918 15164 -910
rect 15373 -1062 15418 -586
rect 15373 -1874 15407 -1062
rect 15438 -1874 15466 -586
rect 15494 -1874 15522 -586
rect 15534 -606 15810 -586
rect 15555 -910 15810 -606
rect 15818 -550 16106 -470
rect 16108 -550 16136 2
rect 16164 -389 16247 2
rect 16164 -550 16192 -389
rect 16213 -448 16247 -389
rect 16689 -401 16723 2
rect 16677 -448 16735 -401
rect 16760 -442 16788 2
rect 16816 -172 16905 2
rect 16816 -392 16926 -172
rect 16816 -401 16844 -392
rect 16856 -401 16926 -392
rect 16816 -448 16926 -401
rect 16985 -448 17019 2
rect 17347 -401 17381 2
rect 17335 -448 17393 -401
rect 16213 -482 17393 -448
rect 16213 -530 16247 -482
rect 16213 -550 16258 -530
rect 16294 -550 16676 -482
rect 16677 -498 16735 -482
rect 16689 -530 16723 -498
rect 16689 -550 16734 -530
rect 16816 -550 16844 -488
rect 16856 -550 16926 -482
rect 16940 -550 17152 -482
rect 17335 -498 17393 -482
rect 17264 -538 17278 -532
rect 17304 -538 17306 -504
rect 17347 -513 17393 -498
rect 17461 -439 17495 2
rect 17502 -405 17529 2
rect 17461 -482 17490 -439
rect 17264 -544 17304 -538
rect 17347 -550 17381 -513
rect 17461 -538 17495 -482
rect 17538 -532 17542 -488
rect 17432 -544 17542 -538
rect 17461 -550 17495 -544
rect 15818 -584 17554 -550
rect 17696 -560 17704 2
rect 18136 -28 21794 6
rect 18136 -96 18376 -28
rect 18386 -96 18433 -49
rect 18136 -130 18433 -96
rect 18136 -424 18376 -130
rect 18403 -189 18448 -178
rect 18414 -365 18448 -189
rect 18386 -424 18433 -377
rect 18136 -450 18433 -424
rect 18502 -450 21794 -28
rect 18136 -484 21794 -450
rect 17832 -512 17952 -510
rect 18136 -526 18376 -484
rect 18502 -526 21794 -484
rect 18136 -530 21794 -526
rect 21806 -530 21828 746
rect 17804 -540 17980 -538
rect 15818 -606 16080 -584
rect 15555 -1062 15600 -910
rect 15818 -918 16030 -606
rect 16031 -1062 16076 -606
rect 15555 -1874 15589 -1062
rect 13986 -1908 15589 -1874
rect 13986 -3206 14020 -1908
rect 14057 -1914 14102 -1908
rect 14118 -1914 14146 -1908
rect 14057 -1929 14146 -1914
rect 14239 -1929 14284 -1908
rect 14715 -1914 14760 -1908
rect 14776 -1914 14804 -1908
rect 14715 -1929 14804 -1914
rect 14832 -1929 14860 -1908
rect 14897 -1929 14942 -1908
rect 14057 -1948 15190 -1929
rect 14057 -2058 14091 -1948
rect 14094 -1970 15190 -1948
rect 14100 -1976 14760 -1970
rect 14773 -1976 15190 -1970
rect 15373 -1976 15407 -1908
rect 14100 -2016 14146 -1976
rect 14150 -2010 14760 -1976
rect 14150 -2016 14174 -2010
rect 14094 -2058 14146 -2016
rect 14057 -2060 14146 -2058
rect 14057 -2069 14164 -2060
rect 14057 -3184 14091 -2069
rect 14100 -2300 14164 -2069
rect 14100 -3045 14146 -2300
rect 14174 -2328 14192 -2032
rect 14239 -2090 14284 -2010
rect 14715 -2016 14760 -2010
rect 14780 -2016 14804 -1976
rect 14808 -2010 15407 -1976
rect 14808 -2016 14860 -2010
rect 14715 -2090 14804 -2016
rect 14094 -3098 14146 -3045
rect 14122 -3144 14146 -3098
rect 14150 -3104 14174 -3098
rect 14239 -3104 14273 -2090
rect 14715 -3104 14749 -2090
rect 14758 -2784 14804 -2090
rect 14832 -2728 14860 -2016
rect 14897 -2090 14942 -2010
rect 15373 -2058 15407 -2010
rect 15438 -2053 15466 -1908
rect 15416 -2058 15466 -2053
rect 15373 -2060 15466 -2058
rect 15494 -2004 15522 -1908
rect 15530 -2004 15589 -1908
rect 15494 -2060 15589 -2004
rect 15373 -2069 15488 -2060
rect 14832 -2784 14876 -2728
rect 14758 -3045 14820 -2784
rect 14752 -3052 14820 -3045
rect 14832 -3052 14848 -2784
rect 14752 -3098 14804 -3052
rect 14832 -3098 14876 -3052
rect 14150 -3138 14749 -3104
rect 14150 -3144 14174 -3138
rect 14094 -3184 14146 -3144
rect 14057 -3200 14146 -3184
rect 14057 -3206 14102 -3200
rect 14118 -3206 14146 -3200
rect 14239 -3184 14273 -3138
rect 14276 -3184 14688 -3138
rect 14239 -3206 14688 -3184
rect 14715 -3184 14749 -3138
rect 14780 -3144 14804 -3098
rect 14808 -3104 14876 -3098
rect 14897 -3104 14931 -2090
rect 15373 -3104 15407 -2069
rect 15416 -2408 15488 -2069
rect 15494 -2408 15516 -2060
rect 15530 -2408 15589 -2060
rect 15416 -3061 15466 -2408
rect 14808 -3138 15407 -3104
rect 14808 -3144 14860 -3138
rect 14752 -3184 14804 -3144
rect 14715 -3200 14804 -3184
rect 14715 -3206 14760 -3200
rect 14776 -3206 14804 -3200
rect 14832 -3206 14860 -3144
rect 14897 -3184 14931 -3138
rect 14897 -3206 14942 -3184
rect 14952 -3206 15334 -3138
rect 15373 -3184 15407 -3138
rect 15373 -3206 15418 -3184
rect 15438 -3206 15466 -3061
rect 15494 -2464 15589 -2408
rect 15494 -3206 15522 -2464
rect 15530 -3184 15589 -2464
rect 15806 -3124 15810 -3116
rect 15530 -3206 15600 -3184
rect 13986 -3240 15600 -3206
rect 14057 -3716 14102 -3240
rect 14057 -4652 14091 -3716
rect 14045 -4699 14104 -4652
rect 14118 -4693 14146 -3240
rect 14239 -3564 14688 -3240
rect 14239 -3716 14284 -3564
rect 14476 -3572 14688 -3564
rect 14715 -3716 14760 -3240
rect 14239 -4652 14273 -3716
rect 14715 -4652 14749 -3716
rect 14239 -4699 14286 -4652
rect 14703 -4699 14762 -4652
rect 14776 -4693 14804 -3240
rect 14832 -4693 14860 -3240
rect 14897 -3716 14942 -3240
rect 14952 -3564 15334 -3240
rect 14952 -3572 15164 -3564
rect 15373 -3716 15418 -3240
rect 14897 -4652 14931 -3716
rect 15373 -4652 15407 -3716
rect 14897 -4699 14944 -4652
rect 15361 -4699 15420 -4652
rect 15438 -4693 15466 -3240
rect 15494 -4693 15522 -3240
rect 15555 -3716 15600 -3240
rect 15818 -3564 15822 -3124
rect 16031 -3184 16065 -1062
rect 16108 -1872 16136 -584
rect 16164 -1872 16192 -584
rect 16213 -1062 16258 -584
rect 16294 -918 16676 -584
rect 16689 -1062 16734 -584
rect 16213 -1872 16247 -1062
rect 16689 -1872 16723 -1062
rect 16816 -1872 16844 -584
rect 16856 -628 16926 -584
rect 16871 -1062 16916 -628
rect 16940 -694 17238 -584
rect 16940 -918 17152 -694
rect 17276 -732 17278 -724
rect 17304 -760 17306 -724
rect 16871 -1872 16905 -1062
rect 16985 -1872 17019 -918
rect 17347 -1872 17381 -584
rect 17461 -1872 17495 -584
rect 18136 -586 21805 -530
rect 18136 -596 18376 -586
rect 18176 -610 18210 -596
rect 18502 -610 21805 -586
rect 17682 -620 17686 -610
rect 17856 -790 17932 -788
rect 17828 -818 17960 -816
rect 17838 -1040 17948 -1020
rect 17876 -1078 17910 -1058
rect 18158 -1062 21805 -610
rect 18158 -1230 21794 -1062
rect 16072 -1906 17554 -1872
rect 16072 -3184 16106 -1906
rect 16108 -2060 16136 -1906
rect 16164 -2056 16192 -1906
rect 16213 -1974 16247 -1906
rect 16689 -1974 16723 -1906
rect 16816 -1927 16844 -1906
rect 16816 -1974 16863 -1927
rect 16213 -2008 16863 -1974
rect 16871 -1974 16905 -1906
rect 16985 -1974 17019 -1906
rect 17347 -1943 17381 -1906
rect 17347 -1958 17393 -1943
rect 17335 -1974 17393 -1958
rect 16871 -2008 17393 -1974
rect 16213 -2056 16247 -2008
rect 16164 -2060 16247 -2056
rect 16175 -2067 16247 -2060
rect 16186 -2316 16247 -2067
rect 16031 -3204 16106 -3184
rect 16108 -3204 16136 -2316
rect 16164 -3043 16247 -2316
rect 16164 -3204 16192 -3043
rect 16213 -3102 16247 -3043
rect 16689 -3102 16723 -2008
rect 16760 -3096 16788 -2014
rect 16816 -2056 16844 -2014
rect 16871 -2056 16905 -2008
rect 16816 -3043 16905 -2056
rect 16816 -3055 16844 -3043
rect 16816 -3102 16863 -3055
rect 16213 -3136 16863 -3102
rect 16871 -3102 16905 -3043
rect 16985 -3102 17019 -2008
rect 17335 -2055 17393 -2008
rect 17461 -1974 17495 -1906
rect 17461 -2017 17490 -1974
rect 17347 -3055 17381 -2055
rect 17335 -3102 17393 -3055
rect 16871 -3136 17393 -3102
rect 16213 -3184 16247 -3136
rect 16213 -3204 16258 -3184
rect 16294 -3204 16676 -3136
rect 16689 -3184 16723 -3136
rect 16689 -3204 16734 -3184
rect 16816 -3204 16844 -3142
rect 16871 -3184 16905 -3136
rect 16871 -3204 16916 -3184
rect 16940 -3204 17152 -3136
rect 17335 -3152 17393 -3136
rect 17347 -3167 17393 -3152
rect 17461 -3093 17495 -2017
rect 17502 -3059 17529 -2051
rect 17674 -2230 17686 -1974
rect 17702 -2176 17742 -1944
rect 18176 -2176 18210 -1230
rect 18290 -1312 18396 -1230
rect 18290 -2176 18324 -1312
rect 18502 -2176 21794 -1230
rect 17702 -2202 21794 -2176
rect 18176 -2358 18210 -2202
rect 18290 -2358 18324 -2202
rect 17642 -2648 17650 -2594
rect 18140 -2612 18376 -2358
rect 18136 -2648 18376 -2612
rect 18502 -2648 21794 -2202
rect 17461 -3136 17490 -3093
rect 17264 -3192 17278 -3186
rect 17264 -3198 17341 -3192
rect 17347 -3204 17381 -3167
rect 17461 -3192 17495 -3136
rect 17538 -3186 17542 -3142
rect 17387 -3198 17542 -3192
rect 17461 -3204 17495 -3198
rect 16031 -3238 17554 -3204
rect 17696 -3214 17704 -2648
rect 18136 -2682 21794 -2648
rect 18136 -2750 18376 -2682
rect 18386 -2750 18433 -2703
rect 18136 -2784 18433 -2750
rect 18136 -3031 18376 -2784
rect 18403 -2843 18448 -2832
rect 18414 -3019 18448 -2843
rect 18136 -3057 18433 -3031
rect 18136 -3078 18376 -3057
rect 18136 -3104 18386 -3078
rect 18502 -3104 21794 -2682
rect 18136 -3138 21794 -3104
rect 17832 -3166 17952 -3164
rect 18136 -3180 18376 -3138
rect 18426 -3166 18428 -3146
rect 18426 -3180 18434 -3174
rect 17804 -3194 17980 -3192
rect 18136 -3206 18466 -3180
rect 18502 -3184 21794 -3138
rect 21806 -3184 21828 -1062
rect 18502 -3206 21805 -3184
rect 16031 -3716 16076 -3238
rect 15555 -4652 15589 -3716
rect 16031 -4652 16065 -3716
rect 15555 -4699 15602 -4652
rect 16019 -4699 16078 -4652
rect 16108 -4693 16136 -3238
rect 16164 -4693 16192 -3238
rect 16213 -3716 16258 -3238
rect 16294 -3290 16676 -3238
rect 16689 -3290 16734 -3238
rect 16294 -3572 16742 -3290
rect 16213 -4652 16247 -3716
rect 16668 -3944 16742 -3572
rect 16689 -4652 16723 -3944
rect 16213 -4699 16260 -4652
rect 16677 -4699 16736 -4652
rect 16816 -4693 16844 -3238
rect 16871 -3716 16916 -3238
rect 16940 -3348 17238 -3238
rect 16940 -3572 17152 -3348
rect 16871 -4652 16905 -3716
rect 16871 -4699 16918 -4652
rect 16985 -4699 17019 -3572
rect 17347 -4652 17381 -3238
rect 17319 -4693 17381 -4652
rect 17313 -4699 17381 -4693
rect 13627 -4733 17381 -4699
rect 13631 -4739 13649 -4733
rect 13581 -4801 13615 -4767
rect 13943 -4801 13977 -4733
rect 14045 -4749 14103 -4733
rect 14057 -4801 14091 -4749
rect 14118 -4801 14146 -4739
rect 14239 -4801 14273 -4733
rect 14703 -4749 14761 -4733
rect 14715 -4801 14749 -4749
rect 14776 -4801 14804 -4739
rect 14832 -4801 14860 -4739
rect 14897 -4801 14931 -4733
rect 15361 -4749 15419 -4733
rect 15373 -4801 15407 -4749
rect 15438 -4801 15466 -4739
rect 15494 -4801 15522 -4739
rect 15555 -4801 15589 -4733
rect 16019 -4749 16077 -4733
rect 16031 -4801 16065 -4749
rect 16108 -4801 16136 -4739
rect 16164 -4801 16192 -4739
rect 16213 -4801 16247 -4733
rect 16677 -4749 16735 -4733
rect 16689 -4801 16723 -4749
rect 16816 -4801 16844 -4739
rect 16871 -4801 16905 -4733
rect 16985 -4801 17019 -4733
rect 17313 -4739 17331 -4733
rect 17341 -4767 17381 -4733
rect 17347 -4801 17381 -4767
rect 13563 -4835 17393 -4801
rect 17399 -4835 17415 -4801
rect 12496 -6642 12616 -6622
rect 12802 -6640 13042 -6088
rect 12802 -6642 13092 -6640
rect 12490 -6670 12644 -6650
rect 12802 -6668 13042 -6642
rect 12802 -6670 13120 -6668
rect 12802 -6726 13042 -6670
rect 13431 -6726 13518 -5834
rect 13467 -7393 13501 -6726
rect 13943 -7353 13977 -4835
rect 14057 -7294 14091 -4835
rect 14118 -5180 14146 -4835
rect 14118 -7347 14146 -6368
rect 14239 -7294 14273 -4835
rect 14715 -7294 14749 -4835
rect 14776 -5180 14804 -4835
rect 14832 -5180 14860 -4835
rect 14776 -7347 14804 -6368
rect 14832 -7347 14860 -6368
rect 14897 -7294 14931 -4835
rect 15373 -7294 15407 -4835
rect 15438 -5180 15466 -4835
rect 15494 -5180 15522 -4835
rect 15438 -7347 15466 -6368
rect 15494 -7347 15522 -6368
rect 15555 -7294 15589 -4835
rect 16031 -7294 16065 -4835
rect 16108 -5180 16136 -4835
rect 16164 -5180 16192 -4835
rect 16108 -7347 16136 -6368
rect 16164 -7347 16192 -6368
rect 16213 -7294 16247 -4835
rect 16689 -7294 16723 -4835
rect 16816 -5180 16844 -4835
rect 16816 -7347 16844 -6368
rect 16871 -7294 16905 -4835
rect 16985 -7353 17019 -4835
rect 13943 -7387 17019 -7353
rect 13943 -7403 13977 -7387
rect 14118 -7400 14146 -7393
rect 14776 -7400 14804 -7393
rect 14832 -7400 14860 -7393
rect 15438 -7400 15466 -7393
rect 15494 -7400 15522 -7393
rect 16108 -7400 16136 -7393
rect 16164 -7400 16192 -7393
rect 16816 -7400 16844 -7393
rect 13943 -7414 13954 -7403
rect 13966 -7414 13977 -7403
rect 16985 -7403 17019 -7387
rect 17461 -7393 17495 -3238
rect 18136 -3240 21805 -3206
rect 18136 -3250 18376 -3240
rect 18502 -3264 21805 -3240
rect 17682 -3274 17686 -3264
rect 18158 -3276 21805 -3264
rect 18538 -3396 18572 -3276
rect 17856 -3444 17932 -3442
rect 17828 -3472 17960 -3470
rect 17798 -3600 18070 -3480
rect 17748 -3694 18070 -3600
rect 17876 -3732 17910 -3712
rect 18510 -3752 18572 -3396
rect 18538 -7370 18572 -3752
rect 18652 -4642 18686 -3276
rect 18718 -3476 18724 -3374
rect 18746 -3448 18752 -3374
rect 18652 -4744 18692 -4642
rect 18702 -4676 18720 -4670
rect 19014 -4676 19048 -3276
rect 19112 -3592 19120 -3276
rect 19128 -3716 19173 -3276
rect 19204 -3648 19232 -3448
rect 19310 -3716 19355 -3276
rect 19372 -3592 19774 -3276
rect 19562 -3596 19774 -3592
rect 19786 -3716 19831 -3276
rect 19128 -4638 19162 -3716
rect 19116 -4676 19174 -4638
rect 19204 -4670 19232 -3848
rect 19310 -4638 19344 -3716
rect 19786 -4638 19820 -3716
rect 19310 -4676 19348 -4638
rect 19774 -4676 19832 -4638
rect 19856 -4670 19884 -3276
rect 19912 -4670 19940 -3276
rect 19968 -3716 20013 -3276
rect 20160 -3592 20422 -3276
rect 20426 -3592 20434 -3282
rect 20160 -3596 20250 -3592
rect 20444 -3716 20489 -3276
rect 19968 -4638 20002 -3716
rect 20444 -4638 20478 -3716
rect 19968 -4676 20006 -4638
rect 20432 -4676 20490 -4638
rect 20514 -4670 20542 -3276
rect 20570 -4670 20598 -3276
rect 20626 -3716 20671 -3276
rect 20686 -3592 21090 -3276
rect 20878 -3598 21090 -3592
rect 21102 -3716 21147 -3276
rect 20626 -4638 20660 -3716
rect 21102 -4638 21136 -3716
rect 20626 -4676 20664 -4638
rect 21090 -4676 21148 -4638
rect 21178 -4670 21206 -3276
rect 21234 -4670 21262 -3276
rect 21284 -3716 21329 -3276
rect 21354 -3598 21734 -3276
rect 21522 -3610 21734 -3598
rect 21742 -3610 21746 -3290
rect 21760 -3716 21805 -3276
rect 21284 -4638 21318 -3716
rect 21760 -4638 21794 -3716
rect 21806 -3752 21828 -3716
rect 21284 -4676 21322 -4638
rect 21748 -4676 21806 -4638
rect 21886 -4670 21914 600
rect 21942 -274 21987 746
rect 21918 -508 22010 -274
rect 22056 -508 22090 746
rect 21918 -732 22210 -508
rect 21942 -3752 21987 -732
rect 21998 -956 22210 -732
rect 21942 -4638 21976 -3752
rect 21942 -4676 21980 -4638
rect 22056 -4676 22090 -956
rect 22418 -4638 22452 746
rect 22532 0 22566 2097
rect 23615 -3180 23649 3435
rect 23779 3402 23782 3422
rect 24334 3402 27958 3497
rect 28438 3467 28636 3497
rect 28650 3467 30023 3497
rect 28342 3464 30023 3467
rect 28342 3436 28376 3464
rect 28308 3429 28410 3436
rect 28600 3435 28620 3464
rect 23751 3368 23754 3394
rect 23779 3389 23846 3402
rect 24294 3389 27958 3402
rect 24334 2120 27958 3389
rect 28342 2966 28376 3429
rect 28480 3395 28495 3429
rect 28511 3396 28536 3429
rect 28538 3396 28569 3429
rect 28518 3386 28533 3396
rect 28547 3386 28556 3396
rect 28585 3395 28594 3429
rect 28650 3402 30023 3464
rect 31220 3434 31254 3502
rect 31334 3472 31368 3502
rect 31372 3472 32884 3502
rect 31322 3434 32946 3472
rect 32960 3434 33498 3472
rect 33566 3468 33604 3472
rect 33566 3434 33606 3468
rect 30836 3402 32946 3434
rect 28620 3389 30023 3402
rect 30032 3394 30100 3402
rect 30166 3394 30242 3402
rect 30690 3394 30758 3402
rect 30824 3400 32946 3402
rect 32998 3400 33606 3434
rect 30824 3394 30906 3400
rect 28502 3362 28572 3386
rect 28523 3348 28557 3352
rect 28489 3314 28490 3319
rect 28511 3315 28569 3348
rect 28600 3346 28620 3389
rect 28445 3303 28490 3314
rect 28456 3127 28490 3303
rect 28489 3111 28490 3127
rect 28523 3115 28557 3315
rect 28584 3314 28591 3319
rect 28573 3303 28618 3314
rect 28584 3127 28618 3303
rect 28511 3102 28570 3115
rect 28584 3111 28591 3127
rect 28511 3034 28590 3102
rect 28511 3018 28569 3034
rect 28523 2966 28557 3000
rect 28650 2966 30023 3389
rect 28342 2932 30023 2966
rect 28650 2882 30023 2932
rect 28324 2262 30023 2882
rect 30690 2392 30826 2502
rect 30690 2366 30842 2392
rect 25045 1666 25079 2120
rect 25045 1346 25516 1666
rect 25045 877 25079 1346
rect 26361 877 26395 2120
rect 26435 877 26469 2120
rect 26549 877 26594 2120
rect 27019 877 27064 2120
rect 27133 1788 27170 2120
rect 27133 877 27167 1788
rect 27831 1350 27846 1560
rect 27859 1322 27874 1588
rect 27831 877 27846 1242
rect 27859 877 27902 1298
rect 28523 877 28557 2262
rect 28600 1696 28602 2120
rect 28650 882 30023 2262
rect 30750 1934 30842 2366
rect 31220 2176 31254 3400
rect 31322 3362 32896 3400
rect 33510 3394 33578 3400
rect 33602 3366 33606 3400
rect 33608 3450 33642 3502
rect 34246 3472 34250 3496
rect 33608 3402 33654 3450
rect 34224 3434 34262 3472
rect 34366 3450 34404 3472
rect 34354 3434 34412 3450
rect 34882 3434 34920 3472
rect 33656 3402 34262 3434
rect 34314 3402 34920 3434
rect 33608 3400 34262 3402
rect 34302 3400 34920 3402
rect 33608 3394 33726 3400
rect 34302 3394 34322 3400
rect 33608 3362 33654 3394
rect 34354 3362 34412 3400
rect 31334 3238 32895 3362
rect 32925 3350 32981 3361
rect 33583 3350 33596 3361
rect 33608 3350 33642 3362
rect 34266 3361 34292 3362
rect 34241 3350 34292 3361
rect 31296 3230 32895 3238
rect 31296 3090 32928 3230
rect 31334 3082 32928 3090
rect 31334 2328 32895 3082
rect 31372 2316 32854 2328
rect 32936 2316 32981 3350
rect 33594 2328 33642 3350
rect 34252 3346 34292 3350
rect 33594 2316 33628 2328
rect 34252 2316 34286 3346
rect 34366 2328 34400 3362
rect 34899 3350 34944 3361
rect 34910 2316 34944 3350
rect 31358 2278 32860 2316
rect 32874 2278 33498 2316
rect 33580 2278 33628 2316
rect 34240 2278 34298 2316
rect 34338 2278 34376 2316
rect 34898 2278 34956 2316
rect 31372 2244 32860 2278
rect 32912 2244 33628 2278
rect 33654 2244 33662 2278
rect 33670 2244 34376 2278
rect 34428 2244 34956 2278
rect 31372 2176 32854 2244
rect 32924 2228 32982 2244
rect 33582 2228 33628 2244
rect 34240 2228 34298 2244
rect 34898 2228 34956 2244
rect 32936 2176 32970 2210
rect 33594 2176 33628 2228
rect 34941 2213 34956 2228
rect 34252 2176 34286 2210
rect 34910 2176 34944 2210
rect 35024 2176 35058 3502
rect 35595 2176 39219 3567
rect 39672 2328 39706 5100
rect 41188 3536 41222 5108
rect 41882 3546 41916 5886
rect 41946 3556 41950 5886
rect 41958 4812 41980 5886
rect 41996 4812 42041 5886
rect 42654 4812 42692 5886
rect 42700 4812 42749 5886
rect 41958 3918 41986 4812
rect 41990 4344 42041 4812
rect 41990 3918 42030 4344
rect 42648 3952 42694 4812
rect 42698 4344 42749 4812
rect 43312 5490 43357 5886
rect 43462 5490 43507 5886
rect 43642 5490 43676 5886
rect 43744 5526 43816 5886
rect 43970 5509 44015 5886
rect 44220 5509 44265 5886
rect 44628 5509 44673 5886
rect 44978 5509 45023 5886
rect 45286 5509 45331 5886
rect 45400 5509 45434 5886
rect 45736 5511 45781 5886
rect 46494 5511 46539 5886
rect 47202 5726 47236 5886
rect 47252 5726 47297 5886
rect 47316 5878 47361 5886
rect 47974 5878 48055 5886
rect 47340 5828 47984 5866
rect 47378 5794 47984 5828
rect 48010 5726 48055 5878
rect 48088 5726 48122 5886
rect 47202 5692 48122 5726
rect 48392 5726 48426 5886
rect 48506 5878 48551 5886
rect 48768 5866 48813 5886
rect 49164 5878 49209 5886
rect 48530 5828 49174 5866
rect 48568 5794 49174 5828
rect 48756 5778 48814 5794
rect 48768 5726 48813 5778
rect 49278 5726 49312 5886
rect 48392 5692 49312 5726
rect 47252 5511 47297 5692
rect 48010 5511 48055 5692
rect 48658 5582 48716 5584
rect 48658 5526 48716 5556
rect 48768 5511 48813 5692
rect 48840 5582 48924 5584
rect 48840 5526 48924 5556
rect 49526 5511 49571 5886
rect 45724 5510 45725 5511
rect 45736 5510 45782 5511
rect 46482 5510 46483 5511
rect 46494 5510 46540 5511
rect 47240 5510 47241 5511
rect 47252 5510 47298 5511
rect 47998 5510 47999 5511
rect 48010 5510 48056 5511
rect 48756 5510 48757 5511
rect 48768 5510 48814 5511
rect 49514 5510 49515 5511
rect 49526 5510 49572 5511
rect 45723 5509 45724 5510
rect 43817 5498 45724 5509
rect 45736 5498 45770 5510
rect 45782 5509 45783 5510
rect 46481 5509 46482 5510
rect 45782 5498 46482 5509
rect 46494 5498 46528 5510
rect 46540 5509 46541 5510
rect 47239 5509 47240 5510
rect 46540 5498 47240 5509
rect 47252 5498 47286 5510
rect 47298 5509 47299 5510
rect 47997 5509 47998 5510
rect 47298 5498 47998 5509
rect 48010 5498 48044 5510
rect 48056 5509 48057 5510
rect 48755 5509 48756 5510
rect 48056 5498 48756 5509
rect 48768 5498 48802 5510
rect 48814 5509 48815 5510
rect 49513 5509 49514 5510
rect 48814 5498 49514 5509
rect 49526 5498 49560 5510
rect 49572 5509 49573 5510
rect 49702 5509 49736 5886
rect 49816 5509 49861 5886
rect 49885 5509 53509 5886
rect 49572 5498 53509 5509
rect 43828 5490 53509 5498
rect 43312 5464 53509 5490
rect 43312 5384 44064 5464
rect 44220 5384 44265 5464
rect 44628 5384 44673 5464
rect 44978 5384 45023 5464
rect 45286 5384 45331 5464
rect 45400 5384 45434 5464
rect 45736 5384 45770 5464
rect 46494 5384 46528 5464
rect 47252 5384 47286 5464
rect 48010 5384 48044 5464
rect 48768 5384 48802 5464
rect 49526 5384 49560 5464
rect 49702 5384 49736 5464
rect 49816 5384 49861 5464
rect 49885 5384 53509 5464
rect 43312 5350 53509 5384
rect 54074 5356 54108 5886
rect 43312 4932 44064 5350
rect 43312 4344 43357 4932
rect 42698 3952 42738 4344
rect 41958 3660 41980 3918
rect 41996 3698 42030 3918
rect 42654 3698 42688 3952
rect 41996 3682 42014 3698
rect 42670 3690 42688 3698
rect 42700 3690 42738 3952
rect 43312 3698 43346 4344
rect 42648 3686 42694 3690
rect 42698 3686 42738 3690
rect 43350 3686 43352 4344
rect 41962 3648 41980 3660
rect 42018 3580 42020 3682
rect 42046 3608 42048 3654
rect 42626 3648 42664 3686
rect 42670 3682 42688 3686
rect 42698 3682 42750 3686
rect 42682 3648 42750 3682
rect 43284 3648 43322 3686
rect 42058 3614 42664 3648
rect 42700 3614 43322 3648
rect 42700 3598 42750 3614
rect 43334 3608 43346 3682
rect 43406 3654 43408 4812
rect 43462 4344 43507 4932
rect 43970 4912 44015 4932
rect 44220 4912 44265 5350
rect 44628 4966 44673 5350
rect 44978 5262 45023 5350
rect 44978 5176 45076 5262
rect 44978 4966 45023 5176
rect 43784 4878 44332 4912
rect 43784 4596 43818 4878
rect 43970 4809 44015 4878
rect 43848 4754 43958 4792
rect 43886 4720 43958 4754
rect 43970 4764 44157 4809
rect 44220 4792 44265 4878
rect 43970 4721 44015 4764
rect 44158 4754 44265 4792
rect 43970 4676 44157 4721
rect 44196 4720 44265 4754
rect 43970 4596 44015 4676
rect 44220 4596 44265 4720
rect 44298 4596 44332 4878
rect 43784 4562 44332 4596
rect 44382 4786 45023 4966
rect 44382 4700 45076 4786
rect 43970 4436 44015 4562
rect 44220 4436 44265 4562
rect 44382 4504 45023 4700
rect 44422 4490 44744 4504
rect 44978 4490 45023 4504
rect 43784 4402 44332 4436
rect 43462 3686 43496 4344
rect 43784 4120 43818 4402
rect 43970 4356 44015 4402
rect 43920 4344 44196 4356
rect 44220 4344 44265 4402
rect 43970 4322 44004 4344
rect 44146 4322 44157 4333
rect 43954 4316 44162 4322
rect 44220 4316 44254 4344
rect 43848 4278 43920 4316
rect 43954 4312 44258 4316
rect 43954 4310 44264 4312
rect 43886 4244 43920 4278
rect 43970 4288 44157 4310
rect 43970 4234 44004 4288
rect 44158 4278 44264 4310
rect 44146 4234 44157 4245
rect 44196 4244 44264 4278
rect 43970 4200 44157 4234
rect 43970 4120 44004 4200
rect 44220 4120 44254 4244
rect 44298 4120 44332 4402
rect 43784 4086 44332 4120
rect 43970 3698 44004 4086
rect 44220 3686 44254 4086
rect 44382 4066 45023 4490
rect 45286 4344 45331 5350
rect 44382 4028 45020 4066
rect 44628 3698 44662 4028
rect 44978 3686 45012 4028
rect 45286 3698 45320 4344
rect 43362 3648 43408 3654
rect 43450 3648 43508 3686
rect 43942 3648 43980 3686
rect 44208 3648 44266 3686
rect 44600 3648 44638 3686
rect 44966 3648 45024 3686
rect 45258 3648 45296 3686
rect 43362 3614 43980 3648
rect 44032 3614 44638 3648
rect 44690 3614 45296 3648
rect 43362 3608 43402 3614
rect 43306 3552 43346 3608
rect 43450 3598 43508 3614
rect 44208 3598 44266 3614
rect 44966 3598 45024 3614
rect 43462 3546 43496 3598
rect 45400 3546 45434 5350
rect 41882 3536 45434 3546
rect 40702 3512 45434 3536
rect 40702 3502 44254 3512
rect 40702 2176 40736 3502
rect 41188 3472 41222 3502
rect 42080 3472 42104 3502
rect 43462 3472 43496 3502
rect 40840 3434 41484 3472
rect 41498 3434 42142 3472
rect 42156 3434 42800 3472
rect 42814 3434 43458 3472
rect 40878 3400 41484 3434
rect 41536 3400 42142 3434
rect 42194 3400 42800 3434
rect 41176 3362 41234 3400
rect 41934 3362 41992 3400
rect 42048 3394 42080 3400
rect 42692 3394 42774 3400
rect 42840 3394 42842 3402
rect 42852 3400 43458 3434
rect 43462 3400 44116 3472
rect 43370 3394 43420 3400
rect 40805 3350 40861 3361
rect 40816 3044 40861 3350
rect 41188 3044 41233 3362
rect 41463 3350 41519 3361
rect 41474 3044 41519 3350
rect 41946 3044 41991 3362
rect 42024 3346 42048 3394
rect 42080 3346 42104 3394
rect 42692 3362 42750 3394
rect 42121 3350 42177 3361
rect 42132 3044 42177 3350
rect 42704 3044 42749 3362
rect 42784 3361 42800 3362
rect 42814 3361 42830 3362
rect 42779 3350 42835 3361
rect 42784 3346 42835 3350
rect 42842 3346 42858 3390
rect 43364 3346 43370 3394
rect 43437 3350 43450 3361
rect 43462 3350 43838 3400
rect 44095 3350 44151 3361
rect 42790 3044 42835 3346
rect 43448 3258 43838 3350
rect 43424 3170 43838 3258
rect 43448 3044 43507 3170
rect 44106 3044 44151 3350
rect 40816 2316 40850 3044
rect 41188 2328 41222 3044
rect 41474 2316 41508 3044
rect 41946 2328 41980 3044
rect 42132 2316 42166 3044
rect 42704 2328 42738 3044
rect 42790 2316 42824 3044
rect 43448 2328 43496 3044
rect 43448 2316 43482 2328
rect 44106 2316 44140 3044
rect 40804 2278 40862 2316
rect 41160 2278 41198 2316
rect 41462 2278 41520 2316
rect 41918 2278 41956 2316
rect 42120 2278 42178 2316
rect 42676 2278 42714 2316
rect 42778 2278 42836 2316
rect 43434 2278 43482 2316
rect 44094 2278 44152 2316
rect 40804 2244 41198 2278
rect 41250 2244 41956 2278
rect 42008 2244 42714 2278
rect 42766 2244 43482 2278
rect 43508 2244 43516 2278
rect 43524 2244 44152 2278
rect 44186 2244 44208 2278
rect 40804 2228 40862 2244
rect 41462 2228 41520 2244
rect 42120 2228 42178 2244
rect 42778 2228 42836 2244
rect 43436 2228 43482 2244
rect 44094 2228 44152 2244
rect 40804 2213 40819 2228
rect 40816 2176 40850 2210
rect 41474 2176 41508 2210
rect 42132 2176 42166 2210
rect 42790 2176 42824 2210
rect 43448 2176 43482 2228
rect 44137 2213 44152 2228
rect 44106 2176 44140 2210
rect 44220 2176 44254 3502
rect 48768 2328 48802 5350
rect 49702 5134 49736 5350
rect 49816 5286 49861 5350
rect 49885 5274 53509 5350
rect 49840 5236 53509 5274
rect 49878 5202 53509 5236
rect 49885 5134 53509 5202
rect 49702 5100 53509 5134
rect 49885 4394 53509 5100
rect 54040 4572 54052 5356
rect 54068 4572 54108 5356
rect 53536 4402 53858 4406
rect 54074 4394 54108 4572
rect 54118 4394 54163 5886
rect 54172 5808 54206 5886
rect 54330 5876 54402 5886
rect 54488 5808 54522 5886
rect 54172 5774 54522 5808
rect 54776 5742 54820 5886
rect 54822 5742 54877 5886
rect 54764 5656 54877 5742
rect 54776 5596 54820 5656
rect 54166 4794 54186 4994
rect 54222 4884 54340 4954
rect 54222 4832 54646 4884
rect 54324 4394 54646 4832
rect 54686 4572 54738 5596
rect 54742 5356 54820 5596
rect 54742 4572 54766 5356
rect 54776 4394 54820 5356
rect 54822 4394 54877 5656
rect 54992 4394 55026 5886
rect 55106 4394 55151 5886
rect 55434 4394 55479 5886
rect 55548 4394 55582 5886
rect 55590 4394 55635 5886
rect 55666 4572 55686 5886
rect 55722 4572 55742 5886
rect 55764 4394 55809 5886
rect 56348 5364 56393 5886
rect 55816 4402 56066 4406
rect 49885 3500 56054 4394
rect 56314 4090 56338 5364
rect 44270 2278 44316 2284
rect 44266 2260 44316 2278
rect 44266 2244 44304 2260
rect 44270 2238 44304 2244
rect 49885 2176 53509 3500
rect 54002 3148 54016 3352
rect 54030 3120 54044 3352
rect 54074 2328 54108 3500
rect 54148 3166 54154 3352
rect 54176 3194 54182 3352
rect 54714 2284 54738 3352
rect 54742 2284 54766 3352
rect 54832 2328 54866 3500
rect 54854 2210 54880 2312
rect 54882 2238 54908 2284
rect 54992 2278 55026 3500
rect 55106 3044 55151 3500
rect 55590 3044 55635 3500
rect 55106 2342 55140 3044
rect 55590 2330 55624 3044
rect 55666 2342 55686 3352
rect 55722 2330 55742 3352
rect 55764 3044 55809 3500
rect 55764 2342 55798 3044
rect 56286 2576 56338 4090
rect 56314 2358 56338 2576
rect 56342 4344 56393 5364
rect 56422 4344 56467 5886
rect 56482 5308 56518 5886
rect 56342 4034 56388 4344
rect 56422 4034 56462 4344
rect 56482 4034 56490 5308
rect 57080 4344 57151 5886
rect 57316 4358 57638 4866
rect 56342 2632 56394 4034
rect 56422 2632 56456 4034
rect 56342 2330 56388 2632
rect 56422 2342 56462 2632
rect 56454 2330 56462 2342
rect 56482 2330 56490 2632
rect 57080 2342 57140 4344
rect 57376 4184 57528 4358
rect 57738 4344 57783 5886
rect 57864 4344 57909 5886
rect 57184 2540 57186 3930
rect 57212 2512 57214 3958
rect 57738 2342 57772 4344
rect 57802 2596 57810 3504
rect 57106 2330 57140 2342
rect 57864 2330 57898 4344
rect 55130 2316 55774 2330
rect 55788 2316 56432 2330
rect 56446 2316 57090 2330
rect 57106 2328 57748 2330
rect 57104 2326 57748 2328
rect 57102 2316 57748 2326
rect 57762 2316 57910 2330
rect 55590 2312 55624 2316
rect 55722 2298 55742 2316
rect 56348 2312 56382 2316
rect 56482 2302 56490 2316
rect 57106 2312 57140 2316
rect 57864 2312 57898 2316
rect 57126 2298 57136 2312
rect 56314 2292 56406 2298
rect 57126 2292 57174 2298
rect 57802 2292 57864 2298
rect 57978 2292 58012 5886
rect 58410 3567 58436 3894
rect 60069 3632 60103 6350
rect 60183 3698 60217 6350
rect 60164 3632 60238 3698
rect 55168 2278 55736 2292
rect 55826 2278 56428 2292
rect 56484 2278 57052 2292
rect 57126 2278 57710 2292
rect 57800 2278 58012 2292
rect 54992 2258 56394 2278
rect 54992 2244 55562 2258
rect 55652 2244 56320 2258
rect 56410 2244 57078 2278
rect 57092 2244 57094 2278
rect 54992 2228 55026 2244
rect 57126 2242 57136 2278
rect 57142 2258 58012 2278
rect 57168 2252 57836 2258
rect 57168 2244 57848 2252
rect 57808 2238 57848 2244
rect 57864 2240 57876 2252
rect 57978 2242 58012 2258
rect 57978 2231 57989 2242
rect 58001 2231 58012 2242
rect 58029 3531 58580 3567
rect 59108 3558 59194 3590
rect 60000 3558 60238 3632
rect 58772 3531 60254 3558
rect 60545 3531 60579 8088
rect 60659 7782 60704 8088
rect 60650 7748 60704 7782
rect 60720 7748 60748 8088
rect 60841 7748 60886 8088
rect 61317 7748 61362 8850
rect 61378 7748 61406 9624
rect 61434 7748 61462 9624
rect 61499 8850 61533 9624
rect 61499 7748 61544 8850
rect 61975 7748 62009 9624
rect 62040 7748 62068 9624
rect 62096 7748 62124 9624
rect 62157 7748 62191 9624
rect 60588 7714 62191 7748
rect 60588 6416 60622 7714
rect 60659 7708 60704 7714
rect 60720 7708 60748 7714
rect 60659 7693 60748 7708
rect 60841 7693 60886 7714
rect 61317 7708 61362 7714
rect 61378 7708 61406 7714
rect 61317 7693 61406 7708
rect 61434 7693 61462 7714
rect 61499 7693 61544 7714
rect 61975 7693 62009 7714
rect 60659 7652 61792 7693
rect 61975 7680 62022 7693
rect 61975 7662 62024 7680
rect 60659 7606 60704 7652
rect 60717 7646 61366 7652
rect 61375 7646 61792 7652
rect 61963 7646 62024 7662
rect 60724 7606 60748 7646
rect 60752 7612 61366 7646
rect 60752 7606 60776 7612
rect 60659 7562 60748 7606
rect 60659 7322 60766 7562
rect 60659 6565 60748 7322
rect 60776 7294 60794 7590
rect 60841 6565 60886 7612
rect 61305 7606 61362 7612
rect 61382 7606 61406 7646
rect 61410 7612 62024 7646
rect 61410 7606 61462 7612
rect 61305 7565 61406 7606
rect 61317 7532 61406 7565
rect 61317 6565 61351 7532
rect 61360 6838 61406 7532
rect 61434 6894 61462 7606
rect 61499 7532 61544 7612
rect 61963 7565 62009 7612
rect 62040 7569 62068 7714
rect 61975 7564 62009 7565
rect 62018 7564 62068 7569
rect 61975 7562 62068 7564
rect 62096 7618 62124 7714
rect 62132 7686 62191 7714
rect 62132 7618 62200 7686
rect 62096 7562 62200 7618
rect 61975 7553 62090 7562
rect 61434 6838 61478 6894
rect 61360 6577 61422 6838
rect 61354 6570 61422 6577
rect 61434 6570 61450 6838
rect 61354 6565 61406 6570
rect 60659 6524 60898 6565
rect 60659 6478 60704 6524
rect 60717 6518 60898 6524
rect 61305 6524 61406 6565
rect 61434 6524 61478 6570
rect 61305 6518 61366 6524
rect 60724 6478 60748 6518
rect 60752 6484 61366 6518
rect 60752 6478 60776 6484
rect 60659 6450 60748 6478
rect 60650 6422 60748 6450
rect 60650 6416 60704 6422
rect 60720 6416 60748 6422
rect 60841 6416 61290 6484
rect 61305 6468 61351 6484
rect 61382 6478 61406 6524
rect 61410 6518 61478 6524
rect 61499 6565 61533 7532
rect 61975 6565 62009 7553
rect 62018 7214 62090 7553
rect 62096 7214 62118 7562
rect 62132 7214 62200 7562
rect 62018 6565 62068 7214
rect 61499 6518 61546 6565
rect 61963 6561 62068 6565
rect 61963 6552 62022 6561
rect 61963 6518 62024 6552
rect 61410 6484 62024 6518
rect 61410 6478 61462 6484
rect 61317 6438 61351 6468
rect 61354 6438 61406 6478
rect 61317 6422 61406 6438
rect 61317 6416 61362 6422
rect 61378 6416 61406 6422
rect 61434 6416 61462 6478
rect 61499 6438 61533 6484
rect 61499 6416 61544 6438
rect 61554 6416 61936 6484
rect 61963 6468 62009 6484
rect 61975 6438 62009 6468
rect 61975 6416 62020 6438
rect 62040 6416 62068 6561
rect 62096 7158 62200 7214
rect 62096 6416 62124 7158
rect 62132 6478 62200 7158
rect 62408 6498 62412 6506
rect 62132 6438 62191 6478
rect 62132 6416 62202 6438
rect 60588 6382 62202 6416
rect 60659 3531 60704 6382
rect 60720 6000 60748 6382
rect 60841 6058 61290 6382
rect 60720 3531 60748 4812
rect 60776 3531 60804 3894
rect 60841 3531 60886 6058
rect 61078 6050 61290 6058
rect 61317 5906 61362 6382
rect 61378 6000 61406 6382
rect 61434 6000 61462 6382
rect 61499 5906 61544 6382
rect 61554 6058 61936 6382
rect 61554 6050 61766 6058
rect 61975 5906 62020 6382
rect 62040 6000 62068 6382
rect 62096 6000 62124 6382
rect 62157 5906 62202 6382
rect 62420 6058 62424 6498
rect 62633 6438 62667 9624
rect 62710 7750 62738 9624
rect 62766 7750 62794 9624
rect 62815 7750 62849 9624
rect 63291 7750 63325 9624
rect 63418 7750 63446 9624
rect 63473 7750 63507 9624
rect 63587 7750 63621 9624
rect 63949 7750 63983 7784
rect 64063 7750 64097 9624
rect 62674 7716 64156 7750
rect 62674 6438 62708 7716
rect 62710 7562 62738 7716
rect 62766 7566 62794 7716
rect 62815 7648 62849 7716
rect 63291 7695 63325 7716
rect 63418 7695 63446 7716
rect 63291 7664 63338 7695
rect 63279 7648 63338 7664
rect 63418 7648 63465 7695
rect 62815 7614 63465 7648
rect 63473 7648 63507 7716
rect 63587 7648 63621 7716
rect 63949 7664 63995 7695
rect 63937 7648 63995 7664
rect 63473 7614 63995 7648
rect 62815 7566 62849 7614
rect 63279 7567 63337 7614
rect 62766 7562 62849 7566
rect 62777 7555 62849 7562
rect 62788 7306 62849 7555
rect 62633 6418 62708 6438
rect 62710 6418 62738 7306
rect 62766 6579 62849 7306
rect 62766 6418 62794 6579
rect 62815 6520 62849 6579
rect 63291 6567 63325 7567
rect 63279 6520 63338 6567
rect 63362 6526 63390 7608
rect 63418 7566 63446 7608
rect 63473 7566 63507 7614
rect 63418 6579 63507 7566
rect 63418 6567 63446 6579
rect 63418 6520 63465 6567
rect 62815 6486 63465 6520
rect 63473 6520 63507 6579
rect 63587 6520 63621 7614
rect 63937 7567 63995 7614
rect 64063 7648 64097 7716
rect 64063 7605 64092 7648
rect 63949 6567 63983 7567
rect 63937 6520 63995 6567
rect 63473 6486 63995 6520
rect 64063 6529 64097 7605
rect 64104 6563 64131 7571
rect 64778 7264 64812 10652
rect 75116 10604 75150 11692
rect 75218 10684 75252 15472
rect 76128 10684 76162 15472
rect 76230 10604 76264 15472
rect 65550 10565 65584 10569
rect 65544 10540 65584 10565
rect 66208 10540 66242 10569
rect 66866 10540 66900 10569
rect 67524 10540 67558 10569
rect 68182 10540 68216 10569
rect 75116 10542 75150 10553
rect 76230 10542 76264 10558
rect 65104 10504 68366 10540
rect 75116 10535 76264 10542
rect 76574 10535 76608 15472
rect 77104 15152 77140 15160
rect 77186 15152 77204 15160
rect 75080 10504 76625 10535
rect 76688 10504 76722 10538
rect 77146 10504 77180 10538
rect 77260 10504 77294 15472
rect 83158 15436 86794 15484
rect 88271 15483 88305 15839
rect 88385 15644 88419 15839
rect 88431 15827 88432 15828
rect 89030 15827 89031 15828
rect 88430 15826 88431 15827
rect 89031 15826 89032 15827
rect 89043 15644 89077 15839
rect 89089 15827 89090 15828
rect 89688 15827 89689 15828
rect 89088 15826 89089 15827
rect 89689 15826 89690 15827
rect 89701 15644 89735 15839
rect 89747 15827 89748 15828
rect 90346 15827 90347 15828
rect 89746 15826 89747 15827
rect 90347 15826 90348 15827
rect 90359 15644 90393 15839
rect 90405 15827 90406 15828
rect 90404 15826 90405 15827
rect 90668 15811 90749 15858
rect 90668 15632 90669 15633
rect 89015 15585 89062 15632
rect 89673 15585 89720 15632
rect 90331 15585 90378 15632
rect 90667 15631 90668 15632
rect 90715 15585 90749 15811
rect 90817 15585 90851 17269
rect 88447 15551 89062 15585
rect 89105 15551 89720 15585
rect 89763 15551 90378 15585
rect 90421 15551 90851 15585
rect 90715 15483 90749 15551
rect 90817 15483 90851 15551
rect 91789 15545 91823 26373
rect 92066 25834 92113 26472
rect 92292 26436 92326 27762
rect 103078 27754 105218 27788
rect 95376 27328 95996 27750
rect 96046 27702 96612 27736
rect 96046 27380 96080 27702
rect 96417 27622 96428 27633
rect 96101 27560 96182 27607
rect 96241 27588 96428 27622
rect 96429 27560 96510 27607
rect 96148 27522 96182 27560
rect 96476 27522 96510 27560
rect 96417 27494 96428 27505
rect 96241 27460 96428 27494
rect 96578 27380 96612 27702
rect 103621 27570 103655 27754
rect 96046 27346 96612 27380
rect 95434 27274 95452 27313
rect 95752 27285 95782 27320
rect 95808 27285 95810 27320
rect 96424 27306 96944 27320
rect 95468 27274 95486 27279
rect 95782 27274 95808 27285
rect 95376 27228 95996 27274
rect 96108 27260 96550 27294
rect 96046 27233 96612 27260
rect 95376 27226 96056 27228
rect 95376 27212 96114 27226
rect 95376 27200 95996 27212
rect 95376 27198 96028 27200
rect 95376 27165 96086 27198
rect 95376 27131 100800 27165
rect 95376 27095 95996 27131
rect 96046 26998 96086 27131
rect 96094 27004 96114 27124
rect 96148 27097 96182 27100
rect 96476 27097 96510 27100
rect 96046 26966 96080 26998
rect 96578 26966 96612 27131
rect 103066 27095 103691 27570
rect 93306 26474 94648 26510
rect 95234 26504 95452 26508
rect 95888 26474 95922 26590
rect 96064 26550 100800 26584
rect 96012 26522 96070 26540
rect 96002 26512 96036 26516
rect 95952 26486 95996 26496
rect 96002 26494 96042 26512
rect 96002 26474 96036 26494
rect 96580 26486 96802 26508
rect 92406 26436 92430 26470
rect 93306 26450 96894 26474
rect 101174 26450 101208 26590
rect 103102 26450 103136 27095
rect 104446 27074 104466 27356
rect 93306 26440 103618 26450
rect 92198 26402 92492 26436
rect 92292 26368 92326 26402
rect 92292 26300 92350 26368
rect 92424 26340 92440 26374
rect 92292 26040 92326 26300
rect 92344 26065 92360 26241
rect 92368 26065 92378 26241
rect 92394 26078 92444 26307
rect 92394 26053 92452 26078
rect 92292 25972 92350 26040
rect 92292 25904 92326 25972
rect 92396 25904 92452 26053
rect 92458 25904 92492 26402
rect 92198 25870 92492 25904
rect 92578 26402 92968 26436
rect 92578 25904 92612 26402
rect 92792 26334 92839 26381
rect 92754 26300 92839 26334
rect 92681 26241 92726 26252
rect 92809 26241 92854 26252
rect 92692 26065 92726 26241
rect 92820 26065 92854 26241
rect 92792 26006 92839 26053
rect 92754 25972 92839 26006
rect 92934 25904 92968 26402
rect 92578 25870 92968 25904
rect 92292 25820 92326 25870
rect 92396 25868 92452 25870
rect 92332 25820 92452 25868
rect 92256 25456 92506 25820
rect 92560 25456 92982 25820
rect 93306 25456 94648 26440
rect 95366 26419 103618 26440
rect 95270 26416 103618 26419
rect 92562 25382 92594 25456
rect 92596 25382 92628 25456
rect 92710 25406 92744 25416
rect 92798 25406 92832 25416
rect 92676 25372 92866 25382
rect 92436 25270 92470 25282
rect 92214 25236 92470 25270
rect 92596 25270 92630 25282
rect 92912 25270 92946 25282
rect 92596 25236 92946 25270
rect 93342 25228 93376 25456
rect 93456 25228 93490 25262
rect 94114 25228 94148 25262
rect 94772 25228 94806 25262
rect 95270 25228 95304 26416
rect 95888 26372 95922 26416
rect 96002 26403 96040 26410
rect 95990 26388 96040 26403
rect 95990 26372 96048 26388
rect 96060 26372 96098 26410
rect 96718 26372 96756 26410
rect 95492 26370 96098 26372
rect 96150 26370 96756 26372
rect 95346 26332 95366 26340
rect 95406 26338 95418 26370
rect 95476 26348 96098 26370
rect 95461 26338 96098 26348
rect 96134 26340 96756 26370
rect 96860 26340 96894 26416
rect 96128 26338 96756 26340
rect 95412 26332 95414 26338
rect 95461 26336 96082 26338
rect 96128 26336 96214 26338
rect 96662 26336 96740 26338
rect 96786 26336 96944 26340
rect 101060 26336 101094 26416
rect 101174 26336 101208 26416
rect 103102 26336 103136 26416
rect 103216 26402 103250 26416
rect 103204 26360 103262 26402
rect 103216 26356 103250 26360
rect 103244 26348 103432 26356
rect 103244 26342 103444 26348
rect 103182 26336 103444 26342
rect 95338 26300 95346 26314
rect 95430 26304 101208 26336
rect 95430 26300 95440 26304
rect 95442 26300 95444 26304
rect 95456 26302 101208 26304
rect 103068 26302 103136 26336
rect 103178 26334 103444 26336
rect 103182 26322 103444 26334
rect 103240 26312 103444 26322
rect 103240 26302 103554 26312
rect 95470 26300 96082 26302
rect 95334 26286 95406 26300
rect 95424 26290 95440 26300
rect 95470 26296 95562 26300
rect 95476 26290 95477 26291
rect 95334 26284 95412 26286
rect 95334 26274 95406 26284
rect 95372 25706 95406 26274
rect 95396 25690 95406 25706
rect 95418 25690 95464 26290
rect 95475 26289 95476 26290
rect 95470 26268 95562 26284
rect 95475 25690 95476 25691
rect 95430 25678 95464 25690
rect 95476 25689 95477 25690
rect 95888 25678 95922 26300
rect 96002 25724 96036 26300
rect 96042 26299 96082 26300
rect 96042 26296 96122 26299
rect 96128 26296 96214 26302
rect 96662 26299 96740 26302
rect 96662 26296 96780 26299
rect 96786 26296 96944 26302
rect 96077 26288 96122 26296
rect 96735 26288 96780 26296
rect 96042 26268 96082 26284
rect 96088 25712 96122 26288
rect 96128 26268 96214 26284
rect 96662 26268 96740 26284
rect 96746 25712 96780 26288
rect 96860 26284 96894 26296
rect 101047 26290 101048 26291
rect 101048 26289 101049 26290
rect 96786 26268 96894 26284
rect 96860 25772 96894 26268
rect 96860 25770 96944 25772
rect 96002 25708 96036 25712
rect 96076 25708 96134 25712
rect 96734 25708 96792 25712
rect 96860 25708 96894 25770
rect 97072 25708 97112 25716
rect 97128 25708 97140 25744
rect 101060 25724 101094 26302
rect 101060 25708 101094 25712
rect 96030 25682 101066 25708
rect 96026 25678 101070 25682
rect 101174 25678 101208 26302
rect 103102 26220 103136 26302
rect 103262 26290 103554 26302
rect 103278 26288 103554 26290
rect 103482 26220 103516 26274
rect 103584 26220 103618 26416
rect 103102 26186 103926 26220
rect 103482 25726 103516 26186
rect 103584 25726 103618 26186
rect 106368 25980 106370 27368
rect 106344 25774 106370 25980
rect 106368 25768 106370 25774
rect 106694 26500 112614 29242
rect 113083 26500 113117 30798
rect 113197 30761 113244 30777
rect 113185 30696 113244 30761
rect 113855 30746 113902 30777
rect 114513 30746 114560 30777
rect 115171 30746 115218 30777
rect 113843 30730 113902 30746
rect 114501 30730 114560 30746
rect 115159 30730 115218 30746
rect 113294 30696 113902 30730
rect 113952 30696 114560 30730
rect 114610 30696 115218 30730
rect 113185 30687 113220 30696
rect 113843 30687 113878 30696
rect 114501 30687 114536 30696
rect 115159 30687 115194 30696
rect 113185 30649 113231 30687
rect 113136 26608 113162 26724
rect 113164 26649 113190 26696
rect 113197 26649 113231 30649
rect 113232 30648 113265 30653
rect 113843 30649 113889 30687
rect 113232 28284 113266 30648
rect 113232 26661 113277 28284
rect 113286 26652 113290 26864
rect 113314 26649 113318 26892
rect 113855 26649 113889 30649
rect 113890 30648 113923 30653
rect 114501 30649 114547 30687
rect 113890 28284 113924 30648
rect 114513 29606 114547 30649
rect 114479 28938 114490 29606
rect 114507 28938 114547 29606
rect 113890 26661 113935 28284
rect 114513 27750 114547 28938
rect 114479 26684 114490 27750
rect 114507 26684 114547 27750
rect 114513 26649 114547 26684
rect 114548 30648 114581 30653
rect 115159 30649 115205 30687
rect 114548 28284 114582 30648
rect 115137 28938 115140 29606
rect 115165 28938 115168 29606
rect 114548 26661 114593 28284
rect 114606 26654 114616 26862
rect 114634 26649 114644 26890
rect 115137 26649 115140 27750
rect 115165 26649 115168 27750
rect 115171 26649 115205 30649
rect 115206 30648 115239 30653
rect 115206 28284 115240 30648
rect 115206 26661 115251 28284
rect 113164 26608 113244 26649
rect 113185 26568 113244 26608
rect 113247 26602 113902 26649
rect 113905 26602 114560 26649
rect 114563 26602 115218 26649
rect 113185 26552 113220 26568
rect 113185 26537 113200 26552
rect 113254 26534 113272 26602
rect 113282 26568 113902 26602
rect 113952 26568 114560 26602
rect 113282 26562 113300 26568
rect 113843 26552 113878 26568
rect 114501 26552 114536 26568
rect 114570 26534 114580 26602
rect 114598 26562 114608 26602
rect 114610 26568 115218 26602
rect 115159 26552 115194 26568
rect 113197 26500 113231 26534
rect 113855 26500 113889 26534
rect 114513 26500 114547 26534
rect 115171 26500 115205 26534
rect 115320 26500 115354 30798
rect 106694 26469 115354 26500
rect 115829 26469 115863 31139
rect 115969 26469 116003 31139
rect 116083 28284 116117 31139
rect 116302 28996 116304 29152
rect 116487 28284 116521 31139
rect 116083 26469 116128 28284
rect 116487 26469 116532 28284
rect 116601 26469 116635 31139
rect 118019 29626 118034 29708
rect 117312 29582 117702 29616
rect 118057 29588 118072 29746
rect 116638 28938 116648 29134
rect 117312 29084 117346 29582
rect 117399 29421 117433 29582
rect 117526 29514 117573 29561
rect 117488 29480 117573 29514
rect 117445 29421 117460 29432
rect 117543 29421 117588 29432
rect 117399 29245 117460 29421
rect 117554 29245 117588 29421
rect 117399 29222 117433 29245
rect 117399 29084 117439 29222
rect 117448 29098 117467 29194
rect 117526 29186 117573 29233
rect 117488 29152 117573 29186
rect 117668 29084 117702 29582
rect 116694 28938 116704 29078
rect 117312 29050 117702 29084
rect 117298 28380 117720 29000
rect 118023 28938 118050 29090
rect 118051 28938 118078 29118
rect 117300 27408 117306 27664
rect 117328 27436 117334 27636
rect 106694 26466 116635 26469
rect 106694 26126 112614 26466
rect 113083 26373 113117 26466
rect 113165 26435 116635 26466
rect 106694 25906 112624 26126
rect 103404 25712 103796 25726
rect 103340 25700 103796 25712
rect 103404 25684 103796 25700
rect 104470 25690 105016 25726
rect 105566 25696 105892 25726
rect 106228 25696 106558 25726
rect 95430 25674 101128 25678
rect 95334 25616 95406 25654
rect 95430 25644 101070 25674
rect 101140 25644 101208 25678
rect 103312 25678 103796 25684
rect 103312 25672 103444 25678
rect 103584 25670 103618 25678
rect 95430 25632 95464 25644
rect 95476 25632 95477 25633
rect 95372 25596 95406 25616
rect 95418 25596 95464 25632
rect 95475 25631 95476 25632
rect 95372 25232 95475 25596
rect 95888 25572 95922 25644
rect 96064 25640 101070 25644
rect 96076 25624 96134 25640
rect 96734 25632 101048 25640
rect 96734 25624 96792 25632
rect 96088 25596 96122 25624
rect 96746 25596 96780 25624
rect 96088 25572 96133 25596
rect 96746 25572 96791 25596
rect 96860 25572 96894 25632
rect 97072 25608 97112 25632
rect 97128 25618 97140 25632
rect 101174 25572 101208 25644
rect 103404 25622 103852 25670
rect 104442 25662 105044 25670
rect 105538 25668 105892 25670
rect 106228 25668 106586 25670
rect 95888 25538 101208 25572
rect 95334 25228 95475 25232
rect 96088 25228 96133 25538
rect 96746 25228 96791 25538
rect 96860 25228 96894 25538
rect 92364 25194 102616 25228
rect 93342 25114 93376 25194
rect 93456 25114 93490 25194
rect 94114 25114 94148 25194
rect 94396 25114 94760 25125
rect 94772 25114 94806 25194
rect 95270 25125 95304 25194
rect 95372 25180 95475 25194
rect 96088 25180 96133 25194
rect 96746 25180 96791 25194
rect 94818 25114 95308 25125
rect 95372 25118 95406 25180
rect 95334 25114 95406 25118
rect 95418 25114 95464 25180
rect 96088 25114 96122 25180
rect 96746 25114 96780 25180
rect 96860 25114 96894 25194
rect 102582 25138 102616 25194
rect 102430 25114 102441 25125
rect 102442 25118 102616 25138
rect 93342 25080 102441 25114
rect 93342 24656 93376 25080
rect 93456 24656 93490 25080
rect 93502 25068 93503 25069
rect 94101 25068 94102 25069
rect 93501 25067 93502 25068
rect 94102 25067 94103 25068
rect 93501 24668 93502 24669
rect 94102 24668 94103 24669
rect 93502 24667 93503 24668
rect 94101 24667 94102 24668
rect 94114 24656 94148 25080
rect 94160 25068 94161 25069
rect 94759 25068 94760 25069
rect 94772 25068 94806 25080
rect 94818 25068 94819 25069
rect 94159 25067 94160 25068
rect 94760 25067 94761 25068
rect 94772 25067 94818 25068
rect 94772 24669 94817 25067
rect 94159 24668 94160 24669
rect 94760 24668 94761 24669
rect 94772 24668 94818 24669
rect 94160 24667 94161 24668
rect 94759 24667 94760 24668
rect 94208 24656 94760 24667
rect 94772 24656 94806 24668
rect 94818 24667 94819 24668
rect 95270 24667 95304 25080
rect 95372 25074 95406 25080
rect 95338 25008 95346 25074
rect 95366 25036 95406 25074
rect 95418 25068 95464 25080
rect 95390 25032 95406 25036
rect 95390 24996 95402 25032
rect 95430 25020 95464 25068
rect 95526 25020 95562 25026
rect 96010 25020 96082 25026
rect 96088 25020 96122 25080
rect 96128 25020 96214 25026
rect 96662 25020 96698 25026
rect 96746 25020 96780 25080
rect 96860 25026 96894 25080
rect 102442 25052 102514 25090
rect 102480 25032 102514 25052
rect 96834 25020 96944 25026
rect 102442 25020 102530 25032
rect 102582 25020 102616 25118
rect 95334 24958 95406 24996
rect 95372 24740 95406 24958
rect 94818 24656 95308 24667
rect 95332 24662 95346 24740
rect 95360 24662 95406 24740
rect 95430 24986 102530 25020
rect 102548 24986 102616 25020
rect 95430 24668 95464 24986
rect 95372 24660 95406 24662
rect 95334 24656 95406 24660
rect 95418 24656 95464 24668
rect 96088 24656 96122 24986
rect 96746 24656 96780 24986
rect 96860 24656 96894 24986
rect 102442 24974 102530 24986
rect 102480 24684 102514 24974
rect 102430 24656 102441 24667
rect 93342 24622 102441 24656
rect 93342 24542 93376 24622
rect 93456 24542 93490 24622
rect 94114 24542 94148 24622
rect 94772 24542 94806 24622
rect 95270 24542 95304 24622
rect 95372 24616 95406 24622
rect 95332 24546 95346 24616
rect 95360 24572 95406 24616
rect 95418 24572 95464 24622
rect 96088 24572 96122 24622
rect 96746 24572 96780 24622
rect 95360 24546 95475 24572
rect 95332 24542 95475 24546
rect 96088 24542 96133 24572
rect 96746 24542 96791 24572
rect 96860 24542 96894 24622
rect 102582 24542 102616 24986
rect 92364 24508 102616 24542
rect 92032 22400 92082 22406
rect 92088 22400 92110 22434
rect 92032 22206 92082 22214
rect 92088 22178 92110 22214
rect 92032 19746 92082 19752
rect 92088 19746 92110 19780
rect 92032 19552 92082 19560
rect 92088 19524 92110 19560
rect 93342 18262 93376 24508
rect 94772 24044 94806 24508
rect 94460 23820 94806 24044
rect 95270 23820 95304 24508
rect 95332 24426 95346 24508
rect 95360 24454 95475 24508
rect 95338 24350 95346 24426
rect 95366 24390 95475 24454
rect 95366 24378 95412 24390
rect 95418 24375 95475 24390
rect 96088 24375 96133 24508
rect 95418 24374 95476 24375
rect 96076 24374 96077 24375
rect 96088 24374 96134 24375
rect 96734 24374 96735 24375
rect 96746 24374 96791 24508
rect 95424 24362 95464 24374
rect 95476 24373 95477 24374
rect 96075 24373 96076 24374
rect 95476 24362 96076 24373
rect 96088 24362 96122 24374
rect 96134 24373 96135 24374
rect 96733 24373 96734 24374
rect 96134 24362 96734 24373
rect 96746 24362 96780 24374
rect 96860 24362 96894 24508
rect 95424 24350 96928 24362
rect 95430 24340 96928 24350
rect 95338 24338 95346 24340
rect 95424 24338 96928 24340
rect 95334 24328 96928 24338
rect 95334 24316 95464 24328
rect 95476 24316 95477 24317
rect 96075 24316 96076 24317
rect 96088 24316 96122 24328
rect 96134 24316 96135 24317
rect 96733 24316 96734 24317
rect 96746 24316 96780 24328
rect 95334 24315 95476 24316
rect 96076 24315 96077 24316
rect 96088 24315 96134 24316
rect 96734 24315 96735 24316
rect 95334 24300 95475 24315
rect 95338 23820 95346 24300
rect 95366 24244 95475 24300
rect 95366 23820 95498 24244
rect 96088 23820 96133 24315
rect 96746 23820 96791 24316
rect 96860 23820 96894 24328
rect 93444 23786 96894 23820
rect 93456 23756 93490 23786
rect 94114 23756 94148 23786
rect 94460 23756 94806 23786
rect 95270 23756 95304 23786
rect 95338 23756 95346 23786
rect 95366 23756 95475 23786
rect 96088 23756 96133 23786
rect 96746 23756 96791 23786
rect 93456 23718 96791 23756
rect 93456 18300 93490 23718
rect 93518 23684 94148 23718
rect 94176 23684 94806 23718
rect 94834 23717 95475 23718
rect 95480 23717 96133 23718
rect 94834 23716 95476 23717
rect 95480 23716 96134 23717
rect 96138 23716 96791 23718
rect 94834 23710 95470 23716
rect 95476 23715 95477 23716
rect 95480 23715 96128 23716
rect 95476 23710 96128 23715
rect 96134 23715 96135 23716
rect 96138 23715 96780 23716
rect 94834 23704 95464 23710
rect 95476 23704 96122 23710
rect 96134 23704 96780 23715
rect 96860 23704 96894 23786
rect 94834 23684 96894 23704
rect 94080 18300 94092 18418
rect 94114 18300 94148 23684
rect 94460 23602 94806 23684
rect 94772 18300 94806 23602
rect 95270 22932 95304 23684
rect 95396 23682 95414 23684
rect 95338 23680 95414 23682
rect 95424 23680 96894 23684
rect 95334 23670 96894 23680
rect 95334 23658 95464 23670
rect 95476 23658 95477 23659
rect 96075 23658 96076 23659
rect 96088 23658 96122 23670
rect 96134 23658 96135 23659
rect 96733 23658 96734 23659
rect 96746 23658 96780 23670
rect 95334 23657 95476 23658
rect 96076 23657 96077 23658
rect 96088 23657 96134 23658
rect 96734 23657 96735 23658
rect 95334 23642 95475 23657
rect 95338 23620 95346 23642
rect 95332 23116 95346 23620
rect 95366 23592 95475 23642
rect 95360 23550 95475 23592
rect 96088 23550 96133 23657
rect 96746 23550 96791 23658
rect 95360 23144 95406 23550
rect 95338 23034 95346 23116
rect 95366 23062 95412 23144
rect 95396 23058 95406 23062
rect 95418 23058 95464 23550
rect 95475 23058 95476 23059
rect 96076 23058 96077 23059
rect 95424 23052 95464 23058
rect 95476 23057 95477 23058
rect 96075 23057 96076 23058
rect 95390 23046 95464 23052
rect 96088 23046 96122 23550
rect 96133 23058 96134 23059
rect 96734 23058 96735 23059
rect 96134 23057 96135 23058
rect 96733 23057 96734 23058
rect 96746 23046 96780 23550
rect 96860 23046 96894 23670
rect 95390 23034 96894 23046
rect 95390 22932 95402 23034
rect 95430 23012 96894 23034
rect 95430 22932 95464 23012
rect 96088 22932 96122 23012
rect 96746 22932 96780 23012
rect 96860 22932 96894 23012
rect 103584 22994 103618 25622
rect 106694 25322 112614 25906
rect 106694 25306 112654 25322
rect 106694 25058 112614 25306
rect 112654 25242 112670 25306
rect 112902 25242 112906 25322
rect 106694 24955 112615 25058
rect 112653 24994 112654 24995
rect 112654 24993 112655 24994
rect 112668 24955 112695 24998
rect 106694 24954 112614 24955
rect 106694 24634 112838 24954
rect 113069 24871 113117 26373
rect 113197 26383 113231 26435
rect 113855 26414 113889 26435
rect 114513 26414 114547 26435
rect 115171 26414 115205 26435
rect 115829 26414 115863 26435
rect 113813 26383 113889 26414
rect 114471 26383 114547 26414
rect 115129 26383 115205 26414
rect 115787 26383 115863 26414
rect 113197 26286 113243 26383
rect 113813 26367 113901 26383
rect 114471 26367 114559 26383
rect 115129 26367 115217 26383
rect 115787 26367 115875 26383
rect 115886 26373 115900 26435
rect 115969 26414 116003 26435
rect 116083 26432 116128 26435
rect 116487 26432 116532 26435
rect 116083 26414 116117 26432
rect 116487 26414 116521 26432
rect 115969 26367 116016 26414
rect 116083 26383 116130 26414
rect 116071 26367 116130 26383
rect 116445 26367 116521 26414
rect 113245 26333 113901 26367
rect 113903 26333 114559 26367
rect 114561 26333 115217 26367
rect 115219 26333 115875 26367
rect 115877 26333 116521 26367
rect 113821 26327 113825 26333
rect 113849 26299 113853 26333
rect 113855 26286 113901 26333
rect 114513 26286 114559 26333
rect 115137 26327 115141 26333
rect 115165 26299 115169 26333
rect 115171 26286 115217 26333
rect 115829 26286 115875 26333
rect 113197 26274 113231 26286
rect 113830 26274 113843 26285
rect 113855 26274 113889 26286
rect 114488 26274 114501 26285
rect 114513 26274 114547 26286
rect 115146 26274 115159 26285
rect 115171 26274 115205 26286
rect 115804 26274 115817 26285
rect 115829 26274 115863 26286
rect 113183 24970 113231 26274
rect 113841 24970 113889 26274
rect 114499 24970 114547 26274
rect 113183 24898 113217 24970
rect 113841 24958 113875 24970
rect 114499 24958 114533 24970
rect 113219 24898 113223 24945
rect 113247 24911 113251 24917
rect 113827 24911 113875 24958
rect 114485 24911 114533 24958
rect 106694 24633 112614 24634
rect 106694 24526 112615 24633
rect 112654 24594 112655 24595
rect 112653 24593 112654 24594
rect 112668 24586 112695 24633
rect 106694 23322 112614 24526
rect 95270 22898 100800 22932
rect 95390 22786 95402 22898
rect 95390 21948 95402 22648
rect 96722 22516 96814 22664
rect 96860 22516 96894 22898
rect 96326 21982 96538 22430
rect 96722 22304 96894 22516
rect 96722 22206 96814 22304
rect 96860 21415 96894 22304
rect 93456 18262 94148 18300
rect 94744 18262 94806 18300
rect 95211 21379 96930 21415
rect 100453 21379 100487 21877
rect 95211 21345 103613 21379
rect 95211 18262 96930 21345
rect 100453 21265 100487 21345
rect 100542 21294 100549 21299
rect 100595 21294 101748 21299
rect 103100 21294 103458 21299
rect 100419 21231 100487 21265
rect 100508 21271 100636 21277
rect 103418 21271 103429 21276
rect 100508 21266 101748 21271
rect 103100 21266 103430 21271
rect 100508 21265 100636 21266
rect 103418 21265 103429 21266
rect 100508 21235 103429 21265
rect 103430 21235 103511 21250
rect 100508 21231 103511 21235
rect 100453 20607 100487 21231
rect 100539 21225 101748 21231
rect 103100 21225 103511 21231
rect 100539 21219 100636 21225
rect 103430 21213 103511 21225
rect 103430 21207 103527 21213
rect 100636 21201 101748 21207
rect 103100 21201 103527 21207
rect 100632 21197 103527 21201
rect 100508 21139 100589 21186
rect 100648 21176 103527 21197
rect 100636 21161 103558 21176
rect 103430 21155 103527 21161
rect 100526 20636 100549 20641
rect 100555 20620 100589 21139
rect 100608 21133 103471 21148
rect 100904 20641 102418 20669
rect 100595 20636 103458 20641
rect 103477 20635 103511 21155
rect 103517 21133 103530 21148
rect 100508 20619 100589 20620
rect 100508 20613 100636 20619
rect 103418 20613 103429 20618
rect 100498 20608 103430 20613
rect 100419 20573 100487 20607
rect 100508 20607 100636 20608
rect 103418 20607 103429 20608
rect 100508 20577 103429 20607
rect 103430 20577 103511 20592
rect 100508 20573 103511 20577
rect 100453 19949 100487 20573
rect 100539 20567 100960 20573
rect 102362 20567 103511 20573
rect 100539 20561 100636 20567
rect 103430 20555 103511 20567
rect 103430 20549 103527 20555
rect 100636 20543 100960 20549
rect 102362 20543 103527 20549
rect 103579 20543 103613 21345
rect 100632 20539 108624 20543
rect 100508 20481 100589 20528
rect 100648 20524 108624 20539
rect 100636 20509 108624 20524
rect 100636 20503 100960 20509
rect 102362 20503 103558 20509
rect 103430 20497 103527 20503
rect 100542 19974 100549 19983
rect 100555 19962 100589 20481
rect 100608 20475 100960 20496
rect 102362 20475 103471 20496
rect 100595 19974 101778 19983
rect 103130 19974 103458 19983
rect 103477 19977 103511 20497
rect 103517 20475 103530 20496
rect 100419 19915 100487 19949
rect 100508 19961 100589 19962
rect 100508 19955 100636 19961
rect 103418 19955 103429 19960
rect 100508 19949 101778 19955
rect 103130 19949 103430 19955
rect 100508 19946 103430 19949
rect 100508 19919 103429 19946
rect 103430 19919 103511 19934
rect 100508 19915 103511 19919
rect 97314 19434 97704 19468
rect 97314 19291 97348 19434
rect 97528 19366 97575 19413
rect 97490 19332 97575 19366
rect 97474 19291 97544 19303
rect 97670 19291 97704 19434
rect 97790 19434 98180 19468
rect 97790 19291 97824 19434
rect 98004 19404 98051 19413
rect 97912 19378 98051 19404
rect 98004 19376 98051 19378
rect 97940 19350 98051 19376
rect 97966 19332 98051 19350
rect 97940 19324 98012 19325
rect 97950 19297 98020 19303
rect 97912 19296 98040 19297
rect 97950 19291 98020 19296
rect 98146 19291 98180 19434
rect 100453 19291 100487 19915
rect 100539 19909 101778 19915
rect 103130 19909 103511 19915
rect 100539 19903 100636 19909
rect 103430 19897 103511 19909
rect 103430 19891 103527 19897
rect 100636 19885 101778 19891
rect 103130 19885 103527 19891
rect 100632 19881 103527 19885
rect 100508 19823 100589 19870
rect 100648 19854 103527 19881
rect 100636 19845 103558 19854
rect 103430 19839 103527 19845
rect 100542 19304 100549 19325
rect 100555 19304 100589 19823
rect 100608 19817 103471 19826
rect 101722 19789 103186 19817
rect 100882 19325 102396 19353
rect 100595 19304 103458 19325
rect 103477 19319 103511 19839
rect 103517 19817 103530 19826
rect 97280 19257 97704 19291
rect 97756 19257 98180 19291
rect 100419 19257 100487 19291
rect 100508 19303 100589 19304
rect 100508 19297 100636 19303
rect 103418 19297 103429 19302
rect 100508 19276 103430 19297
rect 100508 19261 103429 19276
rect 103430 19261 103511 19276
rect 100508 19257 103511 19261
rect 97314 18936 97348 19257
rect 97428 19097 97462 19257
rect 97474 19245 97475 19246
rect 97543 19245 97544 19246
rect 97473 19244 97474 19245
rect 97544 19244 97545 19245
rect 97556 19097 97590 19257
rect 97410 18936 97420 19076
rect 97438 18946 97476 19048
rect 97528 19038 97575 19085
rect 97490 19004 97575 19038
rect 97670 18936 97704 19257
rect 97314 18902 97704 18936
rect 97790 18936 97824 19257
rect 97904 19097 97938 19257
rect 97950 19245 97951 19246
rect 98019 19245 98020 19246
rect 97949 19244 97950 19245
rect 98020 19244 98021 19245
rect 98032 19097 98066 19257
rect 98004 19038 98051 19085
rect 97966 19004 98051 19038
rect 98146 18936 98180 19257
rect 97790 18902 98180 18936
rect 93246 18228 94148 18262
rect 94160 18228 94806 18262
rect 94818 18228 96930 18262
rect 97296 18232 97718 18852
rect 97772 18232 98194 18852
rect 100453 18633 100487 19257
rect 100539 19251 100938 19257
rect 102340 19251 103511 19257
rect 100539 19245 100636 19251
rect 103430 19239 103511 19251
rect 103430 19233 103527 19239
rect 100636 19227 100938 19233
rect 102340 19227 103527 19233
rect 100632 19223 103527 19227
rect 100508 19165 100589 19212
rect 100648 19193 103527 19223
rect 102340 19192 103180 19193
rect 103430 19192 103527 19193
rect 100636 19187 100938 19192
rect 102340 19187 103527 19192
rect 103430 19181 103527 19187
rect 100542 18652 100549 18667
rect 100555 18646 100589 19165
rect 100608 19159 100938 19164
rect 102340 19159 103471 19164
rect 100595 18652 101772 18667
rect 103124 18652 103458 18667
rect 103477 18661 103511 19181
rect 100419 18599 100487 18633
rect 100508 18645 100589 18646
rect 100508 18639 100636 18645
rect 103418 18639 103429 18644
rect 100508 18633 101772 18639
rect 103124 18633 103430 18639
rect 100508 18624 103430 18633
rect 100508 18603 103429 18624
rect 103430 18603 103511 18618
rect 100508 18599 103511 18603
rect 100453 18455 100487 18599
rect 100539 18593 101772 18599
rect 103124 18593 103511 18599
rect 100539 18587 100636 18593
rect 103430 18581 103511 18593
rect 103430 18575 103527 18581
rect 100636 18569 101772 18575
rect 103124 18569 103527 18575
rect 100632 18565 103527 18569
rect 100648 18538 103527 18565
rect 100648 18535 103542 18538
rect 103430 18534 103542 18535
rect 100636 18529 103558 18534
rect 103430 18523 103542 18529
rect 100608 18501 103471 18506
rect 103517 18501 103530 18506
rect 101716 18473 103180 18501
rect 103579 18455 103613 20509
rect 113069 20160 113103 24871
rect 113183 24809 113223 24898
rect 113243 24898 113251 24911
rect 113259 24898 113875 24911
rect 113243 24877 113875 24898
rect 113901 24877 113909 24911
rect 113917 24877 114533 24911
rect 113247 24871 113300 24877
rect 113242 24843 113300 24870
rect 113829 24861 113875 24877
rect 114487 24861 114533 24877
rect 113242 24809 113251 24843
rect 113841 24809 113875 24861
rect 114499 24809 114533 24861
rect 114535 24843 114539 24945
rect 115080 24917 115082 26014
rect 115108 24917 115110 25986
rect 115157 24970 115205 26274
rect 115815 24970 115863 26274
rect 115886 25260 115900 26327
rect 115969 25105 116003 26333
rect 116071 26286 116129 26333
rect 116083 25266 116117 26286
rect 116487 26285 116521 26333
rect 116462 26274 116521 26285
rect 116473 25254 116521 26274
rect 116461 25207 116533 25254
rect 116145 25173 116533 25207
rect 116402 25105 116404 25160
rect 116430 25105 116432 25160
rect 116461 25157 116533 25173
rect 116473 25142 116533 25157
rect 116473 25105 116521 25142
rect 116587 25105 116635 26435
rect 117378 26010 117452 26636
rect 117364 25856 117518 26010
rect 118023 25226 118042 27750
rect 118051 25254 118070 27750
rect 118118 26510 119557 31162
rect 120900 30004 120934 31162
rect 120162 29310 120624 29948
rect 120834 29922 120934 30004
rect 120220 29226 120570 29260
rect 120220 29198 120254 29226
rect 120220 28808 120288 29198
rect 120412 29158 120450 29196
rect 120378 29124 120450 29158
rect 120323 29074 120368 29085
rect 120411 29074 120456 29085
rect 120334 28898 120368 29074
rect 120422 28898 120456 29074
rect 120412 28848 120450 28886
rect 120378 28814 120450 28848
rect 120220 28746 120254 28808
rect 120536 28746 120570 29226
rect 120220 28712 120570 28746
rect 120862 28594 120898 28680
rect 118104 26474 119557 26510
rect 119584 26474 119618 26508
rect 120242 26474 120276 26508
rect 120900 26474 120934 29922
rect 120970 29528 120972 29606
rect 120970 26474 120972 26640
rect 121040 26474 121074 31162
rect 121154 30288 121199 31162
rect 121154 26474 121188 30288
rect 121558 30262 121603 31162
rect 121558 26474 121592 30262
rect 121672 26474 121706 31162
rect 121812 26505 121846 32514
rect 122122 31902 122584 32540
rect 122598 31902 123060 32540
rect 122176 31818 122526 31852
rect 122176 31338 122210 31818
rect 122368 31750 122406 31788
rect 122334 31716 122406 31750
rect 122279 31666 122324 31677
rect 122367 31666 122412 31677
rect 122290 31490 122324 31666
rect 122378 31490 122412 31666
rect 122368 31440 122406 31478
rect 122334 31406 122406 31440
rect 122492 31338 122526 31818
rect 122176 31304 122526 31338
rect 122652 31818 123002 31852
rect 122652 31338 122686 31818
rect 122844 31750 122882 31788
rect 122810 31716 122882 31750
rect 122755 31666 122800 31677
rect 122843 31666 122888 31677
rect 122766 31490 122800 31666
rect 122854 31490 122888 31666
rect 122844 31440 122882 31478
rect 122810 31406 122882 31440
rect 122968 31338 123002 31818
rect 122652 31304 123002 31338
rect 121848 31186 121884 31272
rect 124444 26505 124478 33256
rect 118104 26440 121706 26474
rect 118104 26410 119557 26440
rect 118104 26338 119580 26410
rect 119584 26388 119618 26440
rect 120200 26406 120238 26410
rect 118104 25207 119557 26338
rect 119584 26300 119630 26388
rect 120200 26372 120240 26406
rect 119632 26338 120240 26372
rect 120196 26332 120212 26338
rect 120236 26332 120240 26338
rect 120224 26304 120240 26332
rect 120242 26388 120276 26440
rect 120242 26300 120288 26388
rect 120858 26372 120896 26410
rect 120290 26338 120896 26372
rect 120900 26388 120934 26440
rect 120900 26300 120946 26388
rect 120956 26378 120972 26440
rect 121026 26404 121028 26440
rect 121012 26378 121028 26404
rect 121040 26410 121074 26440
rect 121154 26410 121188 26440
rect 121040 26372 121078 26410
rect 121154 26388 121192 26410
rect 121142 26372 121200 26388
rect 121516 26372 121554 26410
rect 120948 26338 121554 26372
rect 119559 26288 119572 26299
rect 119584 26288 119618 26300
rect 120217 26288 120230 26299
rect 120242 26288 120276 26300
rect 120875 26288 120888 26299
rect 120900 26288 120934 26300
rect 118103 25173 119557 25207
rect 118104 25105 119557 25173
rect 115969 25071 119557 25105
rect 115157 24958 115191 24970
rect 115815 24958 115849 24970
rect 114563 24911 114567 24917
rect 115143 24911 115191 24958
rect 115801 24911 115849 24958
rect 114559 24877 114567 24911
rect 114575 24877 115191 24911
rect 115217 24877 115225 24911
rect 115233 24877 115849 24911
rect 114563 24871 114567 24877
rect 115080 24864 115082 24871
rect 115108 24836 115110 24871
rect 115145 24861 115191 24877
rect 115803 24861 115849 24877
rect 115157 24809 115191 24861
rect 115815 24809 115849 24861
rect 115851 24843 115855 24945
rect 116402 24917 116404 25071
rect 116430 24917 116432 25071
rect 116473 24970 116521 25071
rect 116473 24958 116507 24970
rect 115879 24911 115883 24917
rect 116459 24911 116507 24958
rect 115875 24877 115883 24911
rect 115891 24877 116507 24911
rect 115879 24871 115883 24877
rect 116402 24864 116404 24871
rect 116430 24836 116432 24871
rect 116461 24861 116507 24877
rect 116473 24809 116507 24861
rect 116587 24871 116635 25071
rect 118104 25035 119557 25071
rect 118140 24894 118188 25035
rect 118254 24984 118302 25035
rect 113171 24775 116519 24809
rect 113214 24642 113223 24775
rect 113242 24670 113251 24775
rect 115816 24430 115855 24775
rect 115872 24430 115883 24726
rect 116587 20160 116621 24871
rect 118140 20160 118174 24894
rect 118254 24832 118288 24984
rect 118290 24866 118294 24968
rect 118840 24940 118848 25035
rect 118868 24940 118876 25035
rect 118912 24984 118960 25035
rect 119570 24984 119618 26288
rect 120228 24984 120276 26288
rect 120304 25182 120324 25706
rect 120886 24984 120934 26288
rect 120956 25238 120972 26332
rect 121012 25196 121028 26332
rect 121040 25128 121074 26338
rect 121142 26300 121200 26338
rect 121154 25280 121188 26300
rect 121558 26299 121592 26440
rect 121533 26288 121592 26299
rect 121544 25268 121592 26288
rect 121532 25230 121604 25268
rect 121216 25196 121604 25230
rect 121468 25128 121474 25184
rect 121496 25128 121502 25184
rect 121532 25180 121604 25196
rect 121544 25165 121604 25180
rect 121544 25128 121592 25165
rect 121658 25128 121706 26440
rect 121789 26469 124628 26505
rect 124725 26469 124759 33341
rect 124839 26469 124873 33242
rect 121789 26436 125377 26469
rect 121789 26435 125402 26436
rect 121714 25728 121734 26358
rect 121789 26330 124628 26435
rect 124633 26333 124639 26367
rect 121742 26314 124628 26330
rect 121742 26052 124639 26314
rect 121742 25836 124628 26052
rect 121742 25756 124639 25836
rect 121789 25636 124639 25756
rect 121789 25614 124628 25636
rect 121714 25312 121734 25568
rect 121778 25540 124628 25614
rect 124644 25580 124698 25606
rect 121742 25436 124628 25540
rect 121742 25340 124639 25436
rect 121730 25236 121734 25312
rect 121789 25310 124639 25340
rect 121758 25236 124639 25310
rect 121789 25190 124628 25236
rect 121730 25184 121734 25190
rect 121758 25140 124628 25190
rect 121742 25128 124628 25140
rect 121040 25094 124628 25128
rect 118912 24972 118946 24984
rect 119570 24972 119604 24984
rect 120228 24972 120262 24984
rect 120886 24972 120920 24984
rect 121468 24972 121474 25094
rect 121496 24972 121502 25094
rect 121544 24984 121592 25094
rect 121544 24972 121578 24984
rect 118318 24934 118322 24940
rect 118898 24934 118946 24972
rect 119556 24934 119604 24972
rect 118314 24900 118322 24934
rect 118330 24900 118946 24934
rect 118972 24900 118980 24934
rect 118988 24900 119604 24934
rect 118318 24894 118322 24900
rect 118840 24888 118848 24894
rect 118868 24860 118876 24894
rect 118900 24884 118946 24900
rect 119558 24884 119604 24900
rect 118912 24832 118946 24884
rect 119570 24832 119604 24884
rect 119606 24866 119610 24968
rect 119634 24934 119638 24940
rect 120214 24934 120262 24972
rect 120872 24934 120920 24972
rect 119630 24900 119638 24934
rect 119646 24900 120262 24934
rect 120288 24900 120296 24934
rect 120304 24900 120920 24934
rect 119634 24894 119638 24900
rect 120216 24884 120262 24900
rect 120874 24884 120920 24900
rect 120228 24832 120262 24884
rect 120886 24832 120920 24884
rect 120922 24866 120928 24968
rect 120950 24934 120956 24940
rect 121038 24934 121578 24972
rect 120946 24900 120956 24934
rect 120962 24900 121578 24934
rect 120950 24894 120956 24900
rect 121468 24882 121474 24894
rect 121496 24860 121502 24894
rect 121532 24884 121578 24900
rect 121544 24832 121578 24884
rect 121658 24894 121706 25094
rect 121789 25058 124628 25094
rect 124725 25105 124759 26435
rect 124839 26398 124886 26414
rect 124827 26367 124886 26398
rect 125012 26402 125402 26435
rect 125012 26374 125046 26402
rect 125201 26381 125248 26402
rect 124978 26367 125080 26374
rect 125201 26367 125273 26381
rect 124827 26333 125273 26367
rect 124827 26286 124885 26333
rect 124839 25276 124873 26286
rect 125012 25904 125046 26333
rect 125188 26300 125273 26333
rect 125229 26285 125263 26290
rect 125218 26274 125263 26285
rect 125229 26257 125263 26274
rect 125229 26252 125274 26257
rect 125115 26241 125160 26252
rect 125126 26065 125160 26241
rect 125229 26065 125288 26252
rect 125229 26053 125274 26065
rect 125226 26049 125274 26053
rect 125226 26006 125273 26049
rect 125188 25972 125273 26006
rect 125229 25904 125263 25972
rect 125343 25904 125402 26402
rect 125012 25870 125402 25904
rect 125488 26402 125878 26436
rect 125488 26374 125522 26402
rect 125488 25966 125556 26374
rect 125702 26334 125749 26381
rect 125664 26300 125749 26334
rect 125591 26241 125636 26252
rect 125719 26241 125764 26252
rect 125602 26065 125636 26241
rect 125730 26065 125764 26241
rect 125702 26006 125749 26053
rect 125664 25972 125749 26006
rect 125488 25904 125522 25966
rect 125844 25904 125878 26402
rect 125488 25870 125878 25904
rect 125229 25820 125263 25870
rect 125343 25820 125377 25870
rect 124839 25266 124884 25276
rect 124994 25254 125416 25820
rect 124854 25207 125416 25254
rect 124901 25200 125416 25207
rect 125470 25200 125892 25820
rect 126779 25226 126782 27750
rect 126807 25254 126810 27750
rect 126860 26474 128313 26510
rect 129796 26474 129830 33346
rect 179458 29428 180810 29430
rect 173556 28926 173612 28942
rect 173122 28157 181098 28191
rect 126860 26440 130448 26474
rect 126860 25207 128313 26440
rect 128952 26332 128968 26360
rect 128980 26306 128996 26332
rect 129664 26304 129684 26406
rect 129692 26332 129712 26378
rect 124901 25173 125377 25200
rect 126859 25173 128313 25207
rect 125217 25157 125275 25173
rect 125229 25142 125275 25157
rect 125229 25105 125263 25142
rect 125343 25105 125377 25173
rect 126860 25105 128313 25173
rect 124725 25071 128313 25105
rect 129796 25128 129830 26440
rect 129910 26403 129948 26410
rect 129898 26388 129948 26403
rect 129898 26372 129956 26388
rect 130272 26372 130310 26410
rect 129898 26338 130310 26372
rect 129898 26300 129956 26338
rect 129910 25280 129944 26300
rect 130289 26288 130334 26299
rect 130300 25268 130334 26288
rect 130288 25230 130346 25268
rect 129972 25196 130346 25230
rect 130288 25180 130346 25196
rect 130331 25165 130346 25180
rect 130300 25128 130334 25162
rect 130414 25128 130448 26440
rect 133902 25918 134022 25938
rect 134208 25920 134448 26472
rect 134208 25918 134498 25920
rect 133896 25890 134050 25910
rect 134208 25892 134448 25918
rect 134208 25890 134526 25892
rect 134208 25834 134448 25890
rect 134837 25834 134924 26726
rect 173585 26490 177245 26523
rect 178656 26490 181264 26524
rect 144050 25918 144170 25938
rect 144356 25920 144596 26472
rect 173603 26444 177227 26490
rect 178710 26462 181264 26474
rect 178710 26456 181332 26462
rect 173603 26432 177394 26444
rect 178744 26440 181178 26456
rect 181230 26440 181332 26456
rect 173603 26410 177227 26432
rect 178710 26415 181124 26422
rect 178710 26412 178744 26415
rect 178676 26410 178778 26412
rect 169460 26378 169486 26410
rect 169890 26378 169908 26410
rect 173600 26398 177428 26410
rect 178676 26406 181128 26410
rect 144356 25918 144646 25920
rect 144044 25890 144198 25910
rect 144356 25892 144596 25918
rect 144356 25890 144674 25892
rect 144356 25834 144596 25890
rect 129796 25094 133252 25128
rect 118242 24798 121590 24832
rect 118912 20160 118946 24798
rect 121658 20160 121692 24894
rect 121901 24822 121902 24908
rect 121758 24762 121933 24782
rect 121720 24032 121768 24040
rect 121720 23998 121734 24006
rect 121939 20160 121973 25058
rect 122108 24904 122530 25058
rect 122584 24904 123006 25058
rect 124588 25002 124611 25058
rect 125229 24964 125263 25071
rect 124572 24554 124611 24782
rect 124565 24498 124611 24554
rect 124572 24236 124611 24498
rect 124565 23482 124611 24236
rect 124628 23538 124639 24726
rect 125343 20160 125377 25071
rect 126860 25035 128313 25071
rect 130414 20160 130448 25094
rect 133350 24850 133362 25132
rect 133384 24884 133396 25106
rect 142468 23482 142668 23504
rect 168714 22344 168716 22400
rect 168714 22088 168716 22144
rect 168714 21944 168716 22000
rect 168714 21688 168716 21744
rect 131058 19468 131092 20160
rect 131138 19468 131146 19658
rect 131166 19502 131174 19686
rect 131166 19468 131196 19502
rect 122112 19434 122502 19468
rect 122112 18936 122146 19434
rect 122326 19366 122373 19413
rect 122288 19332 122373 19366
rect 122215 19273 122260 19284
rect 122343 19273 122388 19284
rect 122226 19097 122260 19273
rect 122354 19097 122388 19273
rect 122326 19038 122373 19085
rect 122288 19004 122373 19038
rect 122468 18936 122502 19434
rect 122112 18902 122502 18936
rect 122588 19434 122978 19468
rect 130964 19434 131258 19468
rect 122588 19406 122622 19434
rect 122588 18998 122656 19406
rect 122802 19366 122849 19413
rect 122764 19332 122849 19366
rect 122691 19273 122736 19284
rect 122819 19273 122864 19284
rect 122702 19097 122736 19273
rect 122830 19097 122864 19273
rect 122802 19038 122849 19085
rect 122764 19004 122849 19038
rect 122588 18936 122622 18998
rect 122944 18936 122978 19434
rect 131058 19400 131092 19434
rect 131058 19332 131116 19400
rect 131058 19072 131092 19332
rect 131110 19081 131126 19289
rect 131138 19285 131146 19434
rect 131166 19339 131174 19434
rect 131190 19339 131206 19434
rect 131138 19280 131150 19285
rect 131138 19273 131144 19280
rect 131134 19097 131144 19273
rect 131138 19081 131144 19097
rect 131160 19110 131210 19339
rect 131160 19085 131218 19110
rect 131058 19004 131116 19072
rect 131058 18970 131092 19004
rect 131118 18970 131122 19046
rect 131002 18950 131122 18970
rect 131058 18942 131092 18950
rect 131146 18942 131150 19074
rect 130996 18936 131150 18942
rect 131162 18936 131218 19085
rect 131224 18936 131258 19434
rect 122588 18902 122978 18936
rect 130964 18902 131258 18936
rect 131344 19434 131734 19468
rect 131344 18936 131378 19434
rect 131558 19366 131605 19413
rect 131520 19332 131605 19366
rect 131447 19273 131492 19284
rect 131575 19273 131620 19284
rect 131458 19097 131492 19273
rect 131586 19097 131620 19273
rect 131396 18936 131416 19084
rect 131558 19038 131605 19085
rect 131520 19004 131605 19038
rect 131700 18936 131734 19434
rect 131344 18902 131734 18936
rect 163778 19434 164168 19468
rect 163778 18936 163812 19434
rect 163992 19366 164039 19413
rect 163954 19332 164039 19366
rect 163881 19273 163926 19284
rect 164009 19273 164054 19284
rect 163892 19097 163926 19273
rect 164020 19097 164054 19273
rect 163992 19038 164039 19085
rect 163954 19004 164039 19038
rect 164134 18936 164168 19434
rect 163778 18902 164168 18936
rect 164254 19434 164644 19468
rect 164254 19406 164288 19434
rect 164254 18998 164322 19406
rect 164468 19366 164515 19413
rect 164430 19332 164515 19366
rect 164357 19273 164402 19284
rect 164485 19273 164530 19284
rect 164368 19097 164402 19273
rect 164496 19097 164530 19273
rect 164468 19038 164515 19085
rect 164430 19004 164515 19038
rect 164254 18936 164288 18998
rect 164610 18936 164644 19434
rect 164254 18902 164644 18936
rect 131058 18852 131092 18902
rect 131162 18900 131218 18902
rect 131098 18852 131218 18900
rect 100453 18421 108723 18455
rect 93342 15568 93376 18228
rect 93456 18160 93490 18228
rect 94080 18164 94092 18228
rect 94114 18160 94148 18228
rect 94772 18160 94806 18228
rect 95211 18160 96930 18228
rect 93438 18126 96930 18160
rect 93456 15658 93490 18126
rect 94114 15658 94148 18126
rect 95211 17975 96930 18126
rect 95211 17941 100800 17975
rect 95211 17791 96930 17941
rect 103579 17923 103613 18421
rect 122094 18239 122516 18852
rect 122001 18205 122569 18239
rect 122570 18232 122992 18852
rect 131022 18488 131272 18852
rect 131326 18488 131748 18852
rect 131088 18438 131122 18448
rect 131476 18438 131510 18448
rect 131564 18438 131598 18448
rect 131104 18404 131156 18414
rect 131442 18404 131632 18414
rect 131070 18370 131094 18404
rect 131104 18336 131128 18404
rect 131202 18302 131236 18314
rect 130980 18268 131236 18302
rect 131362 18302 131396 18314
rect 131678 18302 131712 18314
rect 131362 18268 131712 18302
rect 163760 18239 164182 18852
rect 163667 18205 164235 18239
rect 164236 18232 164658 18852
rect 169460 18328 169486 26332
rect 169890 18328 169908 26332
rect 171302 26288 171348 26300
rect 171308 26276 171348 26288
rect 170610 24602 170622 25706
rect 171338 22992 171348 26276
rect 173603 25500 177227 26398
rect 178676 26376 178744 26406
rect 178836 26376 181128 26406
rect 181264 26388 181275 26399
rect 181287 26388 181298 26399
rect 178710 25752 178744 26376
rect 178870 26342 179492 26376
rect 179528 26342 180150 26376
rect 180186 26342 180808 26376
rect 180844 26372 181124 26376
rect 181264 26372 181298 26388
rect 180844 26342 181298 26372
rect 178886 26338 179492 26342
rect 179544 26338 180150 26342
rect 180202 26338 180808 26342
rect 180860 26338 181298 26342
rect 181123 26300 181124 26301
rect 181124 26299 181125 26300
rect 178813 26288 178858 26299
rect 179471 26288 179516 26299
rect 180129 26288 180174 26299
rect 180787 26288 180832 26299
rect 178824 25752 178858 26288
rect 178869 25764 178870 25765
rect 179470 25764 179471 25765
rect 178870 25763 178871 25764
rect 179469 25763 179470 25764
rect 179482 25752 179516 26288
rect 179527 25764 179528 25765
rect 180128 25764 180129 25765
rect 179528 25763 179529 25764
rect 180127 25763 180128 25764
rect 180140 25752 180174 26288
rect 180185 25764 180186 25765
rect 180786 25764 180787 25765
rect 180186 25763 180187 25764
rect 180785 25763 180786 25764
rect 180798 25752 180832 26288
rect 181162 25780 181196 26338
rect 180843 25764 180844 25765
rect 180844 25763 180845 25764
rect 181112 25752 181123 25763
rect 178676 25718 181123 25752
rect 173603 25288 177268 25500
rect 173603 23006 177227 25288
rect 178710 25094 178744 25718
rect 178824 25094 178858 25718
rect 178870 25706 178871 25707
rect 179469 25706 179470 25707
rect 178869 25705 178870 25706
rect 179470 25705 179471 25706
rect 178869 25106 178870 25107
rect 179470 25106 179471 25107
rect 178870 25105 178871 25106
rect 179469 25105 179470 25106
rect 179482 25094 179516 25718
rect 179528 25706 179529 25707
rect 180127 25706 180128 25707
rect 179527 25705 179528 25706
rect 180128 25705 180129 25706
rect 179527 25106 179528 25107
rect 180128 25106 180129 25107
rect 179528 25105 179529 25106
rect 180127 25105 180128 25106
rect 180140 25094 180174 25718
rect 180730 25712 180792 25718
rect 180186 25706 180187 25707
rect 180785 25706 180786 25707
rect 180185 25705 180186 25706
rect 180758 25684 180792 25706
rect 180185 25106 180186 25107
rect 180786 25106 180787 25107
rect 180186 25105 180187 25106
rect 180785 25105 180786 25106
rect 180798 25094 180832 25718
rect 180838 25712 180922 25718
rect 180844 25706 180845 25707
rect 180838 25684 180894 25706
rect 181124 25690 181196 25728
rect 181162 25122 181196 25690
rect 180843 25106 180844 25107
rect 180844 25105 180845 25106
rect 181112 25094 181123 25105
rect 178676 25060 181123 25094
rect 178710 24436 178744 25060
rect 178824 24436 178858 25060
rect 178870 25048 178871 25049
rect 179469 25048 179470 25049
rect 178869 25047 178870 25048
rect 179470 25047 179471 25048
rect 178869 24448 178870 24449
rect 178870 24447 178871 24448
rect 179398 24442 179404 24504
rect 179426 24442 179432 24476
rect 179470 24448 179471 24449
rect 179469 24447 179470 24448
rect 179482 24436 179516 25060
rect 179528 25048 179529 25049
rect 180127 25048 180128 25049
rect 179527 25047 179528 25048
rect 180128 25047 180129 25048
rect 179527 24448 179528 24449
rect 180128 24448 180129 24449
rect 179528 24447 179529 24448
rect 180127 24447 180128 24448
rect 180140 24436 180174 25060
rect 180186 25048 180187 25049
rect 180785 25048 180786 25049
rect 180185 25047 180186 25048
rect 180786 25047 180787 25048
rect 180185 24448 180186 24449
rect 180786 24448 180787 24449
rect 180186 24447 180187 24448
rect 180785 24447 180786 24448
rect 180798 24436 180832 25060
rect 180844 25048 180845 25049
rect 180843 25047 180844 25048
rect 181124 25032 181196 25070
rect 181162 24464 181196 25032
rect 180843 24448 180844 24449
rect 180844 24447 180845 24448
rect 181112 24436 181123 24447
rect 178676 24402 181123 24436
rect 178710 23778 178744 24402
rect 178824 23778 178858 24402
rect 178870 24390 178871 24391
rect 178869 24389 178870 24390
rect 179398 24312 179404 24396
rect 179426 24340 179432 24396
rect 179469 24390 179470 24391
rect 179470 24389 179471 24390
rect 178869 23790 178870 23791
rect 179470 23790 179471 23791
rect 178870 23789 178871 23790
rect 179469 23789 179470 23790
rect 179482 23778 179516 24402
rect 179528 24390 179529 24391
rect 180127 24390 180128 24391
rect 179527 24389 179528 24390
rect 180128 24389 180129 24390
rect 179527 23790 179528 23791
rect 180128 23790 180129 23791
rect 179528 23789 179529 23790
rect 180127 23789 180128 23790
rect 180140 23778 180174 24402
rect 180186 24390 180187 24391
rect 180785 24390 180786 24391
rect 180185 24389 180186 24390
rect 180786 24389 180787 24390
rect 180185 23790 180186 23791
rect 180786 23790 180787 23791
rect 180186 23789 180187 23790
rect 180785 23789 180786 23790
rect 180798 23778 180832 24402
rect 180844 24390 180845 24391
rect 180843 24389 180844 24390
rect 181124 24374 181196 24412
rect 181162 23806 181196 24374
rect 180843 23790 180844 23791
rect 180844 23789 180845 23790
rect 181112 23778 181123 23789
rect 178676 23744 181123 23778
rect 178710 23120 178744 23744
rect 178824 23120 178858 23744
rect 178870 23732 178871 23733
rect 179469 23732 179470 23733
rect 178869 23731 178870 23732
rect 179470 23731 179471 23732
rect 178869 23132 178870 23133
rect 178870 23131 178871 23132
rect 179400 23126 179404 23196
rect 179428 23126 179432 23168
rect 179470 23132 179471 23133
rect 179469 23131 179470 23132
rect 179482 23120 179516 23744
rect 179528 23732 179529 23733
rect 180127 23732 180128 23733
rect 179527 23731 179528 23732
rect 180128 23731 180129 23732
rect 179527 23132 179528 23133
rect 180128 23132 180129 23133
rect 179528 23131 179529 23132
rect 180127 23131 180128 23132
rect 180140 23120 180174 23744
rect 180186 23732 180187 23733
rect 180785 23732 180786 23733
rect 180185 23731 180186 23732
rect 180786 23731 180787 23732
rect 180185 23132 180186 23133
rect 180786 23132 180787 23133
rect 180186 23131 180187 23132
rect 180785 23131 180786 23132
rect 180798 23120 180832 23744
rect 180844 23732 180845 23733
rect 180843 23731 180844 23732
rect 181124 23716 181196 23754
rect 181162 23148 181196 23716
rect 180843 23132 180844 23133
rect 180844 23131 180845 23132
rect 181112 23120 181123 23131
rect 178676 23086 181123 23120
rect 178710 23006 178744 23086
rect 178824 23006 178858 23086
rect 179400 23006 179404 23080
rect 179428 23032 179432 23080
rect 179482 23006 179516 23086
rect 180140 23006 180174 23086
rect 180798 23006 180832 23086
rect 181264 23006 181298 26338
rect 173603 22972 181298 23006
rect 173603 22936 177227 22972
rect 177832 22936 178294 22972
rect 173639 22601 173673 22936
rect 174373 22798 174384 22884
rect 174411 22760 174422 22922
rect 177157 22601 177191 22936
rect 177868 22601 177902 22848
rect 178224 22601 178258 22848
rect 178710 22637 178744 22972
rect 178674 22601 181347 22637
rect 173041 22567 181347 22601
rect 173056 22487 173676 22567
rect 173753 22552 173787 22567
rect 173726 22518 174292 22552
rect 173726 22487 173787 22518
rect 174258 22506 174292 22518
rect 174411 22506 174445 22567
rect 173856 22487 174510 22506
rect 175069 22487 175103 22567
rect 175727 22487 175761 22567
rect 176385 22487 176419 22567
rect 177043 22487 177077 22567
rect 177157 22487 177191 22567
rect 173056 22456 177191 22487
rect 173056 22425 173676 22456
rect 173047 22386 173676 22425
rect 172974 22300 173676 22386
rect 173047 22148 173676 22300
rect 173726 22453 177191 22456
rect 173726 22423 173787 22453
rect 173799 22441 173800 22442
rect 173798 22440 173799 22441
rect 173856 22432 174510 22453
rect 175056 22441 175057 22442
rect 175057 22440 175058 22441
rect 173905 22423 174184 22432
rect 173726 22376 173862 22423
rect 173905 22419 174190 22423
rect 173921 22404 174190 22419
rect 173726 22196 173787 22376
rect 173828 22338 173862 22376
rect 173972 22338 174190 22404
rect 173972 22310 174184 22338
rect 173921 22276 174184 22310
rect 173972 22196 174184 22276
rect 174258 22196 174292 22432
rect 174373 22322 174384 22408
rect 173726 22162 174292 22196
rect 173047 22094 173081 22148
rect 173639 22094 173673 22148
rect 173047 21857 173676 22094
rect 173753 22076 173787 22162
rect 173972 22076 174184 22162
rect 173056 21672 173676 21857
rect 173726 22042 174292 22076
rect 173726 21947 173787 22042
rect 173972 22028 174184 22042
rect 174097 21962 174108 21973
rect 173726 21900 173862 21947
rect 173921 21928 174108 21962
rect 174109 21900 174190 21947
rect 173726 21829 173787 21900
rect 173828 21846 173862 21900
rect 174156 21846 174190 21900
rect 173798 21841 173799 21842
rect 173799 21840 173800 21841
rect 174097 21840 174108 21845
rect 174258 21840 174292 22042
rect 174411 21842 174456 22432
rect 174399 21841 174400 21842
rect 174411 21841 174457 21842
rect 175057 21841 175058 21842
rect 174398 21840 174399 21841
rect 173905 21834 173921 21840
rect 174097 21834 174113 21840
rect 173905 21829 174113 21834
rect 174258 21829 174399 21840
rect 174411 21829 174445 21841
rect 174457 21840 174458 21841
rect 175056 21840 175057 21841
rect 174457 21829 174482 21840
rect 175069 21829 175103 22453
rect 175115 22441 175116 22442
rect 175714 22441 175715 22442
rect 175114 22440 175115 22441
rect 175715 22440 175716 22441
rect 175114 21841 175115 21842
rect 175715 21841 175716 21842
rect 175115 21840 175116 21841
rect 175714 21840 175715 21841
rect 175727 21829 175761 22453
rect 175773 22441 175774 22442
rect 176372 22441 176373 22442
rect 175772 22440 175773 22441
rect 176373 22440 176374 22441
rect 175772 21841 175773 21842
rect 176373 21841 176374 21842
rect 175773 21840 175774 21841
rect 176372 21840 176373 21841
rect 176385 21829 176419 22453
rect 176431 22441 176432 22442
rect 177030 22441 177031 22442
rect 176430 22440 176431 22441
rect 177031 22440 177032 22441
rect 177043 22268 177077 22453
rect 177157 22268 177191 22453
rect 177868 22412 177902 22567
rect 178044 22514 178082 22521
rect 178013 22487 178129 22499
rect 178013 22484 178113 22487
rect 178028 22464 178098 22484
rect 178224 22412 178258 22567
rect 177868 22378 178258 22412
rect 177292 22296 177410 22376
rect 177266 22268 177410 22296
rect 176870 22244 177410 22268
rect 176870 22056 177318 22244
rect 176430 21841 176431 21842
rect 177031 21841 177032 21842
rect 176431 21840 176432 21841
rect 177030 21840 177031 21841
rect 177043 21829 177077 22056
rect 177157 21829 177191 22056
rect 173726 21795 177191 21829
rect 177854 21818 178276 22328
rect 177852 21795 178658 21818
rect 173726 21720 173787 21795
rect 173799 21783 173800 21784
rect 173798 21782 173799 21783
rect 174258 21720 174292 21795
rect 174398 21783 174399 21784
rect 174411 21783 174445 21795
rect 174457 21783 174458 21784
rect 175056 21783 175057 21784
rect 174399 21782 174400 21783
rect 174411 21782 174457 21783
rect 175057 21782 175058 21783
rect 173726 21686 174292 21720
rect 174411 21688 174456 21782
rect 173639 21171 173673 21672
rect 173753 21171 173787 21686
rect 173798 21183 173799 21184
rect 174399 21183 174400 21184
rect 173799 21182 173800 21183
rect 174398 21182 174399 21183
rect 174411 21171 174445 21688
rect 174456 21183 174457 21184
rect 175057 21183 175058 21184
rect 174457 21182 174458 21183
rect 175056 21182 175057 21183
rect 175069 21171 175103 21795
rect 175115 21783 175116 21784
rect 175714 21783 175715 21784
rect 175114 21782 175115 21783
rect 175715 21782 175716 21783
rect 175114 21183 175115 21184
rect 175715 21183 175716 21184
rect 175115 21182 175116 21183
rect 175714 21182 175715 21183
rect 175727 21171 175761 21795
rect 175773 21783 175774 21784
rect 176372 21783 176373 21784
rect 175772 21782 175773 21783
rect 176373 21782 176374 21783
rect 175772 21183 175773 21184
rect 176373 21183 176374 21184
rect 175773 21182 175774 21183
rect 176372 21182 176373 21183
rect 176385 21171 176419 21795
rect 176431 21783 176432 21784
rect 177030 21783 177031 21784
rect 176430 21782 176431 21783
rect 177031 21782 177032 21783
rect 176430 21183 176431 21184
rect 177031 21183 177032 21184
rect 176431 21182 176432 21183
rect 177030 21182 177031 21183
rect 177043 21171 177077 21795
rect 177157 21171 177191 21795
rect 177854 21784 178276 21795
rect 177854 21761 178624 21784
rect 177854 21708 178276 21761
rect 173605 21137 177191 21171
rect 173639 21078 173673 21137
rect 173554 21068 173747 21078
rect 173639 21050 173673 21068
rect 173526 21040 173747 21050
rect 173639 20513 173673 21040
rect 173753 20513 173787 21137
rect 173799 21125 173800 21126
rect 174398 21125 174399 21126
rect 173798 21124 173799 21125
rect 174399 21124 174400 21125
rect 173798 20525 173799 20526
rect 174399 20525 174400 20526
rect 173799 20524 173800 20525
rect 174398 20524 174399 20525
rect 174411 20513 174445 21137
rect 174457 21125 174458 21126
rect 175056 21125 175057 21126
rect 174456 21124 174457 21125
rect 175057 21124 175058 21125
rect 174456 20525 174457 20526
rect 175057 20525 175058 20526
rect 174457 20524 174458 20525
rect 175056 20524 175057 20525
rect 175069 20513 175103 21137
rect 175115 21125 175116 21126
rect 175714 21125 175715 21126
rect 175114 21124 175115 21125
rect 175715 21124 175716 21125
rect 175114 20525 175115 20526
rect 175715 20525 175716 20526
rect 175115 20524 175116 20525
rect 175714 20524 175715 20525
rect 175727 20513 175761 21137
rect 175773 21125 175774 21126
rect 176372 21125 176373 21126
rect 175772 21124 175773 21125
rect 176373 21124 176374 21125
rect 175772 20525 175773 20526
rect 176373 20525 176374 20526
rect 175773 20524 175774 20525
rect 176372 20524 176373 20525
rect 176385 20513 176419 21137
rect 176431 21125 176432 21126
rect 177030 21125 177031 21126
rect 176430 21124 176431 21125
rect 177031 21124 177032 21125
rect 176430 20525 176431 20526
rect 177031 20525 177032 20526
rect 176431 20524 176432 20525
rect 177030 20524 177031 20525
rect 177043 20513 177077 21137
rect 177157 20513 177191 21137
rect 173605 20479 177191 20513
rect 171356 18566 171380 19968
rect 173639 19855 173673 20479
rect 173753 19855 173787 20479
rect 173799 20467 173800 20468
rect 174398 20467 174399 20468
rect 173798 20466 173799 20467
rect 174399 20466 174400 20467
rect 173798 19867 173799 19868
rect 174399 19867 174400 19868
rect 173799 19866 173800 19867
rect 174398 19866 174399 19867
rect 174411 19855 174445 20479
rect 174457 20467 174458 20468
rect 175056 20467 175057 20468
rect 174456 20466 174457 20467
rect 175057 20466 175058 20467
rect 174456 19867 174457 19868
rect 175057 19867 175058 19868
rect 174457 19866 174458 19867
rect 175056 19866 175057 19867
rect 175069 19855 175103 20479
rect 175115 20467 175116 20468
rect 175714 20467 175715 20468
rect 175114 20466 175115 20467
rect 175715 20466 175716 20467
rect 175114 19867 175115 19868
rect 175715 19867 175716 19868
rect 175115 19866 175116 19867
rect 175714 19866 175715 19867
rect 175727 19855 175761 20479
rect 175773 20467 175774 20468
rect 176372 20467 176373 20468
rect 175772 20466 175773 20467
rect 176373 20466 176374 20467
rect 175772 19867 175773 19868
rect 176373 19867 176374 19868
rect 175773 19866 175774 19867
rect 176372 19866 176373 19867
rect 176385 19855 176419 20479
rect 176431 20467 176432 20468
rect 177030 20467 177031 20468
rect 176430 20466 176431 20467
rect 177031 20466 177032 20467
rect 176430 19867 176431 19868
rect 177031 19867 177032 19868
rect 176431 19866 176432 19867
rect 177030 19866 177031 19867
rect 177043 19855 177077 20479
rect 177157 19855 177191 20479
rect 173605 19821 177191 19855
rect 172598 19280 172600 19686
rect 172626 19280 172656 19658
rect 172945 19468 172979 19522
rect 172945 19436 172978 19468
rect 172911 19015 172924 19436
rect 172945 19083 172979 19436
rect 173010 19434 173400 19468
rect 173010 19083 173044 19434
rect 173047 19209 173078 19434
rect 173224 19366 173271 19413
rect 173186 19332 173271 19366
rect 173366 19302 173400 19434
rect 173112 19284 173128 19285
rect 173112 19197 173158 19284
rect 173241 19273 173286 19284
rect 173292 19280 173586 19302
rect 173366 19274 173400 19280
rect 173169 19209 173170 19210
rect 173240 19209 173241 19210
rect 173170 19208 173171 19209
rect 173239 19208 173240 19209
rect 173252 19197 173286 19273
rect 173292 19252 173558 19274
rect 173366 19197 173400 19252
rect 173639 19197 173673 19821
rect 173753 19197 173787 19821
rect 173799 19809 173800 19810
rect 174398 19809 174399 19810
rect 173798 19808 173799 19809
rect 174399 19808 174400 19809
rect 173798 19209 173799 19210
rect 174399 19209 174400 19210
rect 173799 19208 173800 19209
rect 174398 19208 174399 19209
rect 174411 19197 174445 19821
rect 174457 19809 174458 19810
rect 175056 19809 175057 19810
rect 174456 19808 174457 19809
rect 175057 19808 175058 19809
rect 174456 19209 174457 19210
rect 175057 19209 175058 19210
rect 174457 19208 174458 19209
rect 175056 19208 175057 19209
rect 175069 19197 175103 19821
rect 175115 19809 175116 19810
rect 175714 19809 175715 19810
rect 175114 19808 175115 19809
rect 175715 19808 175716 19809
rect 175114 19209 175115 19210
rect 175715 19209 175716 19210
rect 175115 19208 175116 19209
rect 175714 19208 175715 19209
rect 175727 19197 175761 19821
rect 175773 19809 175774 19810
rect 176372 19809 176373 19810
rect 175772 19808 175773 19809
rect 176373 19808 176374 19809
rect 175772 19209 175773 19210
rect 176373 19209 176374 19210
rect 175773 19208 175774 19209
rect 176372 19208 176373 19209
rect 176385 19197 176419 19821
rect 176431 19809 176432 19810
rect 177030 19809 177031 19810
rect 176430 19808 176431 19809
rect 177031 19808 177032 19809
rect 176430 19209 176431 19210
rect 177031 19209 177032 19210
rect 176431 19208 176432 19209
rect 177030 19208 177031 19209
rect 177043 19197 177077 19821
rect 177157 19197 177191 19821
rect 173112 19194 173400 19197
rect 173124 19163 173400 19194
rect 173605 19163 177191 19197
rect 173124 19137 173158 19163
rect 173252 19137 173286 19163
rect 173112 19085 173170 19137
rect 173240 19085 173298 19137
rect 173366 19083 173400 19163
rect 173639 19083 173673 19163
rect 173753 19083 173787 19163
rect 174411 19083 174445 19163
rect 175069 19083 175103 19163
rect 175727 19083 175761 19163
rect 176385 19083 176419 19163
rect 177043 19083 177077 19163
rect 177157 19083 177191 19163
rect 178674 19083 181347 22567
rect 182660 19422 183032 20126
rect 172945 19049 172978 19083
rect 173010 19049 181347 19083
rect 173010 19013 173044 19049
rect 173170 19015 173240 19038
rect 172668 18950 172788 18970
rect 172974 18952 173214 19013
rect 173366 18998 173400 19049
rect 173639 19013 173673 19049
rect 172974 18950 173264 18952
rect 172662 18922 172816 18942
rect 172974 18924 173214 18950
rect 172974 18922 173292 18924
rect 172974 18866 173214 18922
rect 173603 18866 173690 19013
rect 171308 18312 171348 18324
rect 171302 18300 171348 18312
rect 131180 18090 131184 18180
rect 131208 18106 131212 18152
rect 172116 17882 172128 18164
rect 172150 17916 172162 18138
rect 172642 18090 172656 18444
rect 173639 18199 173673 18866
rect 177157 18386 177191 19049
rect 178674 19013 181347 19049
rect 180122 19002 180196 19013
rect 183122 18866 183362 19504
rect 176550 18137 177191 18386
rect 176550 18067 177170 18137
rect 177186 18103 177191 18137
rect 177220 18103 177245 18372
rect 177220 18078 177225 18103
rect 172684 17806 172760 17808
rect 172684 17804 172756 17806
rect 95430 17352 95464 17791
rect 95522 17790 96070 17791
rect 96120 17736 96780 17791
rect 96088 17352 96122 17386
rect 96746 17352 96780 17736
rect 96860 17352 96894 17791
rect 172656 17778 172788 17780
rect 172656 17776 172784 17778
rect 104855 17534 104872 17590
rect 172648 17561 172682 17566
rect 172776 17561 172810 17566
rect 172614 17527 172716 17532
rect 172742 17527 172844 17532
rect 172914 17530 172924 17584
rect 95380 17318 100800 17352
rect 172932 17346 172960 17566
rect 172968 17382 172978 17530
rect 173154 17382 181130 17416
rect 95380 17252 95414 17318
rect 95380 15642 95418 17252
rect 95430 17214 95464 17318
rect 96088 17272 96122 17318
rect 95516 17252 96514 17272
rect 96088 17238 96122 17252
rect 96514 17238 96734 17249
rect 96746 17238 96780 17318
rect 96860 17238 96894 17318
rect 95550 17218 96894 17238
rect 95430 17176 95516 17214
rect 95566 17204 96894 17218
rect 96075 17192 96076 17193
rect 96076 17191 96077 17192
rect 95430 16558 95464 17176
rect 95466 16592 95476 17176
rect 95482 16608 95516 17176
rect 95482 16592 95498 16608
rect 96076 16592 96077 16593
rect 96075 16591 96076 16592
rect 96088 16580 96122 17204
rect 96134 17192 96135 17193
rect 96733 17192 96734 17193
rect 96133 17191 96134 17192
rect 96734 17191 96735 17192
rect 96133 16592 96134 16593
rect 96734 16592 96735 16593
rect 96134 16591 96135 16592
rect 96733 16591 96734 16592
rect 96746 16580 96780 17204
rect 96860 16580 96894 17204
rect 100108 17198 100164 17208
rect 101858 17156 102962 17180
rect 100108 17142 100164 17152
rect 101830 17128 102990 17152
rect 103694 16902 103728 17256
rect 100476 16868 108728 16902
rect 97278 16682 97740 16850
rect 97754 16682 98216 16850
rect 97116 16672 98216 16682
rect 95430 16556 95470 16558
rect 95430 16530 95516 16556
rect 95566 16546 96894 16580
rect 96075 16534 96076 16535
rect 96076 16533 96077 16534
rect 95430 16484 95522 16530
rect 95430 16468 95516 16484
rect 95430 16020 95464 16468
rect 95466 16020 95476 16468
rect 95482 16020 95516 16468
rect 96010 16454 96052 16468
rect 95430 15950 95516 16020
rect 95430 15938 95498 15950
rect 95430 15934 95476 15938
rect 95482 15934 95498 15938
rect 96076 15934 96077 15935
rect 95430 15910 95470 15934
rect 96075 15933 96076 15934
rect 96088 15922 96122 16546
rect 96134 16534 96135 16535
rect 96733 16534 96734 16535
rect 96133 16533 96134 16534
rect 96734 16533 96735 16534
rect 96160 16454 96214 16468
rect 96662 16454 96740 16468
rect 96133 15934 96134 15935
rect 96734 15934 96735 15935
rect 96134 15933 96135 15934
rect 96733 15933 96734 15934
rect 96746 15922 96780 16546
rect 96860 15922 96894 16546
rect 97278 16212 97740 16672
rect 97754 16212 98216 16672
rect 100476 16712 100510 16868
rect 103554 16788 103657 16800
rect 100662 16785 103657 16788
rect 100540 16726 100612 16764
rect 100662 16754 103642 16785
rect 103554 16742 103642 16754
rect 100476 16672 100572 16712
rect 100476 16580 100510 16672
rect 100566 16644 100572 16656
rect 100578 16592 100612 16726
rect 100618 16672 103586 16712
rect 100618 16644 103586 16656
rect 103592 16608 103626 16742
rect 103632 16672 103658 16712
rect 103632 16644 103686 16656
rect 100562 16584 100650 16592
rect 100540 16580 100650 16584
rect 103542 16580 103553 16591
rect 100442 16546 103553 16580
rect 97332 16128 97682 16162
rect 97332 16040 97366 16128
rect 97542 16100 97552 16102
rect 97524 16060 97562 16098
rect 96956 16020 97440 16040
rect 97490 16026 97562 16060
rect 96956 16014 97130 16020
rect 97332 15984 97366 16020
rect 97440 15987 97468 15988
rect 97435 15984 97480 15987
rect 97130 15964 97480 15984
rect 97523 15976 97568 15987
rect 97332 15922 97366 15964
rect 97446 15922 97480 15964
rect 97491 15934 97492 15935
rect 97522 15934 97523 15935
rect 97492 15933 97493 15934
rect 97521 15933 97522 15934
rect 97534 15922 97568 15976
rect 97648 15922 97682 16128
rect 97808 16128 98158 16162
rect 97690 16020 97764 16040
rect 97690 15964 97764 15984
rect 97808 15922 97842 16128
rect 98000 16060 98038 16098
rect 97862 16020 97916 16040
rect 97966 16026 98038 16060
rect 97916 15987 97944 15988
rect 97911 15984 97956 15987
rect 97862 15964 97956 15984
rect 97999 15976 98044 15987
rect 97922 15922 97956 15964
rect 97967 15934 97968 15935
rect 97998 15934 97999 15935
rect 97968 15933 97969 15934
rect 97997 15933 97998 15934
rect 98004 15928 98044 15976
rect 98010 15922 98044 15928
rect 98124 15922 98158 16128
rect 100476 15922 100510 16546
rect 100562 16534 100650 16546
rect 100578 16158 100612 16534
rect 103554 16518 103626 16556
rect 103592 16142 103626 16518
rect 103554 16130 103642 16142
rect 100540 16068 100612 16106
rect 100662 16096 103642 16130
rect 103554 16084 103642 16096
rect 100578 15934 100612 16068
rect 100622 16020 103586 16060
rect 100678 15964 103586 16004
rect 103592 15950 103626 16084
rect 103632 16020 103652 16060
rect 103694 16004 103728 16868
rect 172158 16384 172478 16826
rect 173486 16128 174846 16142
rect 103632 15964 103728 16004
rect 100562 15926 100650 15934
rect 100540 15922 100650 15926
rect 103542 15922 103553 15933
rect 95430 15900 95464 15910
rect 95430 15898 95470 15900
rect 95430 15804 95516 15898
rect 95566 15888 103553 15922
rect 96075 15876 96076 15877
rect 96076 15875 96077 15876
rect 95430 15661 95464 15804
rect 95466 15661 95476 15804
rect 95430 15646 95476 15661
rect 95430 15642 95464 15646
rect 95380 15574 95436 15642
rect 95482 15608 95516 15804
rect 96088 15658 96122 15888
rect 96134 15876 96135 15877
rect 96733 15876 96734 15877
rect 96133 15875 96134 15876
rect 96734 15875 96735 15876
rect 96746 15658 96780 15888
rect 95553 15646 95554 15647
rect 95554 15645 95555 15646
rect 96060 15608 96098 15646
rect 96718 15608 96756 15646
rect 95482 15574 96098 15608
rect 96150 15574 96756 15608
rect 95380 15506 95414 15574
rect 95482 15506 95516 15574
rect 96860 15506 96894 15888
rect 97332 15648 97366 15888
rect 97446 15800 97480 15888
rect 97492 15876 97493 15877
rect 97521 15876 97522 15877
rect 97491 15875 97492 15876
rect 97522 15875 97523 15876
rect 97534 15800 97568 15888
rect 97524 15750 97562 15788
rect 97490 15716 97562 15750
rect 97648 15648 97682 15888
rect 97332 15614 97682 15648
rect 97808 15648 97842 15888
rect 97922 15800 97956 15888
rect 98010 15882 98044 15888
rect 97968 15876 97969 15877
rect 97997 15876 97998 15877
rect 97967 15875 97968 15876
rect 97998 15875 97999 15876
rect 98004 15804 98044 15882
rect 98010 15800 98044 15804
rect 98000 15750 98038 15788
rect 97966 15716 98038 15750
rect 98124 15648 98158 15888
rect 97808 15614 98158 15648
rect 88271 15449 91727 15483
rect 93438 15472 96894 15506
rect 86748 15228 86760 15436
rect 86782 15262 86794 15436
rect 87166 15260 87556 15294
rect 87166 14762 87200 15260
rect 87295 15181 87427 15228
rect 87326 15169 87427 15181
rect 87342 15158 87427 15169
rect 87269 15099 87314 15110
rect 87397 15099 87442 15110
rect 87280 14923 87314 15099
rect 87408 14923 87442 15099
rect 87380 14864 87427 14911
rect 87342 14830 87427 14864
rect 87522 14762 87556 15260
rect 89016 15136 90368 15160
rect 87166 14728 87556 14762
rect 86366 14582 86774 14591
rect 86416 14572 86774 14582
rect 86818 14568 87018 14591
rect 86790 14557 87046 14563
rect 86332 14548 87046 14557
rect 86382 14540 87046 14548
rect 86382 14538 86808 14540
rect 87148 14058 87570 14678
rect 87714 14564 87974 14591
rect 87714 14536 87974 14563
rect 82640 13916 86670 13933
rect 86798 13916 87538 13933
rect 88174 13916 88986 13933
rect 90338 13916 90696 13933
rect 82668 13860 86726 13905
rect 86770 13899 87034 13905
rect 86766 13882 87572 13899
rect 88118 13860 88986 13905
rect 90338 13860 90668 13905
rect 90817 13847 90851 15449
rect 95380 13896 95414 15472
rect 100476 15402 100510 15888
rect 100562 15876 100650 15888
rect 100578 15500 100612 15876
rect 103554 15860 103626 15898
rect 103592 15484 103626 15860
rect 103554 15472 103642 15484
rect 100540 15410 100612 15448
rect 100662 15438 103642 15472
rect 103554 15426 103642 15438
rect 100476 15356 100572 15402
rect 100476 15264 100510 15356
rect 100566 15328 100572 15346
rect 100578 15276 100612 15410
rect 100618 15356 103586 15402
rect 100618 15328 103586 15346
rect 100622 15300 103586 15328
rect 103592 15292 103626 15426
rect 103632 15356 103664 15402
rect 103694 15346 103728 15964
rect 103632 15300 103728 15346
rect 100562 15268 100650 15276
rect 100540 15264 100650 15268
rect 103542 15264 103553 15275
rect 100442 15230 103553 15264
rect 95856 15188 96628 15202
rect 100476 14738 100510 15230
rect 100562 15218 100650 15230
rect 100578 14842 100612 15218
rect 103554 15202 103626 15240
rect 103592 14826 103626 15202
rect 103554 14814 103642 14826
rect 100540 14752 100612 14790
rect 100662 14780 103642 14814
rect 103554 14768 103642 14780
rect 100476 14698 100572 14738
rect 96572 14666 96628 14668
rect 96572 14566 96742 14612
rect 100476 14606 100510 14698
rect 100554 14642 100572 14682
rect 100578 14618 100612 14752
rect 100618 14698 103586 14738
rect 100618 14642 103586 14682
rect 103592 14634 103626 14768
rect 103632 14698 103668 14738
rect 103694 14682 103728 15300
rect 173352 14862 174866 14876
rect 173086 14824 173110 14846
rect 173064 14800 173110 14824
rect 181174 14824 181198 14846
rect 181174 14800 181220 14824
rect 103632 14642 103728 14682
rect 100562 14610 100650 14618
rect 100540 14606 100650 14610
rect 103542 14606 103553 14617
rect 100442 14572 103553 14606
rect 96572 14538 96742 14558
rect 100476 13948 100510 14572
rect 100562 14560 100650 14572
rect 100578 14184 100612 14560
rect 103554 14544 103626 14582
rect 103592 14168 103626 14544
rect 103554 14156 103642 14168
rect 100540 14094 100612 14132
rect 100662 14122 103642 14156
rect 103554 14110 103642 14122
rect 100532 14046 100572 14058
rect 100560 13990 100572 14030
rect 100578 13960 100612 14094
rect 100618 14046 103586 14058
rect 100618 13990 103586 14030
rect 103592 13976 103626 14110
rect 103632 14046 103664 14058
rect 103694 14030 103728 14642
rect 103632 13990 103728 14030
rect 100562 13952 100650 13960
rect 100540 13948 100650 13952
rect 103542 13948 103553 13959
rect 100442 13914 103553 13948
rect 100476 13834 100510 13914
rect 100547 13902 100650 13914
rect 103694 13834 103728 13990
rect 95476 13800 103728 13834
rect 100476 13446 100510 13800
rect 167986 13648 169166 14020
rect 104948 13548 105004 13560
rect 104948 13492 105004 13504
rect 173764 13372 173784 13430
rect 173792 13372 173812 13424
rect 99542 13296 99546 13330
rect 99576 13322 99580 13348
rect 100084 13126 100106 13132
rect 100084 13122 100102 13126
rect 100084 13066 100126 13076
rect 100181 13015 100234 13269
rect 173708 13132 174346 13372
rect 100435 12922 100488 13015
rect 101198 12966 101872 12979
rect 171436 12976 172316 13024
rect 100567 12945 101872 12966
rect 100471 12764 100505 12883
rect 100582 12803 101202 12945
rect 101252 12911 101786 12930
rect 171380 12920 172260 12968
rect 101286 12896 101784 12911
rect 100573 12764 101202 12803
rect 100471 12678 101202 12764
rect 85948 12318 85964 12348
rect 85914 12284 85930 12314
rect 100471 12281 100505 12678
rect 100573 12526 101202 12678
rect 101252 12871 101818 12877
rect 101252 12865 101286 12871
rect 101784 12865 101818 12871
rect 101252 12862 101818 12865
rect 101252 12790 101286 12862
rect 101409 12850 101661 12854
rect 101397 12831 101673 12850
rect 101623 12816 101634 12819
rect 101431 12801 101639 12816
rect 101307 12790 101388 12801
rect 101431 12797 101716 12801
rect 101252 12748 101292 12790
rect 101300 12754 101388 12790
rect 101447 12782 101634 12797
rect 101635 12754 101716 12797
rect 101300 12748 101320 12754
rect 101252 12574 101286 12748
rect 101354 12716 101388 12754
rect 101682 12716 101716 12754
rect 101623 12688 101634 12699
rect 101447 12654 101634 12688
rect 101784 12574 101818 12862
rect 173764 12800 173766 12976
rect 173792 12828 173794 12948
rect 174184 12860 174218 12932
rect 174184 12856 174214 12860
rect 174240 12832 174246 12960
rect 174240 12828 174242 12832
rect 101252 12540 101818 12574
rect 100573 12472 100607 12526
rect 100573 12281 101202 12472
rect 101252 12420 101818 12454
rect 101252 12281 101286 12420
rect 101623 12340 101634 12351
rect 101447 12315 101634 12340
rect 101431 12306 101639 12315
rect 101300 12281 101302 12300
rect 101784 12281 101818 12420
rect 174231 12304 174646 12335
rect 170678 12299 174646 12304
rect 179302 12304 179723 12335
rect 179302 12299 184662 12304
rect 95453 12248 103723 12281
rect 165607 12265 169443 12299
rect 170678 12270 184662 12299
rect 174231 12265 179723 12270
rect 95391 12247 103723 12248
rect 95391 12213 95426 12214
rect 100471 12167 100505 12247
rect 100573 12235 101202 12247
rect 100582 12205 101202 12235
rect 101252 12207 101286 12247
rect 101300 12213 101302 12247
rect 101354 12224 101388 12247
rect 101682 12241 101716 12247
rect 101674 12232 101726 12241
rect 101676 12228 101722 12232
rect 101682 12224 101716 12228
rect 101436 12219 101634 12223
rect 101447 12207 101623 12212
rect 101646 12207 101754 12213
rect 101784 12207 101818 12247
rect 101252 12205 101818 12207
rect 100582 12201 103566 12205
rect 100582 12179 103578 12201
rect 100526 12173 103578 12179
rect 100526 12167 101202 12173
rect 101252 12167 101286 12173
rect 101784 12167 101818 12173
rect 82694 12084 90670 12118
rect 95425 12028 95426 12155
rect 100437 12152 103544 12167
rect 100437 12139 103621 12152
rect 100437 12133 103539 12139
rect 95459 12028 95460 12121
rect 83940 10832 86906 11770
rect 87452 11504 89102 11774
rect 89538 11504 90892 11772
rect 93816 11596 93824 11622
rect 87452 11482 90892 11504
rect 79402 10534 79684 10558
rect 65104 10470 69072 10504
rect 75080 10499 80640 10504
rect 70313 10470 80640 10499
rect 65104 10402 68366 10470
rect 70313 10465 76625 10470
rect 68488 10408 68516 10434
rect 68658 10418 68669 10429
rect 68681 10418 68692 10429
rect 68658 10402 68692 10418
rect 65104 10368 68692 10402
rect 65104 10329 68366 10368
rect 68374 10329 68396 10334
rect 64244 6974 64252 7028
rect 64742 7010 64978 7264
rect 64738 6974 64978 7010
rect 65104 6974 68396 10329
rect 64063 6510 64092 6529
rect 62815 6438 62849 6486
rect 62815 6418 62860 6438
rect 62896 6418 63278 6486
rect 63279 6470 63337 6486
rect 63291 6438 63325 6470
rect 63291 6418 63336 6438
rect 63418 6418 63446 6480
rect 63473 6438 63507 6486
rect 63473 6418 63518 6438
rect 63542 6418 63754 6486
rect 63937 6470 63995 6486
rect 64032 6486 64092 6510
rect 64032 6484 64097 6486
rect 63980 6455 63995 6470
rect 63866 6430 63880 6436
rect 63866 6424 63943 6430
rect 63949 6418 63983 6452
rect 64063 6430 64097 6484
rect 64140 6436 64144 6480
rect 63989 6424 64144 6430
rect 64063 6418 64097 6424
rect 62633 6384 64156 6418
rect 64298 6408 64306 6974
rect 64738 6940 68396 6974
rect 64738 6872 64978 6940
rect 64988 6872 65035 6919
rect 64738 6838 65035 6872
rect 64738 6591 64978 6838
rect 65005 6779 65050 6790
rect 65016 6603 65050 6779
rect 64738 6565 65035 6591
rect 64738 6552 64978 6565
rect 64738 6534 64992 6552
rect 64738 6518 64988 6534
rect 65104 6518 68396 6940
rect 64738 6484 68396 6518
rect 62633 5906 62678 6384
rect 62710 6000 62738 6384
rect 62766 6000 62794 6384
rect 62815 5906 62860 6384
rect 62896 6050 63278 6384
rect 63291 5906 63336 6384
rect 63418 6000 63446 6384
rect 63473 5906 63518 6384
rect 63542 6274 63840 6384
rect 63542 6050 63754 6274
rect 61317 5346 61351 5906
rect 61499 5346 61533 5906
rect 61317 3531 61362 5346
rect 61378 3531 61406 4812
rect 61434 3531 61462 4812
rect 61499 3531 61544 5346
rect 61975 4422 62009 5906
rect 58029 3497 61617 3531
rect 58029 3429 58580 3497
rect 58772 3482 60254 3497
rect 60545 3482 60579 3497
rect 60659 3482 60704 3497
rect 60720 3482 60748 3497
rect 60776 3482 60804 3497
rect 60841 3482 60886 3497
rect 58772 3476 61262 3482
rect 61317 3476 61362 3497
rect 61378 3476 61406 3497
rect 61434 3476 61462 3497
rect 58772 3429 61488 3476
rect 58029 3427 60830 3429
rect 60841 3427 61488 3429
rect 58029 3395 61488 3427
rect 61499 3418 61544 3497
rect 54992 2217 55003 2228
rect 55015 2217 55026 2228
rect 58029 2190 58580 3395
rect 58772 3380 60898 3395
rect 61086 3380 61133 3395
rect 58772 3346 61133 3380
rect 58772 2930 60254 3346
rect 58718 2854 60254 2930
rect 58772 2368 60254 2854
rect 58772 2350 60304 2368
rect 58638 2316 60304 2350
rect 60545 2316 60579 3346
rect 60659 2328 60704 3346
rect 60800 3336 60886 3346
rect 60811 2328 60886 3336
rect 61103 3287 61148 3298
rect 60811 2316 60856 2328
rect 61114 2316 61148 3287
rect 58638 2269 60898 2316
rect 61102 2269 61161 2316
rect 61228 2269 61262 3395
rect 61317 2328 61351 3395
rect 61378 3074 61406 3389
rect 61370 2275 61406 3074
rect 61434 3347 61462 3389
rect 61499 3347 61533 3418
rect 61434 3336 61533 3347
rect 61434 3018 61462 3336
rect 61426 2316 61462 3018
rect 61469 2328 61533 3336
rect 61469 2316 61514 2328
rect 61426 2275 61515 2316
rect 61457 2269 61515 2275
rect 61583 2269 61617 3497
rect 61975 3418 62020 4422
rect 61975 2328 62009 3418
rect 62040 2275 62068 4812
rect 62096 2275 62124 4812
rect 62157 4422 62191 5906
rect 62633 4422 62667 5906
rect 62157 3418 62202 4422
rect 62633 3418 62678 4422
rect 62157 2328 62191 3418
rect 62633 2346 62667 3418
rect 62710 2346 62738 4812
rect 62766 2346 62794 4812
rect 62815 4422 62849 5906
rect 63291 4422 63325 5906
rect 62815 3418 62860 4422
rect 63291 3572 63336 4422
rect 63418 3572 63446 4812
rect 63473 4422 63507 5906
rect 63473 3572 63518 4422
rect 63587 3572 63621 6050
rect 64063 3572 64097 6384
rect 64284 6348 64288 6358
rect 64338 6218 64358 6454
rect 64366 6190 64386 6482
rect 64738 6476 64978 6484
rect 64434 6456 64554 6458
rect 64738 6456 65030 6476
rect 65104 6464 68396 6484
rect 65040 6456 68396 6464
rect 64738 6448 64978 6456
rect 64738 6442 65036 6448
rect 64406 6428 64582 6430
rect 64738 6416 65068 6442
rect 65104 6438 68396 6456
rect 68408 6438 68430 10368
rect 65104 6416 68407 6438
rect 64738 6382 68407 6416
rect 64738 6372 64978 6382
rect 65104 6358 68407 6382
rect 64760 6346 68407 6358
rect 65140 6226 65174 6346
rect 65282 6276 65294 6346
rect 65310 6304 65322 6346
rect 64458 6178 64534 6180
rect 64950 6178 64992 6200
rect 64430 6150 64562 6152
rect 64440 5928 64550 5948
rect 64478 5890 64512 5910
rect 65112 5870 65174 6226
rect 65284 6220 65294 6276
rect 65312 6248 65322 6304
rect 65348 6174 65386 6200
rect 65140 4792 65174 5870
rect 65616 4792 65650 6346
rect 65730 5906 65775 6346
rect 65806 6000 65834 6174
rect 65862 6000 65890 6174
rect 65912 5906 65957 6346
rect 65974 6030 66376 6346
rect 66164 6026 66376 6030
rect 66388 5906 66433 6346
rect 66458 6000 66486 6346
rect 66514 6000 66542 6346
rect 66570 5906 66615 6346
rect 66640 6030 67024 6346
rect 66640 6026 66852 6030
rect 67046 5906 67091 6346
rect 65730 4792 65764 5906
rect 65806 4792 65834 4812
rect 64304 4770 65872 4792
rect 64304 4766 65834 4770
rect 63100 3536 64133 3572
rect 65140 3536 65174 4766
rect 65616 3536 65650 4766
rect 65730 4422 65764 4766
rect 65730 3536 65775 4422
rect 65806 3536 65834 4766
rect 65912 4422 65946 5906
rect 66388 4422 66422 5906
rect 65912 3536 65957 4422
rect 66388 3536 66433 4422
rect 66458 3536 66486 4812
rect 66514 3536 66542 4812
rect 66570 4422 66604 5906
rect 67046 4422 67080 5906
rect 66570 3536 66615 4422
rect 63100 3502 66688 3536
rect 62815 2346 62849 3418
rect 63100 2346 64133 3502
rect 62502 2310 64133 2346
rect 64566 2310 64600 2344
rect 65140 2310 65174 3502
rect 65616 3472 65650 3502
rect 65730 3472 65775 3502
rect 65806 3472 65834 3502
rect 65912 3472 65957 3502
rect 66388 3472 66433 3502
rect 66458 3472 66486 3502
rect 66514 3472 66542 3502
rect 65190 3394 65208 3440
rect 65218 3366 65236 3468
rect 65250 3434 65892 3472
rect 65908 3434 66550 3472
rect 65254 3400 65892 3434
rect 65912 3400 66550 3434
rect 66570 3418 66615 3502
rect 65254 3362 65300 3400
rect 65254 3350 65288 3362
rect 65224 2326 65288 3350
rect 65224 2310 65258 2326
rect 65616 2310 65650 3400
rect 65730 2326 65764 3400
rect 65806 2310 65834 3394
rect 65912 3361 65946 3400
rect 65871 3350 65946 3361
rect 65882 2330 65946 3350
rect 65870 2326 65946 2330
rect 66388 2326 66422 3400
rect 66458 2770 66486 3394
rect 66514 3361 66542 3394
rect 66570 3361 66604 3418
rect 66514 2770 66604 3361
rect 66464 2358 66486 2770
rect 66492 2326 66604 2770
rect 65870 2310 65928 2326
rect 66492 2310 66586 2326
rect 66654 2310 66688 3502
rect 67046 3418 67091 4422
rect 67046 2326 67080 3418
rect 67116 2310 67144 6346
rect 67172 2342 67200 6346
rect 67228 5906 67273 6346
rect 67288 6030 67692 6346
rect 67480 6024 67692 6030
rect 67704 5906 67749 6346
rect 67228 4422 67262 5906
rect 67704 4422 67738 5906
rect 67228 3418 67273 4422
rect 67704 3418 67749 4422
rect 67228 2326 67262 3418
rect 67704 2326 67738 3418
rect 67780 2310 67808 6346
rect 67836 2310 67864 6346
rect 67886 5906 67931 6346
rect 67956 6024 68336 6346
rect 68124 6012 68336 6024
rect 68362 5906 68407 6346
rect 67886 4422 67920 5906
rect 68362 4422 68396 5906
rect 68408 5870 68430 5906
rect 67886 3418 67931 4422
rect 68362 3418 68407 4422
rect 67886 2342 67920 3418
rect 68362 2342 68396 3418
rect 67886 2326 67892 2342
rect 62502 2298 67864 2310
rect 68488 2298 68516 10362
rect 68533 10318 68589 10329
rect 68544 5870 68589 10318
rect 68544 4422 68578 5870
rect 68544 3418 68589 4422
rect 68544 2342 68578 3418
rect 62502 2292 67858 2298
rect 68658 2292 68692 10368
rect 70217 3788 70251 10403
rect 73037 10397 73071 10435
rect 73735 10413 73746 10424
rect 73758 10413 73769 10424
rect 73735 10397 73769 10413
rect 73037 10363 73769 10397
rect 72970 6782 72997 10320
rect 73004 6816 73031 10354
rect 70181 3632 70268 3788
rect 70312 3632 70386 3698
rect 70148 3556 70386 3632
rect 69058 3536 69066 3552
rect 69036 3518 69066 3536
rect 70181 3534 70268 3556
rect 69076 3518 69204 3534
rect 69552 3518 69792 3534
rect 70028 3518 70268 3534
rect 70312 3532 70386 3556
rect 69036 3482 69204 3518
rect 70217 3498 70251 3518
rect 70312 3498 70392 3532
rect 69208 3482 69406 3498
rect 69684 3482 69882 3498
rect 70160 3482 70454 3498
rect 69054 3448 71410 3482
rect 69054 3299 69204 3448
rect 70217 3430 70251 3448
rect 70312 3434 70386 3448
rect 70298 3430 70386 3434
rect 69238 3418 69376 3430
rect 69714 3418 69852 3430
rect 70217 3418 70386 3430
rect 69272 3384 69342 3396
rect 69288 3380 69326 3384
rect 69468 3380 69502 3418
rect 69266 3353 69502 3380
rect 69250 3346 69502 3353
rect 69390 3340 69422 3343
rect 69428 3340 69502 3346
rect 69226 3315 69260 3319
rect 69354 3315 69388 3319
rect 69214 3299 69222 3315
rect 69226 3312 69272 3315
rect 69235 3303 69272 3312
rect 69054 3287 69222 3299
rect 69226 3299 69272 3303
rect 69342 3299 69400 3315
rect 69226 3287 69260 3299
rect 69054 3127 69260 3287
rect 69354 3127 69388 3299
rect 69054 3104 69238 3127
rect 69054 2972 69244 3104
rect 69246 3000 69272 3076
rect 69326 3068 69373 3115
rect 69288 3034 69373 3068
rect 69246 2980 69366 3000
rect 69054 2966 69394 2972
rect 69428 2966 69440 2972
rect 69468 2966 69502 3340
rect 69054 2932 69502 2966
rect 69588 3380 69622 3418
rect 69748 3384 69818 3396
rect 69764 3380 69802 3384
rect 69944 3380 69978 3418
rect 69588 3346 69978 3380
rect 69588 2966 69622 3346
rect 69702 3315 69736 3319
rect 69830 3315 69864 3319
rect 69690 3299 69748 3315
rect 69818 3299 69876 3315
rect 69702 3127 69736 3299
rect 69830 3127 69864 3299
rect 69802 3068 69849 3115
rect 69764 3034 69849 3068
rect 69944 2966 69978 3346
rect 69588 2932 69978 2966
rect 70064 2966 70098 3418
rect 70217 3396 70251 3418
rect 70270 3402 70286 3406
rect 70270 3398 70290 3402
rect 70298 3398 70386 3418
rect 70217 3384 70294 3396
rect 70217 3380 70278 3384
rect 70312 3380 70386 3398
rect 70420 3427 70454 3448
rect 70983 3427 71029 3448
rect 70420 3380 70467 3427
rect 70955 3396 70978 3398
rect 70983 3396 71036 3427
rect 70955 3386 71036 3396
rect 70977 3380 71036 3386
rect 71234 3380 71281 3427
rect 70217 3353 71281 3380
rect 70144 3346 71281 3353
rect 70178 3315 70212 3319
rect 70217 3315 70251 3346
rect 70312 3319 70386 3346
rect 70306 3315 70386 3319
rect 70166 3299 70251 3315
rect 70294 3299 70386 3315
rect 70178 3127 70212 3299
rect 70183 3111 70212 3127
rect 70217 3068 70251 3299
rect 70306 3127 70386 3299
rect 70312 3115 70386 3127
rect 70278 3068 70386 3115
rect 70217 3044 70386 3068
rect 70217 3034 70325 3044
rect 70217 2966 70251 3034
rect 70331 3000 70365 3044
rect 70331 2966 70392 3000
rect 70420 2966 70454 3346
rect 70977 3340 71035 3346
rect 70064 2932 70454 2966
rect 70955 3299 71035 3340
rect 70955 2960 70978 3299
rect 70983 2960 71029 3299
rect 71251 3287 71296 3298
rect 69054 2882 69222 2932
rect 69428 2914 69440 2932
rect 69428 2882 69442 2914
rect 70217 2882 70251 2932
rect 70331 2882 70365 2932
rect 62502 2276 68992 2292
rect 62502 2269 64133 2276
rect 58638 2258 64133 2269
rect 55088 2176 58580 2190
rect 58734 2180 58740 2258
rect 58772 2235 64133 2258
rect 30850 1792 30870 2158
rect 31220 2142 39219 2176
rect 40320 2156 58580 2176
rect 40320 2142 57916 2156
rect 31372 1982 32854 2142
rect 31432 882 31466 1982
rect 31506 882 31540 1982
rect 31620 882 31665 1982
rect 32090 882 32135 1982
rect 32204 1792 32238 1982
rect 32204 1682 32256 1792
rect 32204 882 32238 1682
rect 32278 882 32312 1982
rect 33554 1792 33566 2142
rect 28650 877 34956 882
rect 23717 848 34956 877
rect 23717 843 30023 848
rect 22456 -3470 22464 -3416
rect 23579 -3434 23666 -3180
rect 22474 -4072 22602 -3434
rect 22612 -3853 22620 -3653
rect 22950 -3968 23190 -3434
rect 23426 -3470 23666 -3434
rect 23729 -3470 23763 843
rect 24387 822 24421 843
rect 25045 822 25079 843
rect 25703 822 25737 843
rect 26361 822 26395 843
rect 24359 775 24421 822
rect 25017 775 25079 822
rect 25675 775 25737 822
rect 26333 775 26395 822
rect 26435 822 26469 843
rect 26549 840 26594 843
rect 27019 840 27064 843
rect 26549 822 26583 840
rect 27019 822 27053 840
rect 26435 775 26482 822
rect 26549 775 26596 822
rect 27019 775 27066 822
rect 27133 775 27167 843
rect 27207 822 27241 843
rect 27179 775 27241 822
rect 27831 822 27846 843
rect 27859 822 27902 843
rect 28523 822 28557 843
rect 27831 809 27902 822
rect 28495 809 28557 822
rect 27831 775 27905 809
rect 27915 775 27933 781
rect 28495 775 28572 809
rect 28573 775 28600 781
rect 28650 780 30023 843
rect 30116 818 30150 848
rect 30774 818 30808 848
rect 31432 818 31466 848
rect 31506 818 31540 848
rect 31620 818 31665 848
rect 32090 818 32135 848
rect 32204 818 32238 848
rect 32278 818 32312 848
rect 32936 818 32970 848
rect 33594 818 33628 848
rect 34252 818 34286 848
rect 34910 818 34944 848
rect 30088 814 30150 818
rect 30746 814 30808 818
rect 30088 786 30156 814
rect 30746 786 30814 814
rect 30082 780 30156 786
rect 30166 780 30184 786
rect 30740 780 30814 786
rect 30824 780 30842 786
rect 31220 780 34944 818
rect 28650 775 30156 780
rect 23775 741 24421 775
rect 24433 741 25079 775
rect 25091 741 25737 775
rect 25749 741 26395 775
rect 26407 741 27241 775
rect 27253 741 27905 775
rect 27911 746 30156 775
rect 30162 746 30814 780
rect 30820 746 31472 780
rect 27911 741 30023 746
rect 23426 -3504 23852 -3470
rect 22644 -3988 22764 -3968
rect 22950 -3988 23240 -3968
rect 23426 -3986 23666 -3504
rect 23696 -3538 23712 -3534
rect 23668 -3566 23684 -3562
rect 23668 -3612 23688 -3566
rect 23668 -3614 23684 -3612
rect 23696 -3640 23716 -3538
rect 23717 -3606 23723 -3525
rect 23696 -3642 23712 -3640
rect 23729 -3665 23763 -3504
rect 23704 -3841 23763 -3665
rect 23710 -3924 23714 -3898
rect 23717 -3934 23723 -3853
rect 23426 -3988 23696 -3986
rect 22950 -3996 23190 -3988
rect 22638 -4016 22792 -3996
rect 22950 -4016 23268 -3996
rect 23290 -4014 23314 -3996
rect 23426 -4002 23666 -3988
rect 23729 -4002 23763 -3841
rect 23818 -4002 23852 -3504
rect 23318 -4014 23342 -4008
rect 22950 -4072 23190 -4016
rect 23426 -4036 23852 -4002
rect 23426 -4072 23666 -4036
rect 22532 -4218 22566 -4072
rect 23615 -4086 23649 -4072
rect 23729 -4086 23763 -4036
rect 22528 -4574 22566 -4218
rect 22608 -4270 22798 -4268
rect 22636 -4298 22682 -4296
rect 22724 -4298 22770 -4296
rect 22144 -4676 22452 -4638
rect 18698 -4710 22452 -4676
rect 18702 -4716 18720 -4710
rect 18652 -4778 18686 -4744
rect 19014 -4778 19048 -4710
rect 19116 -4726 19174 -4710
rect 19128 -4774 19162 -4726
rect 19128 -4778 19173 -4774
rect 19204 -4778 19232 -4716
rect 19310 -4774 19344 -4710
rect 19774 -4726 19832 -4710
rect 19786 -4774 19820 -4726
rect 19310 -4778 19355 -4774
rect 19786 -4778 19831 -4774
rect 19856 -4778 19884 -4716
rect 19912 -4778 19940 -4716
rect 19968 -4774 20002 -4710
rect 20432 -4726 20490 -4710
rect 20444 -4774 20478 -4726
rect 19968 -4778 20013 -4774
rect 20444 -4778 20489 -4774
rect 20514 -4778 20542 -4716
rect 20570 -4778 20598 -4716
rect 20626 -4774 20660 -4710
rect 21090 -4726 21148 -4710
rect 21102 -4774 21136 -4726
rect 20626 -4778 20671 -4774
rect 21102 -4778 21147 -4774
rect 21178 -4778 21206 -4716
rect 21234 -4778 21262 -4716
rect 21284 -4774 21318 -4710
rect 21748 -4726 21806 -4710
rect 21760 -4774 21794 -4726
rect 21284 -4778 21329 -4774
rect 21760 -4778 21805 -4774
rect 21886 -4778 21914 -4716
rect 21942 -4774 21976 -4710
rect 21942 -4778 21987 -4774
rect 22056 -4778 22090 -4710
rect 22384 -4716 22402 -4710
rect 22412 -4744 22452 -4710
rect 22418 -4778 22452 -4744
rect 18634 -4812 22486 -4778
rect 19014 -7330 19048 -4812
rect 19128 -5874 19173 -4812
rect 19204 -5180 19232 -4812
rect 19310 -5874 19355 -4812
rect 19680 -5622 19684 -5302
rect 19718 -5622 19722 -5302
rect 19786 -5874 19831 -4812
rect 19856 -5180 19884 -4812
rect 19912 -5180 19940 -4812
rect 19968 -5874 20013 -4812
rect 20444 -5874 20489 -4812
rect 20514 -5180 20542 -4812
rect 20570 -5180 20598 -4812
rect 20626 -5874 20671 -4812
rect 21102 -5686 21147 -4812
rect 21178 -5180 21206 -4812
rect 21234 -5180 21262 -4812
rect 21284 -5686 21329 -4812
rect 19128 -7280 19162 -5874
rect 19204 -7280 19232 -6368
rect 19310 -7280 19344 -5874
rect 19786 -7280 19820 -5874
rect 19856 -7264 19884 -6368
rect 19912 -7264 19940 -6368
rect 19968 -7280 20002 -5874
rect 20444 -7280 20478 -5874
rect 20514 -7324 20542 -6368
rect 20570 -7280 20598 -6368
rect 20626 -7280 20660 -5874
rect 21102 -7280 21136 -5686
rect 21178 -7324 21206 -6368
rect 21234 -7324 21262 -6368
rect 21284 -7280 21318 -5686
rect 21760 -5712 21805 -4812
rect 21886 -5180 21914 -4812
rect 21942 -5712 21987 -4812
rect 21760 -7280 21794 -5712
rect 21830 -6564 21858 -6368
rect 21886 -7324 21914 -6368
rect 21942 -7280 21976 -5712
rect 22056 -7330 22090 -4812
rect 22456 -6124 22464 -6070
rect 22532 -6088 22566 -4574
rect 23579 -4699 23866 -4086
rect 24387 -4652 24421 741
rect 25045 -4652 25079 741
rect 25703 -4652 25737 741
rect 26361 -4652 26395 741
rect 24359 -4665 24421 -4652
rect 25017 -4665 25079 -4652
rect 25675 -4665 25737 -4652
rect 26333 -4665 26395 -4652
rect 24359 -4693 24427 -4665
rect 25017 -4693 25085 -4665
rect 25675 -4693 25743 -4665
rect 26333 -4693 26401 -4665
rect 24353 -4699 24427 -4693
rect 24437 -4699 24455 -4693
rect 25011 -4699 25085 -4693
rect 25095 -4699 25113 -4693
rect 25669 -4699 25743 -4693
rect 25753 -4699 25771 -4693
rect 26327 -4699 26401 -4693
rect 26411 -4699 26429 -4693
rect 26435 -4699 26469 741
rect 26549 -4652 26583 741
rect 26768 -470 26980 -462
rect 26612 -910 26980 -470
rect 26612 -918 26824 -910
rect 26768 -3124 26980 -3116
rect 26612 -3564 26980 -3124
rect 26612 -3572 26824 -3564
rect 27019 -4652 27053 741
rect 27133 388 27167 741
rect 27133 -964 27170 388
rect 26537 -4699 26596 -4652
rect 27019 -4699 27066 -4652
rect 27133 -4699 27167 -964
rect 27207 -4652 27241 741
rect 27831 735 27849 741
rect 27831 600 27846 735
rect 27859 707 27905 741
rect 27915 735 27933 741
rect 28523 707 28572 741
rect 28573 735 28600 741
rect 27859 544 27902 707
rect 27865 6 27899 544
rect 27844 -28 28234 6
rect 27844 -526 27878 -28
rect 28058 -96 28105 -49
rect 28020 -130 28105 -96
rect 27947 -189 27992 -178
rect 28075 -189 28120 -178
rect 27958 -360 27992 -189
rect 27924 -365 27992 -360
rect 28086 -365 28120 -189
rect 27924 -368 27986 -365
rect 27952 -377 27986 -368
rect 27896 -433 27905 -377
rect 27980 -433 27986 -416
rect 28058 -424 28105 -377
rect 28020 -458 28105 -424
rect 28078 -462 28084 -458
rect 28090 -498 28096 -462
rect 28200 -526 28234 -28
rect 27256 -562 27260 -550
rect 27844 -560 28234 -526
rect 27268 -590 27272 -562
rect 27830 -1230 28252 -610
rect 28523 -1226 28557 707
rect 28458 -1312 28557 -1226
rect 28523 -2176 28557 -1312
rect 28600 196 28602 394
rect 28600 -378 28618 196
rect 28600 -1372 28602 -378
rect 28650 -504 30023 741
rect 30082 740 30100 746
rect 30110 712 30156 746
rect 30166 740 30184 746
rect 30740 740 30758 746
rect 30768 712 30814 746
rect 30824 740 30842 746
rect 31398 740 31416 746
rect 31426 712 31472 746
rect 31482 746 32318 780
rect 31482 740 31500 746
rect 28650 -760 30032 -504
rect 30046 -732 30088 -532
rect 28650 -2176 30023 -760
rect 27850 -2202 30023 -2176
rect 27844 -2682 28234 -2648
rect 27844 -3180 27878 -2682
rect 28058 -2750 28105 -2703
rect 28020 -2784 28105 -2750
rect 27947 -2843 27992 -2832
rect 28075 -2843 28120 -2832
rect 27958 -3019 27992 -2843
rect 28086 -3019 28120 -2843
rect 27924 -3059 27932 -3022
rect 27952 -3031 27960 -3022
rect 28058 -3078 28105 -3031
rect 28020 -3112 28105 -3078
rect 28078 -3116 28084 -3112
rect 28090 -3152 28096 -3116
rect 28200 -3180 28234 -2682
rect 28408 -3174 28434 -3032
rect 28436 -3174 28462 -3032
rect 27844 -3214 28234 -3180
rect 27830 -3884 28252 -3264
rect 28408 -3478 28434 -3374
rect 28436 -3478 28462 -3374
rect 28523 -3880 28557 -2202
rect 28600 -3032 28618 -2458
rect 28650 -3158 30023 -2202
rect 28650 -3414 30032 -3158
rect 30074 -3186 30088 -2934
rect 30046 -3216 30088 -3186
rect 30116 -3216 30150 712
rect 30774 42 30808 712
rect 30628 -496 31090 42
rect 30628 -562 31238 -496
rect 30628 -596 31300 -562
rect 30750 -646 30842 -596
rect 31026 -638 31300 -596
rect 31026 -646 31238 -638
rect 30686 -680 31238 -646
rect 30686 -1160 30720 -680
rect 30750 -710 30880 -680
rect 30750 -720 30916 -710
rect 30774 -832 30808 -720
rect 30828 -768 30916 -720
rect 30828 -782 30842 -768
rect 30844 -782 30916 -768
rect 30878 -790 30900 -786
rect 30820 -832 30834 -821
rect 30774 -1008 30834 -832
rect 30854 -990 30870 -792
rect 30906 -818 30928 -786
rect 30882 -821 30898 -820
rect 30877 -832 30922 -821
rect 30882 -1008 30922 -832
rect 31002 -944 31238 -680
rect 31398 -720 31402 -520
rect 31426 -748 31430 -492
rect 31432 -796 31466 712
rect 30774 -1022 30808 -1008
rect 30882 -1018 30898 -1008
rect 30878 -1022 30916 -1020
rect 30774 -1136 30814 -1022
rect 30828 -1108 30842 -1050
rect 30878 -1058 30922 -1022
rect 30844 -1092 30922 -1058
rect 30878 -1108 30894 -1092
rect 30906 -1136 30922 -1092
rect 30774 -1160 30808 -1136
rect 31002 -1160 31036 -944
rect 30686 -1194 31036 -1160
rect 30774 -2612 30808 -1194
rect 31398 -1372 31422 -824
rect 31426 -1400 31466 -796
rect 30878 -2174 30880 -1974
rect 30906 -2202 30908 -1946
rect 30628 -3150 31090 -2612
rect 30628 -3216 31238 -3150
rect 31368 -3174 31394 -3032
rect 31396 -3174 31422 -3032
rect 30046 -3348 30206 -3216
rect 30628 -3250 31300 -3216
rect 31026 -3292 31300 -3250
rect 31026 -3300 31238 -3292
rect 30686 -3334 31238 -3300
rect 30046 -3386 30088 -3348
rect 27844 -3924 27918 -3884
rect 27865 -4652 27899 -3924
rect 28458 -3966 28557 -3880
rect 27179 -4665 27241 -4652
rect 27179 -4693 27247 -4665
rect 27837 -4693 27899 -4652
rect 28408 -4693 28434 -4026
rect 28436 -4693 28462 -4026
rect 28523 -4652 28557 -3966
rect 28600 -4026 28602 -3478
rect 27173 -4699 27247 -4693
rect 27257 -4699 27275 -4693
rect 27831 -4699 27899 -4693
rect 28495 -4699 28557 -4652
rect 28650 -4676 30023 -3414
rect 30074 -4336 30088 -3386
rect 30098 -3936 30172 -3348
rect 30686 -3814 30720 -3334
rect 30774 -3440 30808 -3334
rect 30878 -3402 30916 -3364
rect 30828 -3436 30842 -3402
rect 30844 -3436 30916 -3402
rect 30774 -3472 30814 -3440
rect 30824 -3444 30842 -3440
rect 30878 -3444 30900 -3440
rect 30906 -3472 30928 -3440
rect 30774 -3486 30808 -3472
rect 30820 -3486 30834 -3475
rect 30877 -3486 30922 -3475
rect 30774 -3662 30834 -3486
rect 30888 -3662 30922 -3486
rect 31002 -3598 31238 -3334
rect 31368 -3478 31394 -3374
rect 31396 -3478 31422 -3374
rect 30774 -3814 30808 -3662
rect 30878 -3676 30918 -3674
rect 30878 -3712 30922 -3676
rect 30828 -3746 30842 -3712
rect 30844 -3746 30922 -3712
rect 30878 -3762 30894 -3746
rect 30878 -3774 30890 -3762
rect 30906 -3790 30922 -3746
rect 30906 -3802 30918 -3790
rect 31002 -3814 31036 -3598
rect 30686 -3848 31036 -3814
rect 30116 -4638 30150 -3936
rect 30774 -4638 30808 -3848
rect 31398 -4026 31420 -3808
rect 31368 -4400 31394 -4026
rect 31396 -4372 31422 -4026
rect 30088 -4642 30150 -4638
rect 30088 -4670 30156 -4642
rect 30082 -4676 30156 -4670
rect 30166 -4676 30184 -4670
rect 30746 -4676 30808 -4638
rect 30878 -4670 30880 -4628
rect 30906 -4670 30908 -4600
rect 31432 -4638 31466 -1400
rect 31502 -4372 31504 -2970
rect 31404 -4642 31466 -4638
rect 31404 -4670 31472 -4642
rect 31398 -4676 31472 -4670
rect 31482 -4676 31500 -4670
rect 31506 -4676 31540 746
rect 31620 600 31665 746
rect 32090 600 32135 746
rect 31620 -3254 31654 600
rect 32090 -274 32124 600
rect 32204 132 32238 746
rect 32244 740 32262 746
rect 32272 712 32318 746
rect 32328 746 32976 780
rect 32328 740 32346 746
rect 32902 740 32920 746
rect 32930 712 32976 746
rect 32986 746 33634 780
rect 32986 740 33004 746
rect 33560 740 33578 746
rect 33588 712 33634 746
rect 33644 746 34292 780
rect 33644 740 33662 746
rect 34218 740 34236 746
rect 34246 712 34292 746
rect 34302 746 34944 780
rect 34302 740 34320 746
rect 34876 740 34894 746
rect 34904 712 34944 746
rect 32066 -490 32158 -274
rect 31864 -508 32158 -490
rect 31670 -732 32158 -508
rect 31670 -938 32076 -732
rect 31670 -956 31882 -938
rect 31864 -3162 32076 -3144
rect 31670 -3254 32076 -3162
rect 31604 -3592 32076 -3254
rect 31604 -3610 31882 -3592
rect 31604 -3908 31678 -3610
rect 31620 -4638 31654 -3908
rect 32090 -4638 32124 -732
rect 32204 -972 32256 132
rect 31608 -4676 31666 -4638
rect 32090 -4676 32128 -4638
rect 32204 -4676 32238 -972
rect 32278 -4638 32312 712
rect 32936 0 32970 712
rect 32326 -3460 32350 -3378
rect 32622 -4072 33084 -3434
rect 33098 -4072 33560 -3434
rect 32936 -4122 32970 -4072
rect 32676 -4156 33026 -4122
rect 32676 -4636 32710 -4156
rect 32868 -4224 32906 -4186
rect 32834 -4258 32906 -4224
rect 32866 -4266 32888 -4262
rect 32779 -4308 32824 -4297
rect 32844 -4300 32852 -4270
rect 32894 -4294 32916 -4262
rect 32872 -4297 32880 -4296
rect 32902 -4297 32912 -4294
rect 32867 -4308 32912 -4297
rect 32790 -4484 32824 -4308
rect 32878 -4484 32912 -4308
rect 32902 -4496 32912 -4484
rect 32868 -4500 32912 -4496
rect 32868 -4534 32906 -4500
rect 32834 -4568 32906 -4534
rect 32936 -4636 32970 -4156
rect 32992 -4636 33026 -4156
rect 32676 -4638 33026 -4636
rect 33152 -4156 33502 -4122
rect 33152 -4636 33186 -4156
rect 33344 -4224 33382 -4186
rect 33310 -4258 33382 -4224
rect 33255 -4308 33300 -4297
rect 33343 -4308 33388 -4297
rect 33266 -4484 33300 -4308
rect 33354 -4484 33388 -4308
rect 33344 -4534 33382 -4496
rect 33310 -4568 33382 -4534
rect 33468 -4636 33502 -4156
rect 33152 -4638 33502 -4636
rect 33594 -4638 33628 712
rect 34252 -4638 34286 712
rect 34910 -4638 34944 712
rect 32250 -4670 33506 -4638
rect 33566 -4642 33628 -4638
rect 34224 -4642 34286 -4638
rect 33566 -4670 33634 -4642
rect 34224 -4670 34292 -4642
rect 34882 -4670 34944 -4638
rect 32244 -4676 33506 -4670
rect 33560 -4676 33634 -4670
rect 33644 -4676 33662 -4670
rect 34218 -4676 34292 -4670
rect 34302 -4676 34320 -4670
rect 34876 -4676 34944 -4670
rect 28650 -4699 30156 -4676
rect 23579 -4706 24427 -4699
rect 23615 -5834 23649 -4706
rect 23751 -4767 23769 -4706
rect 23779 -4733 24427 -4706
rect 24433 -4733 25085 -4699
rect 25091 -4733 25743 -4699
rect 25749 -4733 26401 -4699
rect 26407 -4733 27247 -4699
rect 27253 -4733 27899 -4699
rect 27911 -4733 28557 -4699
rect 28569 -4710 30156 -4699
rect 30162 -4710 30808 -4676
rect 30820 -4710 31472 -4676
rect 31478 -4710 32312 -4676
rect 32340 -4710 32976 -4676
rect 28569 -4733 30023 -4710
rect 30082 -4716 30100 -4710
rect 23779 -4739 23797 -4733
rect 24353 -4739 24371 -4733
rect 24381 -4767 24427 -4733
rect 24437 -4739 24455 -4733
rect 25011 -4739 25029 -4733
rect 25039 -4767 25085 -4733
rect 25095 -4739 25113 -4733
rect 25669 -4739 25687 -4733
rect 23729 -4801 23763 -4767
rect 24387 -4801 24421 -4767
rect 25045 -4801 25079 -4767
rect 25166 -4801 25188 -4744
rect 25697 -4767 25743 -4733
rect 25753 -4739 25771 -4733
rect 26327 -4739 26345 -4733
rect 26355 -4767 26401 -4733
rect 26411 -4739 26429 -4733
rect 25703 -4801 25737 -4767
rect 26361 -4801 26395 -4767
rect 26435 -4801 26469 -4733
rect 26537 -4749 26595 -4733
rect 26549 -4801 26583 -4749
rect 27019 -4801 27053 -4733
rect 27133 -4801 27167 -4733
rect 27173 -4739 27191 -4733
rect 27201 -4767 27247 -4733
rect 27257 -4739 27275 -4733
rect 27831 -4739 27849 -4733
rect 27859 -4767 27899 -4733
rect 27207 -4801 27241 -4767
rect 27865 -4801 27899 -4767
rect 28408 -4801 28434 -4739
rect 28436 -4801 28462 -4739
rect 28523 -4801 28557 -4733
rect 28650 -4778 30023 -4733
rect 30110 -4744 30156 -4710
rect 30166 -4716 30184 -4710
rect 30116 -4778 30150 -4744
rect 30774 -4778 30808 -4710
rect 31398 -4716 31416 -4710
rect 30878 -4778 30880 -4716
rect 30906 -4778 30908 -4716
rect 31426 -4744 31472 -4710
rect 31482 -4716 31500 -4710
rect 31432 -4778 31466 -4744
rect 31506 -4778 31540 -4710
rect 31608 -4726 31666 -4710
rect 31620 -4774 31654 -4726
rect 32090 -4774 32124 -4710
rect 31620 -4778 31665 -4774
rect 32090 -4778 32135 -4774
rect 32204 -4778 32238 -4710
rect 32244 -4716 32262 -4710
rect 32272 -4744 32312 -4710
rect 32278 -4778 32312 -4744
rect 32348 -4778 32350 -4710
rect 32898 -4778 32910 -4710
rect 32936 -4744 32976 -4710
rect 32986 -4710 33634 -4676
rect 33640 -4710 34292 -4676
rect 34298 -4710 34944 -4676
rect 32986 -4716 33004 -4710
rect 33560 -4716 33578 -4710
rect 33588 -4744 33634 -4710
rect 33644 -4716 33662 -4710
rect 34218 -4716 34236 -4710
rect 34246 -4744 34292 -4710
rect 34302 -4716 34320 -4710
rect 34876 -4716 34894 -4710
rect 34904 -4744 34944 -4710
rect 32936 -4778 32970 -4744
rect 33594 -4778 33628 -4744
rect 34252 -4778 34286 -4744
rect 34378 -4778 34384 -4744
rect 34910 -4778 34944 -4744
rect 28650 -4801 34978 -4778
rect 23711 -4812 34978 -4801
rect 23711 -4835 30023 -4812
rect 30878 -4828 30880 -4812
rect 23579 -6088 23666 -5834
rect 22474 -6726 22602 -6088
rect 22612 -6507 22620 -6307
rect 22950 -6622 23190 -6088
rect 23426 -6124 23666 -6088
rect 23729 -6124 23790 -6090
rect 23426 -6158 23852 -6124
rect 22644 -6642 22764 -6622
rect 22950 -6642 23240 -6622
rect 23426 -6640 23666 -6158
rect 23717 -6260 23723 -6179
rect 23729 -6319 23763 -6158
rect 23704 -6495 23763 -6319
rect 23710 -6578 23714 -6552
rect 23717 -6588 23723 -6507
rect 23729 -6622 23763 -6495
rect 23426 -6642 23696 -6640
rect 22950 -6650 23190 -6642
rect 22638 -6670 22792 -6650
rect 22950 -6670 23268 -6650
rect 23290 -6668 23314 -6650
rect 23426 -6656 23666 -6642
rect 23729 -6656 23790 -6622
rect 23818 -6656 23852 -6158
rect 23318 -6668 23342 -6662
rect 22950 -6726 23190 -6670
rect 23426 -6690 23852 -6656
rect 23426 -6726 23666 -6690
rect 22532 -6872 22566 -6726
rect 23615 -6740 23649 -6726
rect 22528 -7228 22566 -6872
rect 22608 -6924 22798 -6922
rect 22636 -6952 22682 -6950
rect 22724 -6952 22770 -6950
rect 19014 -7364 22390 -7330
rect 19014 -7380 19048 -7364
rect 20514 -7376 20542 -7370
rect 19014 -7391 19025 -7380
rect 19037 -7391 19048 -7380
rect 21178 -7382 21206 -7370
rect 21234 -7376 21262 -7370
rect 21886 -7382 21914 -7370
rect 22056 -7380 22090 -7364
rect 22532 -7370 22566 -7228
rect 23579 -7360 23866 -6740
rect 25045 -7294 25079 -4835
rect 25166 -5178 25188 -4835
rect 25330 -5024 25720 -4990
rect 25330 -5522 25364 -5024
rect 25544 -5092 25591 -5045
rect 25506 -5126 25591 -5092
rect 25686 -5052 25720 -5024
rect 25433 -5185 25478 -5174
rect 25561 -5185 25606 -5174
rect 25444 -5361 25478 -5185
rect 25572 -5361 25606 -5185
rect 25544 -5420 25591 -5373
rect 25506 -5454 25591 -5420
rect 25686 -5460 25754 -5052
rect 25686 -5522 25720 -5460
rect 25330 -5556 25720 -5522
rect 25312 -6116 25734 -5606
rect 25312 -6226 25736 -6116
rect 25669 -6368 25702 -6226
rect 25703 -6402 25736 -6226
rect 26435 -7353 26469 -4835
rect 26549 -7294 26583 -4835
rect 27019 -7294 27053 -4835
rect 27133 -7353 27167 -4835
rect 28408 -5180 28434 -4835
rect 28436 -5180 28462 -4835
rect 27844 -6254 27918 -5924
rect 27768 -6484 27772 -6368
rect 27844 -6408 28050 -6254
rect 27844 -6578 27918 -6408
rect 28408 -7347 28434 -6368
rect 28436 -6428 28490 -6368
rect 28436 -7347 28462 -6428
rect 28523 -7294 28557 -4835
rect 22056 -7391 22067 -7380
rect 22079 -7391 22090 -7380
rect 16985 -7414 16996 -7403
rect 17008 -7414 17019 -7403
rect 13563 -7489 17399 -7455
rect 18634 -7466 22470 -7432
rect 25040 -7455 26010 -7354
rect 26435 -7387 27167 -7353
rect 26435 -7403 26469 -7387
rect 26435 -7414 26446 -7403
rect 26458 -7414 26469 -7403
rect 27133 -7403 27167 -7387
rect 28408 -7400 28434 -7393
rect 27133 -7414 27144 -7403
rect 27156 -7414 27167 -7403
rect 28436 -7428 28462 -7393
rect 28650 -7432 30023 -4835
rect 30906 -4856 30908 -4812
rect 30074 -6990 30088 -6368
rect 30878 -6428 30890 -6368
rect 30906 -6484 30946 -6368
rect 31368 -7054 31394 -6368
rect 31396 -7026 31422 -6368
rect 31502 -7026 31504 -6368
rect 31506 -7330 31540 -4812
rect 31620 -5874 31665 -4812
rect 32090 -5874 32135 -4812
rect 31620 -7280 31654 -5874
rect 32090 -7280 32124 -5874
rect 32204 -7330 32238 -4812
rect 32278 -7262 32312 -4812
rect 32936 -4826 32948 -4812
rect 34252 -4898 34286 -4812
rect 34194 -4980 34286 -4898
rect 32326 -6114 32350 -6032
rect 32622 -6726 33084 -6088
rect 33098 -6726 33560 -6088
rect 33726 -6554 33738 -6368
rect 32936 -6776 32964 -6742
rect 32676 -6810 33026 -6776
rect 32278 -7280 32326 -7262
rect 32312 -7284 32326 -7280
rect 32676 -7290 32710 -6810
rect 32868 -6878 32906 -6840
rect 32834 -6912 32906 -6878
rect 32866 -6920 32888 -6916
rect 32779 -6962 32824 -6951
rect 32844 -6954 32852 -6924
rect 32894 -6948 32916 -6916
rect 32936 -6924 32946 -6912
rect 32872 -6951 32880 -6950
rect 32902 -6951 32912 -6948
rect 32867 -6962 32912 -6951
rect 32790 -7138 32824 -6962
rect 32878 -7138 32912 -6962
rect 32902 -7150 32912 -7138
rect 32868 -7154 32912 -7150
rect 32868 -7188 32906 -7154
rect 32936 -7176 32950 -6924
rect 32936 -7188 32946 -7176
rect 32834 -7222 32906 -7188
rect 32958 -7256 32970 -6810
rect 32936 -7280 32970 -7256
rect 32958 -7284 32970 -7280
rect 32992 -7290 33026 -6810
rect 32274 -7324 32290 -7296
rect 31506 -7364 32238 -7330
rect 32246 -7330 32262 -7324
rect 32246 -7352 32266 -7330
rect 32258 -7364 32266 -7352
rect 31506 -7380 31540 -7364
rect 31506 -7391 31517 -7380
rect 31529 -7391 31540 -7380
rect 32204 -7380 32238 -7364
rect 32204 -7391 32215 -7380
rect 32227 -7391 32238 -7380
rect 32292 -7398 32300 -7296
rect 32676 -7324 33026 -7290
rect 33152 -6810 33502 -6776
rect 33152 -7290 33186 -6810
rect 33344 -6878 33382 -6840
rect 33310 -6912 33382 -6878
rect 33255 -6962 33300 -6951
rect 33343 -6962 33388 -6951
rect 33266 -7138 33300 -6962
rect 33354 -7138 33388 -6962
rect 33344 -7188 33382 -7150
rect 33310 -7222 33382 -7188
rect 33468 -7290 33502 -6810
rect 34252 -7280 34286 -4980
rect 34378 -5178 34384 -4812
rect 34490 -5592 34952 -4954
rect 34976 -5408 34978 -5364
rect 34544 -5676 34894 -5642
rect 34544 -6156 34578 -5676
rect 34736 -5710 34774 -5706
rect 34728 -5712 34786 -5710
rect 34736 -5744 34774 -5712
rect 34702 -5778 34774 -5744
rect 34647 -5828 34692 -5817
rect 34735 -5828 34780 -5817
rect 34658 -6004 34692 -5828
rect 34746 -6004 34780 -5828
rect 34736 -6054 34774 -6016
rect 34702 -6088 34774 -6054
rect 34860 -6150 34894 -5676
rect 34910 -6116 34928 -5712
rect 34948 -5726 34950 -5618
rect 34976 -5726 34978 -5618
rect 34860 -6156 34898 -6150
rect 34544 -6190 34898 -6156
rect 34876 -6368 34898 -6190
rect 34910 -6402 34932 -6116
rect 33152 -7324 33502 -7290
rect 32340 -7356 32908 -7330
rect 32340 -7364 32910 -7356
rect 32958 -7398 32974 -7324
rect 32986 -7370 33002 -7324
rect 35024 -7370 35058 2142
rect 35595 2106 39219 2142
rect 35631 -3470 35665 2106
rect 38377 877 38411 2106
rect 35733 843 39081 877
rect 35745 822 35779 843
rect 36403 822 36437 843
rect 37061 822 37095 843
rect 37719 822 37753 843
rect 38377 822 38411 843
rect 39035 822 39069 843
rect 35745 775 39069 822
rect 35745 707 35785 775
rect 35795 741 36443 775
rect 35795 735 35813 741
rect 36369 735 36387 741
rect 36397 707 36443 741
rect 36453 741 37101 775
rect 36453 735 36471 741
rect 37027 735 37045 741
rect 37055 707 37101 741
rect 37111 741 37759 775
rect 37111 735 37129 741
rect 37685 735 37703 741
rect 37713 707 37759 741
rect 37769 741 38417 775
rect 37769 735 37787 741
rect 38343 735 38361 741
rect 38371 707 38417 741
rect 38427 741 39069 775
rect 38427 735 38445 741
rect 39001 735 39019 741
rect 39029 707 39069 741
rect 35707 -3460 35708 -3378
rect 35745 -3470 35779 707
rect 35574 -3504 35868 -3470
rect 35631 -3572 35665 -3504
rect 35638 -3615 35665 -3572
rect 35733 -3606 35739 -3525
rect 35597 -3857 35626 -3649
rect 35631 -3891 35665 -3615
rect 35745 -3665 35779 -3504
rect 35720 -3841 35779 -3665
rect 35638 -3934 35665 -3891
rect 35726 -3924 35730 -3898
rect 35733 -3934 35739 -3853
rect 35631 -3968 35665 -3934
rect 35612 -3988 35712 -3968
rect 35631 -3996 35665 -3988
rect 35606 -4002 35712 -3996
rect 35745 -4002 35779 -3841
rect 35834 -4002 35868 -3504
rect 35574 -4036 35868 -4002
rect 35954 -3504 36344 -3470
rect 35954 -4002 35988 -3504
rect 36168 -3572 36215 -3525
rect 36130 -3606 36215 -3572
rect 36057 -3665 36102 -3654
rect 36185 -3665 36230 -3654
rect 36068 -3841 36102 -3665
rect 36196 -3841 36230 -3665
rect 36168 -3900 36215 -3853
rect 36130 -3934 36215 -3900
rect 36310 -4002 36344 -3504
rect 35954 -4036 36344 -4002
rect 35626 -4048 35665 -4036
rect 35631 -4086 35665 -4048
rect 35745 -4086 35779 -4036
rect 35595 -4652 35882 -4086
rect 35936 -4652 36358 -4086
rect 36403 -4652 36437 707
rect 36492 -4014 36502 -3664
rect 36520 -4014 36530 -3636
rect 36492 -4488 36502 -4200
rect 36520 -4516 36530 -4200
rect 37061 -4652 37095 707
rect 37719 -4652 37753 707
rect 38377 -4652 38411 707
rect 39035 -4652 39069 707
rect 35595 -4699 36358 -4652
rect 36375 -4665 36437 -4652
rect 37033 -4665 37095 -4652
rect 37691 -4665 37753 -4652
rect 38349 -4665 38411 -4652
rect 36375 -4693 36443 -4665
rect 37033 -4693 37101 -4665
rect 37691 -4693 37759 -4665
rect 38349 -4693 38417 -4665
rect 39007 -4693 39069 -4652
rect 36369 -4699 36443 -4693
rect 36453 -4699 36471 -4693
rect 37027 -4699 37101 -4693
rect 37111 -4699 37129 -4693
rect 37685 -4699 37759 -4693
rect 37769 -4699 37787 -4693
rect 38343 -4699 38417 -4693
rect 38427 -4699 38445 -4693
rect 39001 -4699 39069 -4693
rect 35595 -4706 36443 -4699
rect 35066 -6008 35074 -5906
rect 35094 -6032 35102 -5934
rect 35631 -6124 35665 -4706
rect 35707 -4788 35730 -4706
rect 35745 -4767 35794 -4706
rect 35795 -4733 36443 -4706
rect 36449 -4733 37101 -4699
rect 37107 -4733 37759 -4699
rect 37765 -4733 38417 -4699
rect 38423 -4733 39069 -4699
rect 35795 -4739 35822 -4733
rect 36369 -4739 36387 -4733
rect 36397 -4767 36443 -4733
rect 36453 -4739 36471 -4733
rect 37027 -4739 37045 -4733
rect 37055 -4767 37101 -4733
rect 37111 -4739 37129 -4733
rect 37685 -4739 37703 -4733
rect 37713 -4767 37759 -4733
rect 37769 -4739 37787 -4733
rect 38343 -4739 38361 -4733
rect 38371 -4767 38417 -4733
rect 38427 -4739 38445 -4733
rect 39001 -4739 39019 -4733
rect 39029 -4767 39069 -4733
rect 35745 -4801 35779 -4767
rect 36403 -4801 36437 -4767
rect 37061 -4801 37095 -4767
rect 37719 -4801 37753 -4767
rect 38377 -4801 38411 -4767
rect 39035 -4801 39069 -4767
rect 35727 -4835 39081 -4801
rect 39087 -4835 39103 -4801
rect 35707 -6114 35708 -6032
rect 35745 -6090 35746 -5994
rect 35745 -6124 35806 -6090
rect 35574 -6158 35868 -6124
rect 35631 -6226 35665 -6158
rect 35638 -6269 35665 -6226
rect 35733 -6260 35739 -6179
rect 35597 -6511 35626 -6303
rect 35631 -6545 35665 -6269
rect 35745 -6319 35779 -6158
rect 35720 -6495 35779 -6319
rect 35638 -6546 35665 -6545
rect 35612 -6564 35712 -6546
rect 35638 -6588 35665 -6564
rect 35726 -6578 35730 -6552
rect 35733 -6588 35739 -6507
rect 35631 -6622 35665 -6588
rect 35745 -6622 35779 -6495
rect 35612 -6642 35712 -6622
rect 35631 -6650 35665 -6642
rect 35606 -6656 35712 -6650
rect 35745 -6656 35806 -6622
rect 35834 -6656 35868 -6158
rect 35574 -6690 35868 -6656
rect 35954 -6158 36344 -6124
rect 35954 -6656 35988 -6158
rect 36168 -6226 36215 -6179
rect 36130 -6260 36215 -6226
rect 36057 -6319 36102 -6308
rect 36185 -6319 36230 -6308
rect 36068 -6495 36102 -6319
rect 36196 -6495 36230 -6319
rect 36168 -6554 36215 -6507
rect 36130 -6588 36215 -6554
rect 36310 -6656 36344 -6158
rect 35954 -6690 36344 -6656
rect 36492 -6668 36502 -6368
rect 36520 -6554 36558 -6368
rect 36520 -6668 36530 -6554
rect 35626 -6702 35665 -6690
rect 35631 -6740 35665 -6702
rect 35595 -7360 35882 -6740
rect 35936 -7360 36358 -6740
rect 36492 -7142 36502 -6854
rect 36520 -7170 36530 -6854
rect 35767 -7421 35794 -7360
rect 35795 -7393 35822 -7360
rect 39149 -7393 39183 2106
rect 40702 -7370 40736 2142
rect 42866 1664 42886 1860
rect 43448 882 43482 2142
rect 40804 848 44152 882
rect 40816 818 40850 848
rect 41474 818 41508 848
rect 42132 818 42166 848
rect 42790 818 42824 848
rect 43448 818 43482 848
rect 44106 818 44140 848
rect 40816 780 44140 818
rect 40816 -4642 40850 780
rect 40878 746 41514 780
rect 41440 740 41458 746
rect 41468 712 41514 746
rect 41524 746 42172 780
rect 41524 740 41542 746
rect 42098 740 42116 746
rect 42126 712 42172 746
rect 42182 746 42830 780
rect 42182 740 42200 746
rect 42756 740 42774 746
rect 42784 712 42830 746
rect 42840 746 43488 780
rect 42840 740 42858 746
rect 43414 740 43432 746
rect 43442 712 43488 746
rect 43498 746 44140 780
rect 43498 740 43516 746
rect 44072 740 44090 746
rect 44100 712 44140 746
rect 40882 -3476 40888 -3220
rect 40910 -3448 40916 -3248
rect 40882 -3876 40888 -3620
rect 40910 -3848 40916 -3648
rect 41474 -4638 41508 712
rect 42132 -4638 42166 712
rect 42790 -4638 42824 712
rect 43448 -4638 43482 712
rect 44106 -4638 44140 712
rect 41446 -4642 41508 -4638
rect 42104 -4642 42166 -4638
rect 42762 -4642 42824 -4638
rect 43420 -4642 43482 -4638
rect 40816 -4744 40856 -4642
rect 41446 -4670 41514 -4642
rect 42104 -4670 42172 -4642
rect 42762 -4670 42830 -4642
rect 43420 -4670 43488 -4642
rect 44078 -4670 44140 -4638
rect 40866 -4676 40884 -4670
rect 41440 -4676 41514 -4670
rect 41524 -4676 41542 -4670
rect 42098 -4676 42172 -4670
rect 42182 -4676 42200 -4670
rect 42756 -4676 42830 -4670
rect 42840 -4676 42858 -4670
rect 43414 -4676 43488 -4670
rect 43498 -4676 43516 -4670
rect 44072 -4676 44140 -4670
rect 40862 -4710 41514 -4676
rect 41520 -4710 42172 -4676
rect 42178 -4710 42830 -4676
rect 42836 -4710 43488 -4676
rect 43494 -4710 44140 -4676
rect 40866 -4716 40884 -4710
rect 41440 -4716 41458 -4710
rect 41468 -4744 41514 -4710
rect 41524 -4716 41542 -4710
rect 42098 -4716 42116 -4710
rect 42126 -4744 42172 -4710
rect 42182 -4716 42200 -4710
rect 42756 -4716 42774 -4710
rect 42784 -4744 42830 -4710
rect 42840 -4716 42858 -4710
rect 43414 -4716 43432 -4710
rect 43442 -4744 43488 -4710
rect 43498 -4716 43516 -4710
rect 44072 -4716 44090 -4710
rect 44100 -4744 44140 -4710
rect 40816 -4778 40850 -4744
rect 41474 -4778 41508 -4744
rect 42132 -4778 42166 -4744
rect 42790 -4778 42824 -4744
rect 43448 -4778 43482 -4744
rect 44106 -4778 44140 -4744
rect 40798 -4812 44174 -4778
rect 41474 -7280 41508 -4812
rect 44220 -7370 44254 2142
rect 49885 2106 53509 2142
rect 58029 2120 58580 2156
rect 58772 2167 60254 2235
rect 60545 2167 60579 2235
rect 60811 2167 60856 2235
rect 61102 2219 61160 2235
rect 61114 2167 61148 2219
rect 61228 2167 61262 2235
rect 61457 2229 61515 2235
rect 61370 2206 61406 2229
rect 61426 2219 61515 2229
rect 61370 2167 61386 2206
rect 61426 2167 61462 2219
rect 61500 2204 61515 2219
rect 61469 2167 61503 2201
rect 61583 2167 61617 2235
rect 62040 2222 62068 2229
rect 62096 2222 62124 2229
rect 62502 2208 64133 2235
rect 64566 2224 64604 2246
rect 64554 2208 64612 2224
rect 65140 2208 65174 2276
rect 65316 2258 68992 2276
rect 69054 2262 69516 2882
rect 69570 2262 69992 2882
rect 70046 2269 70468 2882
rect 70989 2760 71023 2960
rect 70955 2316 70978 2760
rect 70983 2316 71029 2760
rect 71262 2316 71296 3287
rect 70955 2288 71008 2316
rect 70961 2269 71008 2288
rect 71250 2269 71308 2316
rect 70046 2262 71008 2269
rect 65320 2252 65356 2258
rect 65224 2224 65262 2246
rect 65616 2224 65650 2258
rect 65804 2252 66008 2258
rect 66456 2252 66492 2258
rect 65804 2246 65834 2252
rect 65862 2246 66008 2252
rect 65870 2242 65928 2246
rect 66528 2242 67740 2258
rect 67824 2252 67858 2258
rect 65882 2224 65920 2242
rect 66540 2224 66586 2242
rect 66654 2224 66688 2242
rect 67360 2234 67722 2242
rect 67780 2240 67808 2252
rect 67824 2246 67864 2252
rect 67824 2242 67858 2246
rect 67824 2231 67835 2242
rect 67847 2231 67858 2242
rect 68488 2240 68516 2252
rect 68658 2242 68692 2258
rect 68658 2231 68669 2242
rect 68681 2231 68692 2242
rect 65212 2214 67682 2224
rect 65212 2208 67694 2214
rect 62502 2190 66586 2208
rect 66654 2190 66688 2208
rect 67116 2206 67694 2208
rect 67116 2190 67360 2206
rect 67824 2190 67858 2214
rect 69054 2190 69222 2262
rect 62502 2174 69222 2190
rect 62502 2167 64133 2174
rect 58772 2133 64133 2167
rect 64554 2136 64612 2174
rect 65140 2156 69222 2174
rect 70217 2167 70251 2262
rect 70393 2235 71008 2262
rect 71051 2235 71308 2269
rect 71250 2219 71308 2235
rect 71293 2204 71308 2219
rect 71262 2167 71296 2201
rect 71376 2167 71410 3448
rect 72951 2346 73009 2364
rect 73037 2346 73071 10363
rect 73140 10304 73196 10315
rect 73610 10304 73666 10315
rect 73151 6816 73196 10304
rect 73621 6816 73666 10304
rect 73735 10010 73769 10363
rect 75147 10329 75174 10431
rect 75175 10357 75202 10403
rect 73735 8658 73772 10010
rect 73151 4422 73185 6816
rect 73370 6498 73582 6506
rect 73214 6058 73582 6498
rect 73214 6050 73426 6058
rect 73621 4422 73655 6816
rect 73151 3418 73196 4422
rect 73621 3418 73666 4422
rect 73151 2346 73185 3418
rect 73621 2346 73655 3418
rect 73735 2346 73769 8658
rect 73809 2364 73843 10304
rect 75202 9232 75204 10016
rect 75252 9232 76625 10465
rect 76688 10433 76726 10440
rect 76676 10368 76726 10433
rect 77146 10433 77184 10440
rect 77146 10418 77192 10433
rect 77134 10402 77192 10418
rect 76780 10368 77192 10402
rect 76676 10330 76722 10368
rect 77134 10330 77192 10368
rect 73944 9198 76625 9232
rect 73870 8658 73894 8856
rect 73870 7932 73876 8180
rect 73944 6946 73978 9198
rect 74467 9118 74501 9198
rect 75125 9118 75159 9198
rect 75202 9124 75204 9198
rect 75252 9118 76625 9198
rect 73999 9056 74080 9103
rect 74139 9084 76625 9118
rect 74454 9072 74455 9073
rect 74455 9071 74456 9072
rect 74046 7088 74080 9056
rect 74467 7164 74501 9084
rect 74513 9072 74514 9073
rect 75112 9072 75113 9073
rect 74512 9071 74513 9072
rect 75113 9071 75114 9072
rect 75125 7164 75159 9084
rect 75171 9072 75172 9073
rect 75170 9071 75171 9072
rect 75202 8800 75204 9078
rect 74467 7073 74512 7164
rect 75125 7073 75170 7164
rect 74455 7072 74456 7073
rect 74467 7072 74513 7073
rect 75113 7072 75114 7073
rect 75125 7072 75171 7073
rect 74454 7071 74455 7072
rect 74448 7060 74455 7071
rect 74467 7060 74501 7072
rect 74513 7071 74514 7072
rect 75112 7071 75113 7072
rect 74513 7060 75113 7071
rect 75125 7060 75159 7072
rect 75171 7071 75172 7072
rect 75202 7071 75220 7164
rect 75171 7060 75220 7071
rect 75252 7060 76625 9084
rect 76682 10318 76722 10330
rect 76734 10318 76752 10329
rect 76682 7738 76752 10318
rect 76666 7670 76752 7738
rect 76666 7464 76763 7670
rect 77146 7618 77180 10330
rect 77260 9470 77294 10470
rect 78108 10402 78142 10449
rect 78806 10418 78817 10429
rect 78829 10418 78840 10429
rect 78806 10402 78840 10418
rect 78108 10368 78840 10402
rect 77260 9360 77428 9470
rect 77260 9334 77444 9360
rect 77260 7618 77294 9334
rect 77352 8902 77444 9334
rect 78108 9326 78142 10368
rect 78211 10318 78256 10329
rect 78681 10318 78726 10329
rect 78222 9770 78256 10318
rect 78692 9770 78726 10318
rect 78222 9326 78267 9770
rect 78692 9348 78737 9770
rect 78806 9754 78840 10368
rect 79368 10054 79402 10470
rect 79510 10446 79576 10466
rect 79496 10436 79576 10446
rect 79496 10428 79602 10436
rect 79496 10424 79580 10428
rect 79496 10418 79510 10424
rect 79542 10418 79576 10424
rect 79584 10416 79618 10418
rect 79448 10408 79510 10416
rect 79448 10402 79522 10408
rect 79468 10400 79526 10402
rect 79476 10398 79526 10400
rect 79476 10396 79522 10398
rect 79488 10394 79516 10396
rect 79528 10394 79558 10416
rect 79584 10402 79638 10416
rect 79570 10400 79630 10402
rect 79570 10394 79600 10400
rect 79470 10382 79548 10394
rect 79569 10382 79616 10394
rect 79470 10368 79544 10382
rect 79470 10330 79526 10368
rect 79538 10330 79550 10334
rect 79570 10330 79616 10382
rect 79482 10206 79522 10330
rect 79448 10166 79454 10196
rect 79476 10194 79482 10196
rect 79504 10194 79522 10206
rect 79528 10318 79558 10330
rect 79570 10318 79604 10330
rect 79528 10206 79604 10318
rect 79528 10194 79572 10206
rect 79504 10190 79516 10194
rect 79528 10190 79576 10194
rect 79528 10172 79594 10190
rect 79526 10122 79594 10172
rect 79526 10106 79576 10122
rect 79684 10054 79718 10470
rect 80848 10318 80894 10330
rect 80854 10306 80894 10318
rect 79368 10020 79718 10054
rect 78668 9326 78760 9348
rect 78806 9326 78858 9754
rect 77872 8388 80838 9326
rect 81384 9294 81696 9330
rect 82233 9294 82267 10403
rect 82472 10068 85821 10535
rect 87452 10504 89102 11482
rect 89538 10504 90892 11482
rect 93732 11344 93750 11566
rect 93760 11543 93824 11566
rect 93766 11540 93824 11543
rect 95050 11543 95122 11564
rect 95050 11540 95116 11543
rect 95050 11368 95072 11540
rect 87304 10470 90892 10504
rect 87304 10144 87338 10470
rect 87452 10402 89102 10470
rect 89364 10402 89402 10440
rect 89538 10402 90892 10470
rect 87452 10368 89402 10402
rect 89454 10368 90892 10402
rect 87452 10336 89102 10368
rect 89538 10334 90892 10368
rect 90681 10330 90682 10331
rect 90754 10330 90776 10334
rect 90682 10329 90683 10330
rect 87407 10318 87452 10329
rect 88065 10318 88110 10329
rect 88723 10318 88768 10329
rect 89381 10318 89426 10329
rect 90039 10318 90084 10329
rect 87418 10144 87452 10318
rect 87463 10156 87464 10157
rect 88064 10156 88065 10157
rect 87464 10155 87465 10156
rect 88063 10155 88064 10156
rect 88076 10144 88110 10318
rect 88121 10156 88122 10157
rect 88722 10156 88723 10157
rect 88122 10155 88123 10156
rect 88721 10155 88722 10156
rect 88734 10144 88768 10318
rect 88779 10156 88780 10157
rect 89380 10156 89381 10157
rect 88780 10155 88781 10156
rect 89379 10155 89380 10156
rect 89392 10144 89426 10318
rect 89437 10156 89438 10157
rect 90038 10156 90039 10157
rect 89438 10155 89439 10156
rect 90037 10155 90038 10156
rect 90050 10144 90084 10318
rect 90696 10172 90776 10330
rect 90095 10156 90096 10157
rect 90696 10156 90754 10172
rect 90096 10155 90097 10156
rect 90670 10150 90681 10155
rect 90670 10144 90682 10150
rect 87270 10116 90686 10144
rect 90702 10120 90720 10156
rect 90739 10141 90754 10156
rect 90702 10116 90754 10120
rect 87270 10110 90754 10116
rect 87304 10068 87338 10110
rect 87418 10068 87452 10110
rect 87464 10098 87465 10099
rect 88063 10098 88064 10099
rect 87463 10097 87464 10098
rect 88064 10097 88065 10098
rect 82472 9497 87804 10068
rect 88076 9770 88110 10110
rect 88122 10098 88123 10099
rect 88721 10098 88722 10099
rect 88121 10097 88122 10098
rect 88722 10097 88723 10098
rect 88734 9770 88768 10110
rect 88780 10098 88781 10099
rect 89379 10098 89380 10099
rect 88779 10097 88780 10098
rect 89380 10097 89381 10098
rect 87998 9564 88032 9570
rect 88032 9514 88054 9564
rect 88076 9499 88121 9770
rect 88168 9564 88250 9570
rect 88064 9498 88065 9499
rect 88076 9498 88122 9499
rect 88063 9497 88064 9498
rect 82472 9496 88064 9497
rect 88076 9496 88110 9498
rect 88122 9497 88123 9498
rect 88174 9497 88194 9514
rect 88202 9497 88250 9564
rect 88734 9499 88779 9770
rect 88722 9498 88723 9499
rect 88734 9498 88780 9499
rect 89380 9498 89381 9499
rect 88721 9497 88722 9498
rect 88122 9496 88722 9497
rect 82472 9486 88722 9496
rect 88734 9486 88768 9498
rect 88780 9497 88781 9498
rect 89379 9497 89380 9498
rect 88780 9486 89358 9497
rect 89392 9486 89426 10110
rect 89438 10098 89439 10099
rect 90037 10098 90038 10099
rect 89437 10097 89438 10098
rect 90038 10097 90039 10098
rect 89437 9498 89438 9499
rect 90038 9498 90039 9499
rect 89438 9497 89439 9498
rect 90037 9497 90038 9498
rect 90050 9486 90084 10110
rect 90674 10104 90682 10110
rect 90096 10098 90097 10099
rect 90095 10097 90096 10098
rect 90686 10082 90754 10110
rect 90696 9514 90776 10082
rect 90095 9498 90096 9499
rect 90696 9498 90754 9514
rect 90096 9497 90097 9498
rect 90670 9486 90681 9497
rect 82472 9458 90686 9486
rect 90708 9462 90720 9498
rect 90739 9483 90754 9498
rect 90704 9458 90754 9462
rect 82472 9452 90754 9458
rect 82472 9330 87804 9452
rect 88006 9446 88174 9452
rect 88006 9360 88194 9446
rect 88202 9360 88250 9446
rect 88721 9440 88722 9441
rect 88734 9440 88768 9452
rect 88780 9440 88781 9441
rect 89379 9440 89380 9441
rect 88722 9439 88723 9440
rect 88734 9439 88780 9440
rect 89380 9439 89381 9440
rect 88006 9330 88174 9360
rect 88734 9330 88779 9439
rect 82347 9294 82381 9328
rect 82472 9294 89198 9330
rect 81384 9260 89198 9294
rect 78108 7618 78142 8388
rect 78222 7618 78256 8388
rect 78692 7618 78726 8388
rect 78806 7618 78840 8388
rect 80862 7624 80894 9062
rect 80918 7624 80922 9006
rect 81384 7962 81696 9260
rect 82233 9192 82267 9260
rect 82472 9239 89198 9260
rect 82136 8810 82146 9134
rect 82233 9133 82234 9165
rect 82238 9133 82267 9192
rect 82186 9106 82232 9111
rect 82233 9106 82267 9133
rect 82335 9158 89198 9239
rect 82335 9111 82393 9158
rect 82164 9099 82267 9106
rect 82164 9096 82226 9099
rect 82164 8838 82202 9096
rect 82186 8666 82202 8838
rect 82228 8838 82267 9099
rect 82186 8123 82226 8666
rect 82228 8123 82232 8838
rect 82186 8111 82232 8123
rect 82199 8107 82226 8111
rect 82233 8073 82267 8838
rect 82347 8666 82392 9111
rect 82472 8828 89198 9158
rect 89308 8912 89352 8932
rect 89352 8876 89364 8912
rect 89380 8840 89381 8841
rect 89379 8839 89380 8840
rect 89392 8828 89426 9452
rect 89438 9440 89439 9441
rect 90037 9440 90038 9441
rect 89437 9439 89438 9440
rect 90038 9439 90039 9440
rect 89437 8840 89438 8841
rect 90038 8840 90039 8841
rect 89438 8839 89439 8840
rect 90037 8839 90038 8840
rect 90050 8828 90084 9452
rect 90096 9440 90097 9441
rect 90095 9439 90096 9440
rect 90686 9424 90754 9452
rect 90696 8856 90776 9424
rect 90095 8840 90096 8841
rect 90696 8840 90754 8856
rect 90096 8839 90097 8840
rect 90670 8828 90681 8839
rect 82472 8794 90686 8828
rect 82472 8714 89198 8794
rect 89352 8714 89364 8740
rect 89392 8714 89426 8794
rect 90050 8714 90084 8794
rect 90708 8760 90720 8840
rect 90739 8825 90754 8840
rect 82472 8680 90754 8714
rect 82347 8111 82381 8666
rect 82472 8644 89198 8680
rect 82850 8606 82895 8644
rect 82850 8278 82884 8606
rect 82964 8476 82998 8644
rect 83005 8476 83045 8644
rect 83050 8630 83118 8644
rect 83050 8476 83101 8630
rect 83506 8476 83540 8644
rect 83620 8476 83654 8644
rect 83663 8476 83697 8644
rect 83818 8626 84040 8644
rect 84216 8608 84232 8644
rect 84278 8476 84312 8644
rect 84321 8476 84361 8644
rect 84372 8476 84389 8644
rect 84930 8608 84970 8644
rect 84936 8476 84970 8608
rect 84979 8476 85008 8644
rect 85050 8476 85084 8644
rect 85610 8484 85678 8644
rect 85712 8484 85737 8644
rect 85751 8484 85785 8644
rect 87268 8492 89198 8644
rect 89352 8632 89364 8680
rect 82942 8278 83934 8476
rect 82614 8111 83934 8278
rect 82238 8064 82267 8073
rect 82335 8064 82394 8111
rect 82472 8109 83934 8111
rect 82472 8064 84040 8109
rect 82238 8062 84040 8064
rect 84132 8062 85124 8476
rect 82238 8030 85124 8062
rect 82233 7962 82267 8030
rect 82335 8014 82393 8030
rect 82614 8028 85124 8030
rect 82335 7999 82350 8014
rect 82347 7962 82381 7996
rect 82614 7962 83948 8028
rect 81384 7960 83948 7962
rect 83970 7960 84008 8020
rect 84062 7972 84086 8018
rect 84076 7960 84086 7972
rect 84132 7960 85124 8028
rect 81384 7928 85124 7960
rect 81384 7892 81696 7928
rect 76688 7446 76763 7464
rect 76662 7218 76808 7446
rect 76688 7208 76763 7218
rect 76628 7178 76634 7208
rect 76656 7206 76763 7208
rect 76790 7206 76814 7208
rect 76666 7148 76763 7206
rect 76818 7178 76842 7208
rect 74139 7026 76625 7060
rect 76654 7034 76660 7076
rect 76682 7074 76763 7148
rect 76682 7062 76688 7074
rect 76718 7062 76763 7074
rect 76850 7062 79158 7618
rect 74467 6974 74501 7026
rect 74446 6946 74836 6974
rect 75125 6946 75159 7026
rect 75202 6946 75220 7020
rect 75252 6946 76625 7026
rect 76714 7024 79158 7062
rect 76718 6990 79158 7024
rect 76718 6974 76764 6990
rect 73944 6922 76625 6946
rect 76850 6922 79158 6990
rect 73944 6912 79158 6922
rect 74446 6442 74480 6912
rect 74660 6872 74707 6912
rect 74622 6838 74707 6872
rect 74549 6779 74594 6790
rect 74677 6779 74722 6790
rect 74560 6603 74594 6779
rect 74688 6603 74722 6779
rect 74660 6544 74707 6591
rect 74622 6510 74707 6544
rect 74680 6506 74686 6510
rect 74692 6470 74698 6506
rect 74802 6442 74836 6912
rect 75008 6754 75016 6784
rect 74980 6726 75016 6728
rect 74446 6408 74836 6442
rect 74432 5738 74854 6358
rect 75125 5742 75159 6912
rect 75202 6590 75220 6912
rect 75252 6888 79158 6912
rect 75230 6754 75246 6784
rect 75252 6728 76625 6888
rect 76712 6820 76716 6876
rect 75230 6726 76625 6728
rect 75202 6582 75218 6590
rect 75252 6464 76625 6726
rect 75252 6208 76634 6464
rect 76648 6236 76690 6436
rect 75060 5656 75159 5742
rect 75010 4792 75036 5596
rect 75038 4792 75064 5596
rect 75125 4792 75159 5656
rect 75202 5596 75204 6144
rect 75252 4792 76625 6208
rect 76850 6180 79158 6888
rect 79428 7554 81696 7624
rect 79428 6256 81700 7554
rect 79428 6186 81696 6256
rect 76960 6030 77172 6180
rect 77288 5996 77322 6180
rect 77346 5996 77356 6180
rect 77376 6150 77416 6180
rect 77426 6178 77444 6180
rect 77480 6178 77502 6180
rect 77508 6150 77530 6180
rect 77376 6136 77410 6150
rect 77422 6136 77447 6147
rect 77479 6136 77535 6147
rect 77376 5996 77447 6136
rect 77490 5996 77535 6136
rect 77604 6024 77840 6180
rect 77604 5996 77638 6024
rect 74452 4766 76625 4792
rect 74446 3368 74520 3698
rect 74446 3214 74652 3368
rect 74446 3044 74520 3214
rect 73797 2346 73855 2364
rect 74455 2346 74513 2364
rect 75010 2346 75036 4766
rect 75038 2346 75064 4766
rect 75125 2364 75159 4766
rect 75113 2346 75171 2364
rect 75252 2346 76625 4766
rect 76910 5962 77830 5996
rect 76910 4682 76944 5962
rect 77288 5894 77322 5962
rect 77346 5932 77356 5962
rect 77376 5960 77447 5962
rect 77490 5960 77535 5962
rect 77376 5948 77410 5960
rect 77416 5948 77430 5956
rect 77496 5948 77508 5956
rect 77376 5946 77518 5948
rect 77376 5932 77524 5946
rect 77604 5932 77638 5962
rect 77346 5894 77692 5932
rect 77086 5860 77692 5894
rect 77013 5810 77058 5821
rect 77024 4834 77058 5810
rect 77288 5808 77322 5860
rect 77346 5842 77356 5860
rect 77364 5842 77422 5860
rect 77346 5822 77422 5842
rect 77346 5814 77421 5822
rect 77350 5808 77421 5814
rect 77604 5808 77638 5860
rect 77671 5810 77727 5821
rect 77288 5774 77638 5808
rect 77376 4822 77421 5774
rect 77682 4834 77727 5810
rect 77346 4784 77692 4822
rect 77086 4750 77692 4784
rect 77364 4734 77422 4750
rect 77376 4682 77410 4734
rect 77796 4682 77830 5962
rect 78000 5596 78024 6144
rect 77912 5468 77922 5574
rect 78008 5470 78018 5574
rect 78028 4744 78052 6172
rect 78108 5996 78142 6180
rect 78222 5996 78267 6180
rect 78272 6030 78678 6180
rect 78272 6012 78484 6030
rect 78692 5996 78726 6180
rect 78806 5996 78840 6180
rect 82233 6052 82267 7928
rect 82614 7926 85124 7928
rect 82614 7856 83948 7926
rect 82942 7802 83948 7856
rect 82614 7448 83948 7802
rect 83970 7508 84008 7926
rect 84076 7914 84086 7926
rect 82614 7380 83934 7448
rect 82942 7056 83934 7380
rect 84132 7056 85124 7926
rect 82351 6052 82381 7039
rect 85442 7005 86434 8484
rect 86610 8460 89198 8492
rect 89392 8460 89426 8494
rect 90050 8460 90084 8494
rect 90708 8460 90742 8494
rect 90822 8460 90856 10334
rect 93768 8576 93806 11344
rect 93824 8632 93834 11344
rect 95321 8693 95520 12028
rect 100471 11509 100505 12133
rect 100557 12121 101202 12133
rect 100573 12050 101202 12121
rect 101252 12127 101308 12133
rect 101252 12098 101286 12127
rect 101784 12098 101818 12133
rect 103540 12105 103621 12139
rect 101252 12064 101818 12098
rect 100573 11577 100607 12050
rect 100950 11602 101080 11618
rect 101280 11602 102408 11618
rect 100978 11574 101080 11590
rect 101280 11574 102380 11590
rect 101802 11555 102380 11574
rect 103587 11561 103621 12105
rect 101802 11549 103266 11555
rect 103540 11549 103637 11561
rect 103689 11549 103723 12247
rect 100666 11543 108642 11549
rect 100437 11475 100505 11509
rect 100526 11521 100607 11522
rect 100526 11509 100641 11521
rect 100650 11515 108642 11543
rect 100526 11503 100607 11509
rect 100616 11503 103544 11509
rect 100526 11494 103544 11503
rect 100526 11481 103621 11494
rect 100526 11475 103539 11481
rect 100471 10851 100505 11475
rect 100557 11463 100654 11475
rect 100573 10919 100607 11463
rect 101080 11446 101280 11456
rect 103540 11447 103621 11481
rect 101052 11418 101308 11428
rect 103587 10903 103621 11447
rect 103540 10891 103637 10903
rect 100666 10885 103637 10891
rect 100437 10817 100505 10851
rect 100526 10863 100607 10864
rect 100650 10863 103637 10885
rect 100526 10851 100641 10863
rect 100650 10857 103578 10863
rect 100526 10845 100607 10851
rect 100616 10845 103544 10851
rect 100526 10836 103544 10845
rect 100526 10823 103621 10836
rect 100526 10817 103539 10823
rect 100471 10193 100505 10817
rect 100557 10805 100654 10817
rect 100573 10261 100607 10805
rect 103540 10789 103621 10823
rect 101888 10768 103240 10786
rect 101860 10740 103268 10758
rect 100928 10280 102386 10298
rect 100956 10252 102358 10270
rect 103587 10245 103621 10789
rect 103540 10233 103637 10245
rect 100666 10227 103637 10233
rect 100437 10159 100505 10193
rect 100526 10205 100607 10206
rect 100650 10205 103637 10227
rect 100526 10193 100641 10205
rect 100650 10199 103578 10205
rect 100526 10187 100607 10193
rect 100616 10187 103544 10193
rect 100526 10178 103544 10187
rect 100526 10165 103621 10178
rect 100526 10159 103539 10165
rect 100471 9461 100505 10159
rect 100557 10147 100654 10159
rect 100573 9603 100607 10147
rect 103540 10131 103621 10165
rect 103587 9587 103621 10131
rect 103540 9575 103637 9587
rect 100666 9569 103637 9575
rect 100650 9547 103637 9569
rect 100650 9541 103578 9547
rect 100616 9507 103544 9535
rect 100628 9503 103528 9507
rect 103587 9473 103621 9495
rect 103689 9461 103723 11515
rect 163952 10499 163986 11642
rect 165511 10499 165545 12203
rect 165987 12197 166021 12235
rect 169029 12213 169040 12224
rect 169052 12213 169063 12224
rect 169029 12197 169063 12213
rect 165687 12163 169363 12197
rect 165987 10499 166021 12163
rect 166090 12104 166146 12115
rect 166272 12104 166328 12115
rect 166748 12104 166804 12115
rect 166930 12104 166986 12115
rect 167406 12104 167451 12115
rect 167588 12104 167633 12115
rect 168064 12104 168109 12115
rect 168246 12104 168291 12115
rect 168722 12104 168767 12115
rect 168904 12104 168949 12115
rect 166101 11848 166822 12104
rect 166101 10499 166146 11848
rect 166162 10499 166190 11780
rect 166283 10499 166328 11848
rect 166759 10499 166804 11848
rect 166820 10499 166848 11780
rect 166876 10499 166904 11780
rect 166941 10499 166986 12104
rect 163643 10465 167195 10499
rect 108667 9553 108674 9626
rect 108701 9587 108708 9660
rect 100471 9427 108741 9461
rect 103689 8825 103723 9427
rect 151710 9198 151744 9930
rect 152482 9292 152516 9326
rect 153140 9292 153174 9326
rect 154312 9294 154322 9348
rect 154428 9294 154436 9328
rect 155060 9294 155094 9328
rect 155718 9294 155752 9328
rect 156376 9294 156410 9328
rect 156490 9294 156524 9936
rect 152262 9258 153840 9292
rect 151710 8756 151754 9198
rect 103104 8732 103362 8744
rect 151720 8476 151754 8756
rect 152262 8694 152296 9258
rect 152398 9122 152422 9224
rect 152482 9206 152529 9237
rect 152426 9190 152450 9196
rect 152470 9190 152529 9206
rect 153006 9190 153053 9237
rect 152426 9156 153053 9190
rect 152426 9150 152450 9156
rect 152470 9109 152528 9156
rect 153056 9122 153074 9224
rect 153140 9206 153187 9237
rect 153084 9190 153102 9196
rect 153128 9190 153187 9206
rect 153664 9190 153711 9237
rect 153806 9230 153840 9258
rect 153772 9196 153840 9230
rect 154366 9238 154376 9294
rect 154390 9260 157822 9294
rect 154390 9238 154400 9260
rect 153084 9156 153711 9190
rect 153084 9154 153102 9156
rect 153128 9154 153186 9156
rect 153084 9150 153186 9154
rect 153128 9126 153186 9150
rect 153104 9122 153186 9126
rect 152365 9097 152410 9108
rect 152376 8843 152410 9097
rect 152482 8855 152516 9109
rect 153023 9097 153068 9108
rect 153034 8843 153068 9097
rect 153076 8928 153098 9104
rect 153104 8900 153126 9122
rect 153128 9109 153186 9122
rect 153140 8855 153174 9109
rect 153681 9097 153726 9108
rect 153692 8843 153726 9097
rect 153806 8889 153866 9196
rect 153798 8855 153866 8889
rect 152364 8796 152423 8843
rect 152454 8802 152501 8843
rect 152446 8796 152501 8802
rect 153022 8796 153081 8843
rect 153112 8802 153159 8843
rect 153100 8796 153159 8802
rect 153680 8796 153738 8843
rect 152364 8762 152501 8796
rect 152544 8762 153159 8796
rect 153202 8762 153738 8796
rect 153772 8762 153786 8796
rect 152364 8746 152422 8762
rect 152446 8756 152466 8762
rect 152364 8731 152379 8746
rect 152474 8728 152494 8762
rect 153022 8746 153080 8762
rect 153100 8756 153124 8762
rect 153128 8728 153152 8762
rect 153680 8746 153738 8762
rect 153723 8731 153738 8746
rect 153806 8694 153840 8855
rect 154366 8700 154400 9238
rect 154402 8845 154434 9238
rect 155060 9208 155107 9239
rect 155048 9192 155107 9208
rect 155110 9192 155157 9239
rect 155718 9208 155765 9239
rect 155706 9192 155765 9208
rect 155768 9192 155815 9239
rect 156376 9208 156422 9239
rect 156364 9192 156422 9208
rect 156490 9192 156524 9260
rect 154542 9158 155157 9192
rect 155200 9158 155815 9192
rect 155858 9158 156422 9192
rect 156426 9158 156444 9192
rect 154446 9110 154470 9139
rect 155048 9111 155106 9158
rect 155706 9152 155780 9158
rect 155706 9132 155764 9152
rect 155706 9124 155790 9132
rect 155706 9111 155764 9124
rect 156364 9122 156422 9158
rect 156490 9133 156496 9165
rect 156500 9133 156524 9192
rect 156364 9111 156444 9122
rect 154474 9110 154498 9111
rect 154446 9099 154514 9110
rect 154446 8856 154470 9099
rect 154474 8849 154514 9099
rect 155060 8892 155100 9111
rect 155127 9106 155172 9110
rect 155110 9099 155172 9106
rect 155110 8920 155128 9099
rect 155060 8861 155094 8892
rect 155138 8849 155172 9099
rect 155718 8861 155752 9111
rect 155785 9099 155830 9110
rect 155796 8849 155830 9099
rect 156376 8872 156416 9111
rect 156420 8900 156444 9111
rect 156376 8861 156410 8872
rect 154468 8802 154527 8849
rect 155032 8802 155079 8849
rect 155126 8802 155185 8849
rect 155690 8802 155737 8849
rect 155784 8802 155843 8849
rect 156348 8802 156395 8849
rect 154468 8768 155079 8802
rect 155122 8768 155737 8802
rect 155780 8768 156395 8802
rect 154468 8752 154526 8768
rect 155126 8752 155184 8768
rect 155784 8752 155842 8768
rect 154468 8737 154483 8752
rect 156454 8700 156462 8734
rect 156490 8700 156524 9133
rect 151806 8660 153850 8694
rect 154366 8666 156524 8700
rect 152262 8556 152296 8660
rect 152156 8536 152818 8556
rect 152198 8516 152764 8536
rect 152262 8512 152296 8516
rect 152226 8488 152764 8512
rect 152262 8476 152296 8488
rect 153806 8476 153840 8660
rect 154366 8484 154400 8666
rect 86610 8426 91262 8460
rect 86610 8358 89198 8426
rect 89208 8358 89246 8396
rect 89392 8374 89430 8396
rect 89380 8358 89438 8374
rect 89866 8358 89904 8396
rect 90050 8374 90088 8396
rect 90038 8358 90096 8374
rect 90524 8358 90562 8396
rect 90708 8389 90746 8396
rect 90708 8374 90754 8389
rect 90696 8358 90754 8374
rect 86610 8324 89246 8358
rect 89298 8324 89904 8358
rect 89956 8324 90562 8358
rect 90614 8324 90754 8358
rect 86610 7041 89198 8324
rect 89225 8274 89270 8285
rect 89236 7041 89270 8274
rect 89274 7041 89308 8318
rect 89330 7041 89364 8318
rect 89380 8286 89438 8324
rect 89392 7041 89426 8286
rect 89883 8274 89928 8285
rect 89894 7041 89928 8274
rect 89932 7041 89972 8318
rect 89988 7041 90028 8318
rect 90038 8286 90096 8324
rect 90050 7041 90084 8286
rect 90541 8274 90586 8285
rect 90552 7041 90586 8274
rect 90652 7041 90680 8318
rect 90696 8286 90754 8324
rect 90708 7041 90742 8286
rect 86610 7005 90787 7041
rect 82385 6971 90787 7005
rect 82385 6052 82419 6971
rect 82936 6891 82993 6902
rect 83005 6891 83039 6971
rect 83629 6924 83634 6926
rect 83657 6924 83662 6954
rect 83051 6896 83651 6902
rect 83663 6896 83697 6971
rect 84321 6952 84361 6971
rect 84287 6902 84306 6924
rect 83709 6896 83936 6902
rect 83051 6891 83950 6896
rect 84134 6891 84309 6902
rect 84315 6897 84361 6952
rect 84368 6902 84389 6956
rect 84321 6891 84355 6897
rect 84367 6891 84967 6902
rect 84979 6891 85013 6971
rect 85442 6912 86434 6971
rect 86462 6940 90787 6971
rect 86462 6912 86496 6940
rect 85025 6891 85134 6902
rect 85442 6891 86530 6912
rect 86610 6906 90787 6940
rect 86604 6904 90787 6906
rect 86591 6891 90787 6904
rect 82440 6829 82521 6876
rect 82580 6857 90787 6891
rect 82992 6845 82993 6846
rect 83005 6845 83039 6857
rect 83051 6845 83052 6846
rect 82993 6844 82994 6845
rect 83005 6844 83051 6845
rect 82487 6261 82521 6829
rect 83005 6246 83050 6844
rect 83248 6836 83950 6857
rect 84321 6851 84355 6857
rect 83112 6776 83122 6802
rect 83084 6748 83122 6774
rect 83248 6624 83606 6836
rect 83629 6774 83634 6816
rect 83657 6774 83662 6816
rect 83663 6246 83708 6836
rect 84287 6816 84306 6851
rect 84308 6845 84309 6846
rect 84315 6845 84361 6851
rect 84368 6846 84389 6851
rect 84367 6845 84389 6846
rect 84966 6845 84967 6846
rect 84979 6845 85013 6857
rect 85025 6845 85026 6846
rect 84309 6844 84310 6845
rect 84315 6844 84367 6845
rect 84315 6788 84366 6844
rect 84321 6246 84366 6788
rect 84368 6774 84389 6845
rect 84967 6844 84968 6845
rect 84979 6844 85025 6845
rect 84979 6246 85024 6844
rect 85442 6672 86434 6857
rect 86462 6672 86496 6857
rect 86610 6790 90787 6857
rect 86565 6779 90787 6790
rect 86576 6672 90787 6779
rect 85442 6472 90787 6672
rect 85442 6464 86758 6472
rect 82993 6245 82994 6246
rect 83005 6245 83051 6246
rect 83651 6245 83652 6246
rect 83663 6245 83709 6246
rect 84309 6245 84310 6246
rect 84321 6245 84367 6246
rect 84967 6245 84968 6246
rect 84979 6245 85025 6246
rect 85610 6245 85682 6464
rect 85724 6326 85785 6464
rect 85800 6336 86070 6464
rect 86310 6460 86758 6464
rect 85724 6322 85792 6326
rect 82992 6244 82993 6245
rect 82936 6233 82993 6244
rect 83005 6233 83039 6245
rect 83051 6244 83052 6245
rect 83650 6244 83651 6245
rect 83051 6233 83651 6244
rect 83663 6233 83697 6245
rect 83709 6244 83710 6245
rect 84308 6244 84309 6245
rect 83709 6233 83936 6244
rect 84134 6233 84309 6244
rect 84321 6233 84355 6245
rect 84367 6244 84368 6245
rect 84966 6244 84967 6245
rect 84367 6233 84967 6244
rect 84979 6233 85013 6245
rect 85025 6244 85026 6245
rect 85610 6244 85678 6245
rect 85025 6233 85134 6244
rect 85428 6233 85678 6244
rect 85724 6244 85785 6322
rect 86382 6246 86427 6460
rect 86428 6374 86440 6460
rect 86462 6442 86496 6460
rect 86818 6442 86852 6472
rect 87040 6458 87085 6472
rect 87268 6458 90787 6472
rect 86462 6408 86852 6442
rect 86370 6245 86371 6246
rect 86382 6245 86428 6246
rect 86369 6244 86370 6245
rect 85724 6233 86370 6244
rect 86382 6233 86416 6245
rect 86428 6244 86429 6245
rect 86448 6244 86870 6358
rect 86944 6280 90787 6458
rect 86970 6254 87034 6267
rect 86944 6244 86970 6254
rect 87000 6248 87034 6254
rect 87040 6248 87130 6280
rect 87040 6246 87085 6248
rect 87028 6245 87029 6246
rect 87040 6245 87086 6246
rect 87027 6244 87028 6245
rect 86428 6233 86440 6244
rect 86448 6239 87028 6244
rect 87040 6239 87080 6245
rect 87086 6244 87087 6245
rect 87268 6244 90787 6280
rect 87086 6239 90787 6244
rect 86448 6233 87034 6239
rect 87040 6233 87074 6239
rect 87080 6233 90787 6239
rect 82440 6171 82521 6218
rect 82580 6199 90787 6233
rect 82992 6187 82993 6188
rect 83005 6187 83039 6199
rect 83051 6187 83052 6188
rect 83650 6187 83651 6188
rect 83663 6187 83697 6199
rect 83709 6187 83710 6188
rect 84308 6187 84309 6188
rect 84321 6187 84355 6199
rect 84367 6187 84368 6188
rect 84966 6187 84967 6188
rect 84979 6187 85013 6199
rect 85025 6187 85026 6188
rect 85610 6187 85678 6199
rect 82993 6186 82994 6187
rect 83005 6186 83051 6187
rect 83651 6186 83652 6187
rect 83663 6186 83709 6187
rect 84309 6186 84310 6187
rect 84321 6186 84367 6187
rect 84967 6186 84968 6187
rect 84979 6186 85025 6187
rect 82487 6052 82521 6171
rect 83005 6052 83050 6186
rect 83566 6116 83570 6166
rect 83594 6116 83598 6138
rect 83663 6052 83708 6186
rect 84321 6052 84366 6186
rect 84979 6052 85024 6186
rect 78880 5996 78914 6030
rect 79538 6004 79572 6038
rect 80196 6004 80230 6038
rect 80854 6012 80888 6046
rect 78100 5962 79020 5996
rect 78066 5900 78068 5934
rect 76910 4648 77830 4682
rect 78100 4682 78142 5962
rect 78222 5910 78267 5962
rect 78692 5932 78726 5962
rect 78222 5822 78268 5910
rect 78692 5894 78730 5932
rect 78806 5894 78840 5962
rect 78880 5956 78914 5962
rect 78874 5932 78914 5956
rect 78844 5894 78914 5932
rect 78276 5860 78914 5894
rect 78222 5821 78267 5822
rect 78203 5810 78267 5821
rect 78214 4834 78267 5810
rect 78222 4822 78267 4834
rect 78692 4822 78726 5860
rect 78806 5156 78840 5860
rect 78846 5854 78856 5860
rect 78874 5826 78914 5860
rect 78872 5822 78914 5826
rect 78866 5821 78914 5822
rect 78861 5810 78914 5821
rect 78866 5798 78914 5810
rect 78806 4846 78862 5156
rect 78872 4846 78914 5798
rect 78222 4734 78268 4822
rect 78692 4784 78730 4822
rect 78806 4784 78840 4846
rect 78866 4822 78914 4846
rect 78844 4784 78914 4822
rect 78276 4750 78914 4784
rect 78222 4682 78267 4734
rect 78692 4686 78726 4750
rect 78692 4682 78737 4686
rect 78806 4682 78840 4750
rect 78846 4744 78856 4750
rect 78874 4688 78914 4750
rect 78880 4682 78914 4688
rect 78986 4682 79020 5962
rect 78100 4648 79020 4682
rect 79410 5970 80330 6004
rect 76676 3456 76690 4034
rect 76676 3400 76716 3456
rect 77376 3402 77410 4648
rect 77508 3402 77548 3450
rect 77970 3402 77996 4026
rect 77998 3402 78024 3998
rect 78104 3402 78106 3998
rect 78108 3402 78142 4648
rect 78222 3402 78267 4648
rect 78692 3402 78737 4648
rect 78806 3402 78840 4648
rect 79410 4090 79444 5970
rect 79538 5918 79572 5970
rect 80154 5936 80192 5940
rect 79448 5568 79454 5854
rect 79538 5830 79584 5918
rect 80154 5902 80194 5936
rect 79586 5868 80194 5902
rect 80162 5862 80166 5868
rect 80190 5834 80194 5868
rect 79476 5596 79482 5826
rect 79513 5818 79526 5829
rect 79538 5818 79572 5830
rect 80171 5818 80184 5829
rect 80196 5818 80230 5970
rect 79524 4242 79572 5818
rect 80182 4242 80230 5818
rect 79538 4230 79572 4242
rect 79538 4142 79584 4230
rect 80154 4226 80192 4230
rect 80154 4192 80194 4226
rect 79586 4158 80194 4192
rect 80162 4152 80166 4158
rect 79538 4090 79572 4142
rect 80190 4124 80194 4158
rect 80196 4090 80230 4242
rect 80296 4090 80330 5970
rect 79410 4056 80330 4090
rect 80578 5978 81498 6012
rect 80578 4098 80612 5978
rect 80854 5926 80892 5948
rect 80842 5910 80900 5926
rect 81322 5910 81360 5948
rect 80754 5876 81360 5910
rect 80722 5837 80776 5870
rect 80681 5826 80776 5837
rect 80692 4250 80776 5826
rect 80722 4206 80776 4250
rect 80778 4206 80804 5870
rect 80842 5838 80900 5876
rect 80854 4238 80888 5838
rect 81339 5826 81384 5837
rect 81350 4250 81384 5826
rect 80842 4200 80900 4238
rect 81322 4200 81360 4238
rect 80754 4166 81360 4200
rect 80842 4150 80900 4166
rect 80854 4098 80888 4150
rect 81464 4098 81498 5978
rect 81512 4104 81532 6046
rect 82197 5575 85326 6052
rect 85610 5587 85682 6187
rect 85610 5586 85678 5587
rect 85428 5575 85678 5586
rect 85724 5586 85785 6199
rect 86369 6187 86370 6188
rect 86382 6187 86416 6199
rect 86428 6187 86429 6188
rect 86370 6186 86371 6187
rect 86382 6186 86428 6187
rect 86382 5588 86427 6186
rect 86448 5738 86870 6199
rect 86944 6193 87034 6199
rect 87040 6193 87074 6199
rect 87080 6193 87130 6199
rect 87027 6187 87028 6188
rect 87040 6187 87080 6193
rect 87086 6187 87087 6188
rect 87028 6186 87029 6187
rect 87040 6186 87086 6187
rect 87040 6144 87085 6186
rect 87040 6137 87130 6144
rect 87040 5742 87085 6137
rect 87040 5656 87112 5742
rect 86480 5596 86600 5609
rect 87012 5596 87034 5609
rect 87040 5588 87085 5656
rect 86370 5587 86371 5588
rect 86382 5587 86428 5588
rect 87028 5587 87029 5588
rect 87040 5587 87086 5588
rect 86369 5586 86370 5587
rect 85724 5575 86370 5586
rect 86382 5575 86416 5587
rect 86428 5586 86429 5587
rect 87027 5586 87028 5587
rect 86428 5575 86440 5586
rect 86600 5581 87028 5586
rect 86600 5575 87034 5581
rect 87040 5575 87074 5587
rect 87086 5586 87087 5587
rect 87268 5586 90787 6199
rect 87086 5575 90787 5586
rect 82197 5541 90787 5575
rect 82197 4928 85326 5541
rect 85610 5535 85718 5541
rect 85724 5535 85816 5541
rect 85610 5529 85678 5535
rect 85610 5516 85682 5529
rect 85724 5516 85785 5535
rect 86369 5529 86370 5530
rect 86382 5529 86416 5541
rect 86428 5529 86429 5530
rect 87027 5529 87028 5530
rect 87040 5529 87074 5541
rect 87086 5529 87087 5530
rect 86370 5528 86371 5529
rect 86382 5528 86428 5529
rect 87028 5528 87029 5529
rect 87040 5528 87086 5529
rect 85610 5507 85718 5516
rect 85724 5507 85788 5516
rect 85610 5454 85705 5507
rect 85610 4962 85682 5454
rect 85724 5123 85785 5507
rect 86382 5123 86427 5528
rect 87040 5123 87085 5528
rect 85751 5111 85785 5123
rect 87268 5111 90787 5541
rect 85739 5064 86401 5111
rect 86600 5064 90787 5111
rect 85751 4962 85785 5064
rect 85786 5030 86401 5064
rect 86444 5052 87059 5064
rect 87102 5052 90787 5064
rect 86444 5048 90787 5052
rect 90822 5048 90856 8426
rect 91204 6000 91206 6239
rect 91210 5098 91244 8274
rect 151698 7892 151790 8476
rect 152226 8080 152690 8476
rect 152226 7890 152704 8080
rect 152708 8028 152764 8046
rect 152818 8028 152870 8046
rect 100494 6240 100528 7812
rect 108672 7136 108674 7760
rect 108706 7148 108708 7748
rect 152666 7448 152704 7890
rect 152726 7508 152764 8020
rect 152818 8000 152842 8018
rect 152888 7890 153876 8476
rect 101276 6496 101628 6582
rect 101276 6478 102024 6496
rect 108672 6478 108674 7102
rect 108706 6490 108708 7090
rect 100800 6444 108656 6478
rect 154330 6464 155190 8484
rect 155366 6472 156358 8492
rect 156526 8262 157954 8496
rect 156526 7934 157976 8262
rect 101276 6422 102024 6444
rect 101276 6308 101628 6422
rect 99768 6206 103224 6240
rect 100494 6172 100528 6206
rect 100472 6138 100528 6172
rect 100596 6138 100630 6206
rect 101074 6138 101112 6176
rect 101732 6138 101770 6176
rect 102390 6138 102428 6176
rect 103048 6138 103086 6176
rect 100494 6104 101112 6138
rect 101164 6104 101770 6138
rect 101822 6104 102428 6138
rect 102480 6104 103086 6138
rect 100476 6062 100484 6066
rect 100494 6062 100528 6104
rect 100410 6000 100436 6062
rect 100476 6000 100528 6062
rect 97356 5312 97373 5344
rect 97356 5242 97374 5312
rect 86444 5030 91866 5048
rect 86980 5028 91866 5030
rect 87268 5024 91866 5028
rect 86450 5006 86706 5022
rect 86980 5014 91866 5024
rect 86478 4978 86678 4994
rect 86980 4972 90787 5014
rect 87268 4962 90787 4972
rect 85610 4946 90787 4962
rect 90822 4946 90856 5014
rect 85610 4928 91262 4946
rect 82197 4917 85625 4928
rect 85637 4917 85671 4928
rect 85751 4917 85785 4928
rect 82197 4883 85819 4917
rect 87268 4912 91262 4928
rect 82197 4259 85326 4883
rect 85624 4871 85625 4872
rect 85637 4871 85671 4883
rect 85625 4870 85626 4871
rect 85637 4444 85682 4871
rect 85625 4271 85626 4272
rect 85624 4270 85625 4271
rect 85637 4259 85671 4444
rect 85751 4259 85785 4883
rect 86478 4794 86678 4812
rect 86450 4766 86706 4784
rect 82197 4225 85785 4259
rect 80578 4064 81498 4098
rect 78890 3470 78914 3628
rect 78928 3508 78952 3590
rect 79224 3402 79686 3534
rect 79700 3402 80162 3534
rect 80762 3406 80776 4054
rect 80854 3406 80888 4064
rect 81814 3508 81834 3590
rect 81852 3470 81872 3628
rect 82197 3612 85326 4225
rect 85624 4213 85625 4214
rect 85625 4212 85626 4213
rect 85637 3846 85671 4225
rect 85625 3613 85626 3614
rect 85637 3613 85682 3846
rect 85624 3612 85625 3613
rect 82197 3601 85625 3612
rect 85637 3601 85671 3613
rect 85751 3601 85785 4225
rect 87268 3660 90787 4912
rect 82197 3567 85819 3601
rect 85821 3567 90787 3660
rect 90822 3567 90856 4912
rect 98796 4604 98854 4634
rect 98830 4570 98854 4600
rect 96298 4398 96680 4498
rect 95512 4026 96692 4398
rect 100494 4390 100528 6000
rect 100596 5848 100630 6104
rect 100668 6066 100669 6067
rect 100667 6065 100668 6066
rect 101091 6054 101136 6065
rect 101749 6054 101794 6065
rect 102407 6054 102452 6065
rect 103065 6054 103110 6065
rect 101090 5832 101091 5833
rect 101089 5831 101090 5832
rect 101102 5820 101136 6054
rect 101147 5832 101148 5833
rect 101748 5832 101749 5833
rect 101148 5831 101149 5832
rect 101747 5831 101748 5832
rect 101760 5820 101794 6054
rect 101805 5832 101806 5833
rect 102406 5832 102407 5833
rect 101806 5831 101807 5832
rect 102405 5831 102406 5832
rect 102418 5820 102452 6054
rect 102463 5832 102464 5833
rect 103064 5832 103065 5833
rect 102464 5831 102465 5832
rect 103063 5831 103064 5832
rect 103076 5820 103110 6054
rect 103190 5820 103224 6206
rect 107928 5904 107984 5916
rect 108672 5820 108674 6444
rect 108706 5832 108708 6432
rect 154506 6294 154520 6464
rect 154534 6322 154548 6464
rect 100558 5758 100630 5796
rect 100680 5786 103224 5820
rect 101089 5774 101090 5775
rect 101090 5773 101091 5774
rect 100596 5346 100630 5758
rect 101102 5346 101136 5786
rect 101148 5774 101149 5775
rect 101747 5774 101748 5775
rect 101147 5773 101148 5774
rect 101748 5773 101749 5774
rect 101760 5346 101794 5786
rect 101806 5774 101807 5775
rect 102405 5774 102406 5775
rect 101805 5773 101806 5774
rect 102406 5773 102407 5774
rect 102418 5346 102452 5786
rect 102464 5774 102465 5775
rect 103063 5774 103064 5775
rect 102463 5773 102464 5774
rect 103064 5773 103065 5774
rect 100596 5190 100668 5346
rect 101102 5175 101147 5346
rect 101760 5252 101805 5346
rect 102418 5252 102463 5346
rect 101310 5180 102490 5252
rect 101362 5175 102463 5180
rect 101090 5174 101091 5175
rect 101102 5174 101148 5175
rect 101362 5174 102464 5175
rect 103064 5174 103065 5175
rect 101089 5173 101090 5174
rect 100669 5162 101090 5173
rect 101102 5162 101136 5174
rect 101148 5173 101149 5174
rect 101362 5173 102452 5174
rect 101148 5162 102452 5173
rect 102464 5173 102465 5174
rect 103063 5173 103064 5174
rect 102464 5162 103008 5173
rect 103076 5162 103110 5786
rect 103190 5162 103224 5786
rect 107928 5724 107984 5744
rect 107928 5668 107984 5688
rect 108672 5162 108674 5786
rect 108706 5224 108708 5774
rect 108700 5202 108724 5224
rect 108700 5178 108746 5202
rect 108706 5174 108708 5178
rect 100558 5100 100668 5138
rect 100680 5128 108656 5162
rect 101089 5116 101090 5117
rect 101102 5116 101136 5128
rect 101148 5116 101149 5117
rect 101362 5116 102452 5128
rect 102464 5116 102465 5117
rect 103063 5116 103064 5117
rect 101090 5115 101091 5116
rect 101102 5115 101148 5116
rect 101362 5115 102464 5116
rect 103064 5115 103065 5116
rect 100596 4532 100668 5100
rect 101102 4517 101147 5115
rect 101362 5106 102463 5115
rect 101310 4880 102490 5106
rect 101760 4517 101805 4880
rect 102418 4517 102463 4880
rect 101090 4516 101091 4517
rect 101102 4516 101148 4517
rect 101748 4516 101749 4517
rect 101760 4516 101806 4517
rect 102406 4516 102407 4517
rect 102418 4516 102464 4517
rect 101089 4515 101090 4516
rect 100669 4504 101090 4515
rect 101102 4504 101136 4516
rect 101148 4515 101149 4516
rect 101747 4515 101748 4516
rect 101148 4504 101748 4515
rect 101760 4504 101794 4516
rect 101806 4515 101807 4516
rect 102405 4515 102406 4516
rect 101806 4504 102406 4515
rect 102418 4504 102452 4516
rect 102464 4515 102465 4516
rect 103042 4515 103066 4600
rect 102464 4504 103066 4515
rect 103076 4504 103110 5128
rect 103190 4504 103224 5128
rect 108672 4504 108674 5128
rect 108706 4516 108708 5116
rect 153864 4956 153890 5880
rect 153898 4956 153924 5846
rect 155796 5123 155830 6472
rect 156500 5030 156516 5064
rect 156526 4892 157954 7934
rect 163643 7406 163677 10465
rect 163838 10413 163884 10444
rect 163826 10397 163884 10413
rect 163819 10363 163884 10397
rect 163826 10316 163884 10363
rect 163746 10304 163791 10315
rect 163757 7555 163791 10304
rect 163838 7567 163872 10316
rect 163745 7508 163804 7555
rect 163810 7508 163857 7555
rect 163745 7474 163857 7508
rect 163745 7458 163803 7474
rect 163745 7443 163760 7458
rect 163757 7406 163791 7440
rect 163952 7406 163986 10465
rect 161280 7372 163986 7406
rect 100680 4470 103224 4504
rect 101102 4390 101136 4470
rect 101760 4390 101794 4470
rect 102418 4390 102452 4470
rect 103076 4390 103110 4470
rect 103190 4390 103224 4470
rect 100494 4356 108746 4390
rect 97308 4062 98300 4074
rect 98476 4056 99468 4074
rect 82197 3534 85326 3567
rect 82044 3487 85326 3534
rect 85637 3487 85671 3567
rect 85751 3487 85785 3567
rect 85821 3531 90892 3567
rect 85821 3497 92143 3531
rect 85821 3487 90892 3497
rect 82044 3453 90892 3487
rect 91372 3476 91570 3497
rect 91368 3467 91570 3476
rect 91848 3467 92046 3497
rect 76648 3200 76660 3400
rect 76676 3200 76688 3400
rect 76676 3144 76716 3200
rect 76676 3056 76690 3144
rect 76676 3000 76716 3056
rect 76648 2800 76660 3000
rect 76676 2800 76688 3000
rect 76782 2896 80162 3402
rect 80272 2954 80284 3274
rect 80294 3238 81696 3406
rect 81702 3238 81944 3406
rect 76782 2862 79748 2896
rect 76676 2744 76716 2800
rect 76676 2632 76690 2744
rect 76776 2672 79748 2862
rect 76748 2632 79748 2672
rect 76748 2616 76752 2632
rect 76782 2464 79748 2632
rect 79754 2812 80104 2846
rect 76712 2364 76716 2400
rect 72650 2310 76625 2346
rect 76706 2330 76764 2364
rect 77364 2330 77422 2364
rect 72650 2305 78006 2310
rect 72650 2299 76717 2305
rect 76753 2299 77375 2305
rect 77411 2299 78006 2305
rect 72650 2287 76706 2299
rect 76764 2287 77364 2299
rect 77422 2287 78006 2299
rect 72650 2276 76717 2287
rect 76753 2276 77375 2287
rect 77411 2276 78006 2287
rect 71642 2167 72612 2268
rect 72650 2266 76625 2276
rect 72650 2242 76706 2266
rect 76764 2242 77364 2266
rect 77422 2242 77888 2266
rect 77972 2242 78006 2276
rect 72650 2224 76625 2242
rect 77508 2234 77870 2242
rect 72650 2214 77830 2224
rect 72650 2208 77842 2214
rect 72650 2190 76625 2208
rect 77480 2206 77842 2208
rect 77830 2190 77842 2206
rect 77858 2190 77870 2234
rect 77972 2231 77983 2242
rect 77995 2231 78006 2242
rect 78108 2292 78142 2464
rect 78222 2342 78267 2464
rect 78692 2342 78737 2464
rect 78806 2292 78840 2464
rect 79278 2332 79312 2464
rect 79398 2434 79508 2464
rect 79538 2446 79552 2464
rect 79436 2400 79508 2434
rect 79538 2342 79566 2366
rect 79594 2332 79628 2464
rect 78876 2298 78892 2326
rect 79278 2298 79628 2332
rect 79754 2332 79788 2812
rect 79874 2744 79984 2782
rect 79912 2710 79984 2744
rect 79857 2660 79913 2671
rect 79945 2660 80001 2671
rect 79868 2484 79913 2660
rect 79956 2484 80001 2660
rect 79874 2434 79984 2472
rect 79912 2400 79984 2434
rect 80070 2332 80104 2812
rect 80272 2480 80284 2768
rect 80294 2502 81944 3238
rect 82044 3370 85326 3453
rect 85751 3370 85785 3453
rect 85821 3417 90892 3453
rect 91276 3464 91666 3467
rect 91276 3436 91310 3464
rect 91340 3436 91356 3448
rect 91242 3435 91356 3436
rect 91368 3435 91384 3464
rect 91242 3429 91344 3435
rect 87268 3402 88108 3406
rect 88651 3402 90892 3417
rect 87268 3370 90892 3402
rect 91276 3370 91310 3429
rect 91394 3412 91421 3445
rect 91532 3435 91554 3464
rect 91560 3435 91582 3448
rect 91632 3436 91666 3464
rect 91752 3464 92101 3467
rect 91752 3436 91786 3464
rect 91598 3429 91700 3436
rect 91718 3429 91820 3436
rect 91976 3435 92008 3448
rect 92032 3435 92036 3464
rect 91356 3389 91368 3402
rect 91436 3396 91463 3412
rect 91340 3370 91356 3389
rect 91368 3370 91384 3389
rect 91436 3370 91490 3396
rect 91495 3395 91528 3429
rect 91554 3389 91560 3402
rect 91532 3370 91554 3389
rect 91560 3370 91582 3389
rect 91632 3370 91666 3429
rect 91752 3395 92063 3429
rect 91752 3370 91786 3395
rect 91928 3370 91966 3395
rect 92008 3389 92032 3395
rect 91976 3370 92008 3389
rect 92032 3370 92036 3389
rect 92108 3370 92133 3402
rect 82044 3336 92056 3370
rect 82044 2896 85326 3336
rect 85637 3284 85683 3315
rect 85625 3268 85683 3284
rect 85354 3234 85683 3268
rect 85625 3187 85683 3234
rect 82197 2846 85326 2896
rect 82098 2812 85326 2846
rect 82098 2502 82132 2812
rect 82197 2512 85326 2812
rect 85637 2512 85671 3187
rect 82197 2502 85337 2512
rect 79754 2298 80104 2332
rect 80294 2468 85337 2502
rect 80294 2432 81944 2468
rect 78108 2258 78840 2292
rect 78848 2270 78864 2298
rect 78942 2266 79510 2292
rect 78942 2258 79512 2266
rect 78108 2242 78142 2258
rect 78108 2231 78119 2242
rect 78131 2231 78142 2242
rect 78806 2242 78840 2258
rect 78806 2231 78817 2242
rect 78829 2231 78840 2242
rect 79560 2224 79576 2298
rect 79588 2252 79604 2298
rect 77972 2190 78006 2214
rect 80294 2190 81878 2432
rect 82098 2394 82132 2468
rect 82197 2432 85337 2468
rect 72650 2182 81878 2190
rect 82197 2262 82484 2432
rect 82530 2316 82960 2432
rect 83005 2328 83050 2432
rect 83188 2316 83233 2432
rect 83663 2328 83708 2432
rect 83756 2316 83780 2432
rect 83784 2316 83836 2432
rect 83846 2316 83891 2432
rect 82518 2269 83892 2316
rect 72650 2167 81696 2182
rect 70217 2156 81696 2167
rect 65212 2136 65270 2156
rect 65870 2136 65928 2156
rect 58029 2106 58048 2120
rect 58145 1844 58168 2000
rect 57968 1800 58168 1844
rect 58173 1788 58196 2028
rect 58772 1982 60254 2133
rect 57940 1772 58196 1788
rect 58180 1222 58213 1266
rect 58214 1256 58247 1266
rect 58837 -186 58871 1982
rect 58898 1690 58922 1792
rect 58942 1150 58976 1982
rect 59056 1311 59101 1982
rect 59495 1299 59540 1982
rect 60153 1299 60198 1982
rect 60811 1299 60856 2133
rect 61114 1311 61148 2133
rect 59071 1252 60898 1299
rect 61086 1252 61133 1299
rect 59118 1218 61133 1252
rect 59483 1202 59541 1218
rect 60141 1202 60199 1218
rect 60799 1202 60857 1218
rect 59495 1150 59529 1184
rect 60153 1150 60187 1184
rect 60811 1150 60845 1184
rect 61228 1150 61262 2133
rect 58942 1116 61262 1150
rect 61583 888 61617 2133
rect 62502 2097 64133 2133
rect 63136 1196 63170 2097
rect 63250 1336 63284 2097
rect 63908 1336 63942 2097
rect 64566 1336 64600 2136
rect 65224 1336 65269 2136
rect 65882 1336 65927 2136
rect 66492 1788 66512 2156
rect 66528 2136 66586 2156
rect 66282 1346 66286 1666
rect 66320 1346 66324 1666
rect 66540 1336 66585 2136
rect 63238 1298 63296 1336
rect 63896 1298 63954 1336
rect 64554 1298 64612 1336
rect 65138 1298 66586 1336
rect 63238 1264 66586 1298
rect 63238 1248 63296 1264
rect 63896 1248 63954 1264
rect 64554 1248 64612 1264
rect 65212 1248 65270 1264
rect 65870 1248 65928 1264
rect 66528 1248 66586 1264
rect 63238 1233 63253 1248
rect 66571 1233 66586 1248
rect 63250 1196 63284 1230
rect 63908 1196 63942 1230
rect 64566 1196 64600 1230
rect 65224 1196 65258 1230
rect 65882 1196 65916 1230
rect 66540 1196 66574 1230
rect 66654 1196 66688 2156
rect 67698 2131 67756 2136
rect 67824 1258 67858 2156
rect 69054 2120 69204 2156
rect 70217 2133 76625 2156
rect 77858 2140 77870 2156
rect 69090 1212 69124 2120
rect 69170 1364 69182 2120
rect 69204 1398 69216 2120
rect 69170 1261 69196 1364
rect 69204 1295 69230 1398
rect 71376 1212 71410 2133
rect 71642 2097 72612 2133
rect 72650 2097 76625 2133
rect 77846 2131 77904 2136
rect 76460 2000 76488 2097
rect 72086 1836 72158 1844
rect 72086 1834 72154 1836
rect 77972 1694 78006 2156
rect 80294 2120 81696 2156
rect 80758 2106 80920 2108
rect 82197 2097 82198 2262
rect 82369 2201 82396 2262
rect 82397 2229 82450 2262
rect 82416 2184 82450 2229
rect 82518 2235 83024 2269
rect 83067 2235 83682 2269
rect 82518 2222 82576 2235
rect 82518 2212 82596 2222
rect 83176 2212 83234 2235
rect 82480 2190 82596 2212
rect 83126 2206 83282 2212
rect 82518 2185 82576 2190
rect 83176 2185 83234 2206
rect 83687 2197 83694 2269
rect 83725 2235 83892 2269
rect 83834 2229 83892 2235
rect 83756 2194 83780 2229
rect 83784 2222 83892 2229
rect 83818 2212 83892 2222
rect 83818 2196 83912 2212
rect 83820 2188 83910 2196
rect 83834 2185 83892 2188
rect 82408 2172 82628 2184
rect 83126 2172 83282 2184
rect 83780 2173 83784 2184
rect 83790 2172 83940 2184
rect 82408 2168 83940 2172
rect 82408 2167 83938 2168
rect 83960 2167 83994 2432
rect 84520 2184 84554 2432
rect 84634 2316 84679 2432
rect 84979 2328 85024 2432
rect 85292 2316 85337 2432
rect 85637 2328 85682 2512
rect 84622 2269 85656 2316
rect 84622 2235 84998 2269
rect 85041 2235 85656 2269
rect 84622 2219 84680 2235
rect 85280 2219 85338 2235
rect 84622 2204 84637 2219
rect 84398 2167 84628 2184
rect 84634 2167 84668 2201
rect 84674 2167 84734 2184
rect 85230 2167 85286 2184
rect 85292 2167 85326 2201
rect 85332 2167 85384 2184
rect 85751 2167 85785 3336
rect 86514 3228 86668 3336
rect 87062 3332 90892 3336
rect 87268 3315 90892 3332
rect 91276 3315 91310 3336
rect 91433 3315 91479 3336
rect 91632 3315 91666 3336
rect 91752 3315 91786 3336
rect 92008 3333 92056 3336
rect 86966 3284 86977 3295
rect 86989 3284 87000 3295
rect 86966 3268 87000 3284
rect 87268 3268 91820 3315
rect 91866 3314 91913 3315
rect 92022 3314 92056 3333
rect 91855 3303 91913 3314
rect 91983 3303 92056 3314
rect 91866 3302 91913 3303
rect 91866 3268 91914 3302
rect 86966 3264 87238 3268
rect 87268 3264 91269 3268
rect 86966 3234 91269 3264
rect 86514 3214 86688 3228
rect 86656 3194 86688 3214
rect 86656 3176 86682 3194
rect 82329 2138 85785 2167
rect 82329 2133 83198 2138
rect 83212 2133 85785 2138
rect 82416 2098 82450 2133
rect 83250 2104 83818 2133
rect 83960 2098 83994 2133
rect 80796 2068 80882 2070
rect 81074 2004 81572 2032
rect 84520 1970 84554 2133
rect 85950 1970 85984 3175
rect 86584 3010 86682 3176
rect 86712 3171 86716 3228
rect 86584 2996 86662 3010
rect 86582 2826 86750 2996
rect 85990 2368 86610 2790
rect 86626 2352 86642 2810
rect 86966 2776 87000 3234
rect 87142 3230 90892 3234
rect 87268 3187 90892 3230
rect 87254 3183 90892 3187
rect 91276 3209 91310 3268
rect 91312 3234 91914 3268
rect 91276 3186 91318 3209
rect 87069 3171 87114 3182
rect 87255 3175 90892 3183
rect 91239 3175 91318 3186
rect 87080 2776 87114 3171
rect 86660 2742 87226 2776
rect 86660 2420 86694 2742
rect 86966 2662 87000 2742
rect 87080 2679 87114 2742
rect 87192 2683 87226 2742
rect 87266 2683 90892 3175
rect 87031 2662 87042 2673
rect 86715 2600 86796 2647
rect 86855 2628 87042 2662
rect 86762 2562 86796 2600
rect 86966 2534 87000 2628
rect 87043 2600 87124 2647
rect 87192 2636 90892 2683
rect 87126 2602 90892 2636
rect 87090 2546 87124 2600
rect 87031 2534 87042 2545
rect 87192 2534 87226 2602
rect 87254 2586 90892 2602
rect 87266 2534 90892 2586
rect 86855 2500 90892 2534
rect 87192 2420 87226 2500
rect 86660 2386 87226 2420
rect 87266 2464 90892 2500
rect 86528 2238 86536 2268
rect 86556 2238 86564 2240
rect 86684 2038 86700 2238
rect 86712 2010 86728 2266
rect 87266 2120 88108 2464
rect 88651 2140 90892 2464
rect 91250 3028 91318 3175
rect 91390 3187 91467 3234
rect 91390 3127 91424 3187
rect 91399 3111 91424 3127
rect 91433 3115 91467 3187
rect 91518 3127 91552 3234
rect 91433 3102 91479 3115
rect 91418 3068 91479 3102
rect 91490 3068 91537 3115
rect 91433 3034 91537 3068
rect 91250 2966 91310 3028
rect 91433 3018 91479 3034
rect 91433 2966 91467 3018
rect 91632 2966 91666 3234
rect 91250 2932 91666 2966
rect 91752 2966 91786 3234
rect 91866 3186 91900 3234
rect 91908 3186 91934 3191
rect 91866 3175 91942 3186
rect 91866 3127 91900 3175
rect 91874 3111 91900 3127
rect 91908 3102 91942 3175
rect 91994 3127 92056 3303
rect 91894 3068 91942 3102
rect 91966 3068 92013 3115
rect 91908 3034 92013 3068
rect 91908 2966 91942 3034
rect 92022 2966 92056 3127
rect 92108 3028 92159 3370
rect 92108 2966 92137 3028
rect 92205 2990 92239 3435
rect 92274 3404 92275 3567
rect 94844 3536 94878 3964
rect 94958 3536 94992 3570
rect 95616 3536 95650 3570
rect 95730 3536 95764 3964
rect 96034 3536 96068 3964
rect 96148 3536 96182 3570
rect 96806 3536 96840 3570
rect 96920 3536 96954 3964
rect 93854 3502 97214 3536
rect 94844 3406 94878 3502
rect 95610 3472 95612 3476
rect 94946 3406 95198 3472
rect 95212 3434 95662 3472
rect 95250 3406 95662 3434
rect 95730 3406 95764 3502
rect 96034 3406 96068 3502
rect 96136 3406 96514 3472
rect 96528 3434 96852 3472
rect 96566 3406 96852 3434
rect 96920 3406 96954 3502
rect 97344 3406 97364 3590
rect 98230 3406 98264 3424
rect 92528 2990 92529 3404
rect 93722 2990 94178 3404
rect 94632 3402 98264 3406
rect 94452 3394 94514 3402
rect 94580 3394 98264 3402
rect 92182 2966 94178 2990
rect 91752 2932 92137 2966
rect 91250 2882 91284 2932
rect 91433 2882 91467 2932
rect 91908 2882 91942 2932
rect 92022 2882 92056 2932
rect 91250 2830 91680 2882
rect 91734 2830 92156 2882
rect 91250 2684 92156 2830
rect 91250 2262 91680 2684
rect 91734 2262 92156 2684
rect 91250 2199 91295 2262
rect 91433 2187 91528 2262
rect 91908 2199 91953 2262
rect 90910 2140 91927 2187
rect 88651 2120 91269 2140
rect 87266 1970 87300 2120
rect 90478 2038 90512 2120
rect 90654 2106 91269 2120
rect 91312 2106 91927 2140
rect 90763 2090 90821 2106
rect 91421 2090 91479 2106
rect 91976 2038 92008 2048
rect 92022 2038 92056 2262
rect 90478 2004 92056 2038
rect 87302 1970 87334 2002
rect 82380 1966 84030 1970
rect 75760 1298 78042 1694
rect 78550 1528 79776 1562
rect 81342 1558 81356 1586
rect 72862 1264 78042 1298
rect 62634 1162 67762 1196
rect 58882 852 61653 888
rect 63136 852 63170 1162
rect 63250 852 63284 886
rect 63908 852 63942 886
rect 64566 852 64600 886
rect 65224 852 65258 886
rect 65882 852 65916 886
rect 66540 852 66574 886
rect 66654 852 66688 1162
rect 75760 1126 78042 1264
rect 71950 874 71984 886
rect 72108 880 72142 899
rect 79146 888 79180 1469
rect 81342 1266 81356 1456
rect 81342 1258 81366 1266
rect 81330 1256 81366 1258
rect 81342 1224 81366 1256
rect 81304 1222 81366 1224
rect 81342 1192 81366 1222
rect 72266 874 72300 886
rect 75760 852 78068 888
rect 58882 818 78068 852
rect 58882 166 61653 818
rect 63136 738 63170 818
rect 63250 738 63284 818
rect 63908 738 63942 818
rect 64566 738 64600 818
rect 65224 738 65258 818
rect 65882 738 65916 818
rect 66540 738 66574 818
rect 66654 738 66688 818
rect 71950 778 72300 804
rect 69218 756 69266 772
rect 63136 704 66688 738
rect 63136 280 63170 704
rect 63250 280 63284 704
rect 63296 692 63297 693
rect 63895 692 63896 693
rect 63295 691 63296 692
rect 63896 691 63897 692
rect 63295 292 63296 293
rect 63896 292 63897 293
rect 63296 291 63297 292
rect 63895 291 63896 292
rect 63908 280 63942 704
rect 63954 692 63955 693
rect 64553 692 64554 693
rect 63953 691 63954 692
rect 64554 691 64555 692
rect 63953 292 63954 293
rect 64554 292 64555 293
rect 63954 291 63955 292
rect 64553 291 64554 292
rect 64566 280 64600 704
rect 64612 692 64613 693
rect 65211 692 65212 693
rect 64611 691 64612 692
rect 65212 691 65213 692
rect 64611 292 64612 293
rect 65212 292 65213 293
rect 64612 291 64613 292
rect 65211 291 65212 292
rect 65224 280 65258 704
rect 65270 692 65271 693
rect 65869 692 65870 693
rect 65269 691 65270 692
rect 65870 691 65871 692
rect 65269 292 65270 293
rect 65870 292 65871 293
rect 65270 291 65271 292
rect 65869 291 65870 292
rect 65882 280 65916 704
rect 65928 692 65929 693
rect 66527 692 66528 693
rect 65927 691 65928 692
rect 66528 691 66529 692
rect 65927 292 65928 293
rect 66528 292 66529 293
rect 65928 291 65929 292
rect 66527 291 66528 292
rect 66540 280 66574 704
rect 66654 280 66688 704
rect 69066 723 69092 750
rect 69218 738 69232 756
rect 69240 738 69266 750
rect 75760 738 78068 818
rect 69096 723 69100 726
rect 67182 308 67766 322
rect 63136 246 66688 280
rect 69066 281 69100 723
rect 69232 723 69236 726
rect 69240 723 78068 738
rect 69232 704 78068 723
rect 69130 688 69164 692
rect 69124 608 69164 688
rect 69130 292 69164 608
rect 69168 292 69202 692
rect 69232 314 69266 704
rect 69066 258 69092 281
rect 69096 258 69100 281
rect 69218 281 69266 314
rect 69218 280 69236 281
rect 69232 258 69236 280
rect 69240 280 69266 281
rect 68978 246 69092 258
rect 63136 166 63170 246
rect 63250 166 63284 246
rect 63908 166 63942 246
rect 64566 166 64600 246
rect 65224 166 65258 246
rect 65882 166 65916 246
rect 66540 166 66574 246
rect 66654 166 66688 246
rect 69066 234 69092 246
rect 69240 246 69286 280
rect 75760 256 78068 704
rect 78338 262 79450 888
rect 79770 482 79798 600
rect 69240 234 69266 246
rect 69012 212 69066 224
rect 58882 132 79318 166
rect 58882 96 61653 132
rect 63136 0 63170 132
rect 66654 0 66688 132
rect 82408 92 82442 1838
rect 84484 1694 88108 1970
rect 88651 1700 90792 1970
rect 82884 532 84286 546
rect 84484 256 88216 1694
rect 88486 1576 90792 1700
rect 88486 1248 90809 1576
rect 90816 1286 90847 1538
rect 88486 262 90792 1248
rect 91433 877 91467 911
rect 91976 877 92008 2004
rect 92032 877 92036 2004
rect 92091 877 92125 911
rect 92205 877 92239 2966
rect 92528 1966 92529 2966
rect 93722 2713 94178 2966
rect 94632 2738 98264 3394
rect 98656 3346 98666 3958
rect 101102 3918 101122 3952
rect 100636 3884 101184 3918
rect 100636 3602 100670 3884
rect 101116 3822 101136 3856
rect 100811 3804 101009 3815
rect 101016 3810 101030 3818
rect 100700 3760 100810 3798
rect 100822 3770 101009 3804
rect 101012 3798 101030 3810
rect 101010 3760 101120 3798
rect 100738 3726 100810 3760
rect 100811 3716 101009 3727
rect 100822 3682 101009 3716
rect 101012 3678 101030 3760
rect 101040 3726 101120 3760
rect 101040 3706 101058 3726
rect 101090 3710 101098 3726
rect 101044 3684 101058 3706
rect 101102 3688 101120 3726
rect 101016 3656 101030 3678
rect 101102 3602 101122 3636
rect 101138 3602 101142 3608
rect 101150 3602 101184 3884
rect 100636 3568 101184 3602
rect 101234 3567 101872 3972
rect 98799 3429 99468 3567
rect 99636 3429 102899 3567
rect 98799 3395 102899 3429
rect 94632 2736 98256 2738
rect 94632 2713 98264 2736
rect 93336 2677 93370 2711
rect 93722 2704 98264 2713
rect 98512 2730 98546 2736
rect 98799 2730 99468 3395
rect 99514 3354 99542 3395
rect 99486 3346 99514 3354
rect 99542 3346 99570 3354
rect 99636 3347 102899 3395
rect 99514 3298 99542 3346
rect 99596 3336 102899 3347
rect 103070 3346 103072 3448
rect 98512 2718 99468 2730
rect 99607 2726 102899 3336
rect 103190 2788 103224 4356
rect 103190 2726 103224 2731
rect 99607 2718 103224 2726
rect 98512 2713 103224 2718
rect 93722 2682 98256 2704
rect 98512 2696 103260 2713
rect 98799 2682 103260 2696
rect 93722 2677 103260 2682
rect 103544 2677 103578 3684
rect 104310 3572 104324 3597
rect 103870 3536 107132 3572
rect 114018 3536 115391 3567
rect 103870 3502 107838 3536
rect 114018 3531 120330 3536
rect 109079 3502 120330 3531
rect 103870 3434 107132 3502
rect 109079 3497 115391 3502
rect 107254 3440 107282 3466
rect 107424 3450 107435 3461
rect 107447 3450 107458 3461
rect 107424 3434 107458 3450
rect 103870 3400 107458 3434
rect 103870 3361 107132 3400
rect 107226 3394 107254 3400
rect 103870 2713 107173 3361
rect 107254 3346 107282 3394
rect 107299 3350 107355 3361
rect 103658 2677 103692 2711
rect 103870 2682 107249 2713
rect 107310 2682 107355 3350
rect 107424 2682 107458 3400
rect 107702 3394 107770 3402
rect 107786 2682 107820 2716
rect 107900 2682 107934 3440
rect 111803 3429 111837 3467
rect 112501 3445 112512 3456
rect 112524 3445 112535 3456
rect 112501 3429 112535 3445
rect 109147 3389 109214 3402
rect 109662 3389 109739 3402
rect 109805 3389 109872 3402
rect 110320 3389 110397 3402
rect 111803 3395 112535 3429
rect 111803 2718 111837 3395
rect 111906 3336 111951 3347
rect 112376 3336 112421 3347
rect 111917 2718 111951 3336
rect 108947 2682 112320 2718
rect 103870 2677 112320 2682
rect 93037 2668 112320 2677
rect 93037 2643 97346 2668
rect 93037 2036 93071 2643
rect 93513 2622 93547 2643
rect 93722 2622 97346 2643
rect 93166 2575 97346 2622
rect 93213 2541 97346 2575
rect 93324 2494 93382 2541
rect 93140 2482 93196 2493
rect 93151 2185 93196 2482
rect 93336 2197 93381 2494
rect 93513 2185 93547 2541
rect 93616 2482 93672 2493
rect 93722 2482 97346 2541
rect 98072 2648 112320 2668
rect 98072 2522 98256 2648
rect 98799 2643 107249 2648
rect 98584 2580 98618 2627
rect 98799 2622 102172 2643
rect 102239 2622 102284 2643
rect 102353 2622 102387 2643
rect 98799 2580 102761 2622
rect 98584 2575 102761 2580
rect 98584 2546 102584 2575
rect 98584 2522 98618 2546
rect 98799 2541 102584 2546
rect 102627 2541 102761 2575
rect 98799 2522 102172 2541
rect 98072 2486 102172 2522
rect 93627 2226 97346 2482
rect 93627 2185 93672 2226
rect 93722 2185 97346 2226
rect 93139 2138 97346 2185
rect 93139 2104 93355 2138
rect 93398 2104 97346 2138
rect 93139 2088 93197 2104
rect 93139 2073 93154 2088
rect 93268 2036 93276 2098
rect 93513 2036 93547 2104
rect 93627 2036 93672 2104
rect 93688 2036 93716 2098
rect 93722 2036 97346 2104
rect 92660 2002 97346 2036
rect 93037 877 93071 2002
rect 93268 877 93276 2002
rect 93513 877 93547 2002
rect 93627 877 93672 2002
rect 93688 877 93716 2002
rect 93722 918 97346 2002
rect 97398 2452 102172 2486
rect 97398 2158 97432 2452
rect 98072 2400 102172 2452
rect 98060 2384 102172 2400
rect 97574 2350 102172 2384
rect 98060 2303 102172 2350
rect 97501 2291 97546 2302
rect 97398 1944 97454 2158
rect 97476 2000 97482 2158
rect 97398 1154 97432 1944
rect 97450 1676 97454 1944
rect 97450 1476 97456 1676
rect 97450 1247 97454 1476
rect 97512 1315 97546 2291
rect 97652 1766 97844 1818
rect 98072 1766 102172 2303
rect 97628 1698 102172 1766
rect 98072 1303 102172 1698
rect 98060 1256 102172 1303
rect 97574 1222 102172 1256
rect 98060 1206 102172 1222
rect 98072 1154 102172 1206
rect 97398 1120 102172 1154
rect 97408 918 97412 1120
rect 98072 1084 102172 1120
rect 98072 918 98256 1084
rect 93722 882 98256 918
rect 98584 882 98618 1084
rect 98698 882 98743 1084
rect 98774 882 102172 1084
rect 93722 877 102172 882
rect 102239 877 102284 2541
rect 102353 877 102387 2541
rect 102703 2494 102761 2541
rect 102554 2482 102610 2493
rect 102565 877 102610 2482
rect 102644 1638 102650 2158
rect 102672 1666 102706 2158
rect 102682 877 102706 1666
rect 102715 877 102760 2494
rect 102829 877 102863 2643
rect 103544 2575 103578 2643
rect 103661 2622 103695 2643
rect 103870 2622 107249 2643
rect 103646 2618 107249 2622
rect 107310 2618 107355 2648
rect 107424 2618 107458 2648
rect 103646 2615 107646 2618
rect 103627 2581 107646 2615
rect 103646 2575 107646 2581
rect 107660 2580 107832 2618
rect 103285 2546 107646 2575
rect 107698 2546 107832 2580
rect 103285 2541 107249 2546
rect 103223 877 103257 911
rect 103544 877 103578 2541
rect 103646 2494 103726 2541
rect 103658 877 103726 2494
rect 103764 2482 103820 2493
rect 103775 877 103820 2482
rect 103870 882 107249 2541
rect 107310 882 107355 2546
rect 107424 882 107458 2546
rect 107774 2508 107832 2546
rect 107625 2496 107681 2507
rect 107636 882 107681 2496
rect 107738 1988 107758 2158
rect 107710 1638 107728 1932
rect 107738 1666 107784 1988
rect 107762 882 107784 1666
rect 107786 882 107831 2508
rect 107900 882 107934 2648
rect 108732 2580 108766 2627
rect 108947 2580 112320 2648
rect 108732 2546 112320 2580
rect 108294 882 108328 916
rect 108732 882 108766 2546
rect 108947 2507 112320 2546
rect 108835 2496 108880 2507
rect 108941 2496 112320 2507
rect 108846 1970 108880 2496
rect 108846 882 108886 1970
rect 108912 882 108914 1914
rect 108947 882 112320 2496
rect 103870 877 112320 882
rect 80744 58 84200 92
rect 59495 -186 59529 0
rect 60153 -186 60187 0
rect 82408 -10 82442 58
rect 82510 -10 82544 0
rect 82708 -10 82746 28
rect 83366 -10 83404 28
rect 84024 -10 84062 28
rect 82408 -44 82746 -10
rect 82798 -44 83404 -10
rect 83456 -44 84062 -10
rect 80756 -88 80802 -82
rect 80756 -94 80828 -88
rect 80762 -106 80828 -94
rect 58772 -1762 60254 -186
rect 80796 -494 80828 -106
rect 80796 -1598 80802 -494
rect 80852 -522 80856 -60
rect 82072 -94 82118 -82
rect 82072 -106 82112 -94
rect 81480 -1542 81494 -1296
rect 81508 -1598 81550 -1296
rect 82072 -1342 82096 -434
rect 82408 -1584 82442 -44
rect 82510 -126 82544 -44
rect 82702 -70 82804 -54
rect 83360 -60 83462 -54
rect 83330 -70 83488 -60
rect 84018 -70 84120 -54
rect 82582 -82 82583 -81
rect 82581 -83 82582 -82
rect 82730 -83 82776 -82
rect 83388 -83 83434 -82
rect 84046 -83 84092 -82
rect 82725 -94 82776 -83
rect 83383 -88 83434 -83
rect 82730 -98 82776 -94
rect 83358 -98 83460 -88
rect 84041 -94 84092 -83
rect 84046 -98 84092 -94
rect 82724 -142 82725 -141
rect 82723 -143 82724 -142
rect 82736 -154 82770 -98
rect 82781 -142 82782 -141
rect 83382 -142 83383 -141
rect 82782 -143 82783 -142
rect 83381 -143 83382 -142
rect 83394 -154 83428 -98
rect 83439 -142 83440 -141
rect 84040 -142 84041 -141
rect 83440 -143 83441 -142
rect 84039 -143 84040 -142
rect 84052 -154 84086 -98
rect 84166 -154 84200 58
rect 82472 -216 82544 -178
rect 82594 -188 84200 -154
rect 82723 -200 82724 -199
rect 82724 -201 82725 -200
rect 82510 -784 82544 -216
rect 82724 -800 82725 -799
rect 82723 -801 82724 -800
rect 82736 -812 82770 -188
rect 82782 -200 82783 -199
rect 83381 -200 83382 -199
rect 82781 -201 82782 -200
rect 83382 -201 83383 -200
rect 82781 -800 82782 -799
rect 83382 -800 83383 -799
rect 82782 -801 82783 -800
rect 83381 -801 83382 -800
rect 83394 -812 83428 -188
rect 83440 -200 83441 -199
rect 84039 -200 84040 -199
rect 83439 -201 83440 -200
rect 84040 -201 84041 -200
rect 83439 -800 83440 -799
rect 84040 -800 84041 -799
rect 83440 -801 83441 -800
rect 84039 -801 84040 -800
rect 84052 -812 84086 -188
rect 84166 -812 84200 -188
rect 82472 -874 82544 -836
rect 82594 -846 84200 -812
rect 82723 -858 82724 -857
rect 82724 -859 82725 -858
rect 82510 -1442 82544 -874
rect 82724 -1458 82725 -1457
rect 82723 -1459 82724 -1458
rect 82736 -1470 82770 -846
rect 82782 -858 82783 -857
rect 83381 -858 83382 -857
rect 82781 -859 82782 -858
rect 83382 -859 83383 -858
rect 82781 -1458 82782 -1457
rect 83382 -1458 83383 -1457
rect 82782 -1459 82783 -1458
rect 83381 -1459 83382 -1458
rect 83394 -1470 83428 -846
rect 83440 -858 83441 -857
rect 84039 -858 84040 -857
rect 83439 -859 83440 -858
rect 84040 -859 84041 -858
rect 83439 -1458 83440 -1457
rect 84040 -1458 84041 -1457
rect 83440 -1459 83441 -1458
rect 84039 -1459 84040 -1458
rect 84052 -1470 84086 -846
rect 84166 -1470 84200 -846
rect 84484 -1032 88108 256
rect 88651 128 90792 262
rect 91169 848 112320 877
rect 91169 843 98256 848
rect 91169 128 91203 843
rect 91344 781 91356 843
rect 91433 791 91480 822
rect 91421 775 91480 791
rect 91913 775 91960 822
rect 91976 781 92008 843
rect 92032 794 92036 843
rect 92032 781 92064 794
rect 92091 791 92137 822
rect 92079 775 92137 791
rect 91345 741 91960 775
rect 92003 741 92137 775
rect 91272 682 91317 693
rect 91283 128 91317 682
rect 91344 128 91356 735
rect 91421 694 91479 741
rect 91433 128 91467 694
rect 91930 682 91975 693
rect 91941 128 91975 682
rect 91976 388 92008 735
rect 92032 444 92064 735
rect 92079 694 92137 741
rect 91976 128 92026 388
rect 92032 128 92082 444
rect 92091 128 92125 694
rect 92205 128 92239 843
rect 93037 128 93071 843
rect 93212 822 93220 843
rect 93268 837 93276 843
rect 93268 822 93297 837
rect 93513 822 93547 843
rect 93627 822 93672 843
rect 93688 822 93716 843
rect 93722 822 98256 843
rect 93139 818 98256 822
rect 98332 818 98368 842
rect 98584 818 98618 848
rect 98698 818 98743 848
rect 98774 843 107249 848
rect 98774 818 102172 843
rect 93139 786 102172 818
rect 93139 775 98340 786
rect 98352 782 102172 786
rect 102239 840 102284 843
rect 102239 782 102273 840
rect 102353 782 102387 843
rect 102565 840 102610 843
rect 102565 782 102599 840
rect 102632 836 102650 837
rect 102682 782 102706 843
rect 102715 840 102760 843
rect 102715 782 102749 840
rect 102829 782 102863 843
rect 103223 822 103257 843
rect 102922 782 103018 822
rect 98352 780 103018 782
rect 103195 809 103257 822
rect 103195 781 103263 809
rect 93139 741 93276 775
rect 93319 746 98340 775
rect 98390 775 103018 780
rect 103189 775 103263 781
rect 103273 775 103291 781
rect 103544 775 103578 843
rect 103658 775 103726 843
rect 103775 840 103820 843
rect 103775 822 103809 840
rect 103870 822 107249 843
rect 103775 791 103822 822
rect 103763 775 103822 791
rect 103853 818 107249 822
rect 107310 818 107355 848
rect 107424 818 107458 848
rect 107636 818 107681 848
rect 107702 828 107728 842
rect 107762 818 107784 848
rect 107786 818 107831 848
rect 107900 818 107934 848
rect 108294 818 108328 848
rect 103853 780 108674 818
rect 108732 780 108766 848
rect 108846 796 108886 848
rect 108912 814 108914 848
rect 108947 818 112320 848
rect 108924 814 112320 818
rect 108912 810 112320 814
rect 108834 786 108892 796
rect 108924 786 112320 810
rect 108834 780 112320 786
rect 103853 775 107681 780
rect 98390 748 103263 775
rect 98390 746 102599 748
rect 93319 741 98312 746
rect 93139 735 93241 741
rect 93268 735 93269 741
rect 93139 694 93220 735
rect 93268 694 93297 735
rect 93151 394 93220 694
rect 93251 693 93297 694
rect 93246 682 93302 693
rect 93251 394 93302 682
rect 93151 128 93196 394
rect 93257 128 93302 394
rect 93513 128 93547 741
rect 93627 128 93672 741
rect 93722 740 98312 741
rect 93722 708 98268 740
rect 98332 712 98340 746
rect 93722 706 98267 708
rect 93722 320 98256 706
rect 98317 696 98362 707
rect 98328 320 98362 696
rect 98584 320 98618 746
rect 98698 706 98743 746
rect 98799 741 102599 746
rect 102611 741 103263 748
rect 103269 746 107681 775
rect 107698 746 108334 780
rect 103269 741 107249 746
rect 98698 320 98732 706
rect 98799 680 102172 741
rect 102184 680 102231 727
rect 98799 646 102231 680
rect 102239 680 102273 741
rect 102353 680 102387 741
rect 102565 727 102599 741
rect 102632 735 102682 741
rect 102565 696 102612 727
rect 102553 680 102612 696
rect 102682 686 102688 735
rect 102715 727 102749 741
rect 102632 680 102682 686
rect 102715 680 102762 727
rect 102829 680 102863 741
rect 102239 646 102863 680
rect 93722 128 98772 320
rect 88651 80 98772 128
rect 88468 46 98772 80
rect 88468 -154 88502 46
rect 88651 -22 98772 46
rect 88644 -56 98772 -22
rect 88548 -70 88650 -66
rect 88576 -95 88622 -94
rect 88571 -98 88622 -95
rect 88571 -106 88616 -98
rect 88582 -154 88616 -106
rect 88620 -148 88638 -98
rect 88651 -154 98772 -56
rect 88434 -188 98772 -154
rect 88468 -812 88502 -188
rect 88582 -812 88616 -188
rect 88620 -286 88638 -194
rect 88651 -618 98772 -188
rect 98799 -448 102172 646
rect 102239 598 102273 646
rect 102201 587 102273 598
rect 102212 -389 102273 587
rect 102184 -448 102231 -401
rect 98799 -482 102231 -448
rect 102239 -448 102273 -389
rect 102353 -448 102387 646
rect 102553 599 102611 646
rect 102565 -134 102599 599
rect 102548 -448 102618 -134
rect 102715 -401 102749 646
rect 102829 598 102863 646
rect 102870 598 102897 603
rect 102829 587 102904 598
rect 102715 -448 102762 -401
rect 102829 -448 102863 587
rect 102870 -389 102904 587
rect 102870 -405 102897 -389
rect 102239 -482 102863 -448
rect 98799 -550 102172 -482
rect 102239 -530 102273 -482
rect 102239 -550 102284 -530
rect 102308 -550 102520 -482
rect 102548 -550 102618 -482
rect 102650 -488 102682 -482
rect 102682 -538 102706 -488
rect 102715 -530 102749 -482
rect 102650 -544 102682 -538
rect 102715 -550 102760 -530
rect 102829 -550 102863 -482
rect 102984 -550 103018 741
rect 103189 735 103207 741
rect 103217 707 103263 741
rect 103273 735 103291 741
rect 103223 6 103257 707
rect 103544 6 103578 741
rect 103658 98 103726 741
rect 103763 694 103821 741
rect 103775 196 103809 694
rect 103775 98 103820 196
rect 103658 16 103820 98
rect 103658 6 103726 16
rect 103775 6 103820 16
rect 103870 6 107249 741
rect 98799 -584 103018 -550
rect 103064 -28 103454 6
rect 103064 -526 103098 -28
rect 103206 -96 103223 -62
rect 103224 -96 103269 -80
rect 103278 -96 103325 -49
rect 103224 -130 103325 -96
rect 103224 -139 103269 -130
rect 103288 -138 103304 -130
rect 103172 -178 103186 -177
rect 103189 -178 103212 -173
rect 103167 -189 103212 -178
rect 103178 -365 103212 -189
rect 103172 -377 103186 -368
rect 103189 -381 103212 -365
rect 103223 -177 103269 -139
rect 103223 -377 103257 -177
rect 103295 -189 103340 -178
rect 103306 -365 103340 -189
rect 103223 -390 103269 -377
rect 103206 -415 103269 -390
rect 103206 -424 103223 -415
rect 103224 -416 103269 -415
rect 103278 -416 103325 -377
rect 103224 -458 103325 -416
rect 103224 -474 103269 -458
rect 103288 -498 103320 -458
rect 103316 -510 103320 -498
rect 103200 -512 103217 -510
rect 103263 -512 103320 -510
rect 103344 -526 103348 -391
rect 103420 -526 103454 -28
rect 103064 -560 103454 -526
rect 103540 -28 107249 6
rect 103540 -526 103578 -28
rect 103658 -96 103726 -28
rect 103775 -49 103809 -28
rect 103754 -96 103809 -49
rect 103658 -130 103809 -96
rect 103658 -178 103726 -130
rect 103643 -189 103726 -178
rect 103654 -331 103726 -189
rect 103627 -365 103726 -331
rect 103658 -391 103726 -365
rect 103775 -173 103809 -130
rect 103775 -189 103820 -173
rect 103775 -365 103816 -189
rect 103775 -377 103820 -365
rect 103754 -381 103820 -377
rect 103661 -526 103695 -391
rect 103754 -403 103809 -381
rect 103754 -424 103822 -403
rect 103700 -450 103822 -424
rect 103870 -450 107249 -28
rect 103700 -458 107249 -450
rect 103704 -484 107249 -458
rect 103775 -490 103809 -484
rect 103775 -526 103815 -490
rect 103832 -526 103843 -490
rect 103870 -526 107249 -484
rect 103540 -560 107249 -526
rect 88620 -806 88622 -734
rect 88627 -800 88628 -799
rect 88628 -801 88629 -800
rect 88651 -812 98267 -618
rect 88434 -846 98267 -812
rect 85968 -1242 86002 -1032
rect 86082 -1090 86116 -1032
rect 86740 -1090 86774 -1032
rect 86712 -1140 86750 -1102
rect 86144 -1174 86750 -1140
rect 86854 -1242 86888 -1032
rect 85968 -1276 86888 -1242
rect 87158 -1242 87192 -1032
rect 87272 -1090 87306 -1032
rect 87930 -1090 87964 -1032
rect 87902 -1140 87940 -1102
rect 87334 -1174 87940 -1140
rect 88044 -1242 88078 -1032
rect 87158 -1276 88078 -1242
rect 87330 -1386 87880 -1384
rect 87358 -1414 87852 -1412
rect 88468 -1470 88502 -846
rect 88582 -1470 88616 -846
rect 88620 -938 88622 -852
rect 88628 -858 88629 -857
rect 88627 -859 88628 -858
rect 88651 -1032 98267 -846
rect 98288 -956 98318 -618
rect 98288 -980 98290 -956
rect 98288 -990 98322 -980
rect 88620 -1464 88622 -1386
rect 88627 -1458 88628 -1457
rect 88628 -1459 88629 -1458
rect 88651 -1470 97101 -1032
rect 97108 -1392 97134 -1042
rect 97162 -1062 97207 -1032
rect 82594 -1504 97101 -1470
rect 82736 -1584 82770 -1504
rect 83394 -1584 83428 -1504
rect 84052 -1584 84086 -1504
rect 84166 -1584 84200 -1504
rect 88468 -1584 88502 -1504
rect 88582 -1584 88616 -1504
rect 88620 -1584 88622 -1510
rect 88651 -1584 97101 -1504
rect 82408 -1618 97101 -1584
rect 44808 -3988 44928 -3968
rect 45114 -3986 45354 -3434
rect 45114 -3988 45404 -3986
rect 44802 -4016 44956 -3996
rect 45114 -4014 45354 -3988
rect 45114 -4016 45432 -4014
rect 45114 -4072 45354 -4016
rect 58837 -4640 58871 -1762
rect 59495 -4640 59529 -1762
rect 60153 -4640 60187 -1762
rect 78236 -2484 78260 -1790
rect 78270 -2484 78294 -1824
rect 83310 -2002 83328 -1618
rect 83366 -2002 83384 -1670
rect 82550 -2090 83098 -2056
rect 82550 -2372 82584 -2090
rect 82736 -2170 82770 -2090
rect 82912 -2170 82923 -2159
rect 82614 -2214 82686 -2176
rect 82652 -2248 82686 -2214
rect 82736 -2204 82923 -2170
rect 82723 -2216 82724 -2215
rect 82724 -2217 82725 -2216
rect 82724 -2246 82725 -2245
rect 82723 -2247 82724 -2246
rect 82736 -2258 82770 -2204
rect 82924 -2214 82996 -2176
rect 82782 -2216 82783 -2215
rect 82781 -2217 82782 -2216
rect 82781 -2246 82782 -2245
rect 82782 -2247 82783 -2246
rect 82912 -2258 82923 -2247
rect 82962 -2248 82996 -2214
rect 82736 -2292 82923 -2258
rect 82736 -2372 82770 -2292
rect 83064 -2372 83098 -2090
rect 82550 -2406 83098 -2372
rect 83148 -2464 83786 -2002
rect 83310 -2478 83328 -2464
rect 83366 -2478 83384 -2464
rect 82550 -2566 83098 -2532
rect 82550 -2848 82584 -2566
rect 82736 -2646 82770 -2566
rect 82912 -2646 82923 -2635
rect 82614 -2686 82686 -2652
rect 82736 -2680 82923 -2646
rect 82614 -2690 82694 -2686
rect 82652 -2724 82694 -2690
rect 82723 -2692 82724 -2691
rect 82724 -2693 82725 -2692
rect 82724 -2722 82725 -2721
rect 82723 -2723 82724 -2722
rect 82668 -2740 82694 -2724
rect 82724 -2742 82730 -2728
rect 82736 -2734 82770 -2680
rect 82924 -2690 82996 -2652
rect 82782 -2692 82783 -2691
rect 82781 -2693 82782 -2692
rect 82781 -2722 82782 -2721
rect 82782 -2723 82783 -2722
rect 82776 -2734 82830 -2728
rect 82912 -2734 82923 -2723
rect 82962 -2724 82996 -2690
rect 82736 -2768 82923 -2734
rect 82736 -2848 82770 -2768
rect 83064 -2848 83098 -2566
rect 82550 -2882 83098 -2848
rect 83148 -2940 83786 -2478
rect 84046 -2668 84048 -1654
rect 84166 -3360 84200 -1618
rect 88468 -1772 88502 -1618
rect 88620 -1694 88622 -1618
rect 88651 -1654 97101 -1618
rect 88651 -1904 89424 -1654
rect 67242 -3988 67362 -3968
rect 67548 -3986 67788 -3434
rect 67548 -3988 67838 -3986
rect 67236 -4016 67390 -3996
rect 67548 -4014 67788 -3988
rect 67548 -4016 67866 -4014
rect 67548 -4072 67788 -4016
rect 88801 -4640 88835 -1904
rect 89425 -3412 89430 -1824
rect 89459 -3412 89464 -1790
rect 89600 -1896 90592 -1654
rect 90117 -4640 90151 -1896
rect 90760 -3492 97101 -1654
rect 97108 -1866 97134 -1578
rect 91169 -4801 91203 -3492
rect 91283 -3924 91328 -3492
rect 91283 -4652 91317 -3924
rect 91340 -4406 91356 -3492
rect 91271 -4699 91330 -4652
rect 91344 -4693 91356 -4406
rect 91433 -3924 91478 -3492
rect 91502 -3564 91714 -3492
rect 91941 -3924 91986 -3492
rect 92002 -3876 92008 -3616
rect 91433 -4640 91467 -3924
rect 91941 -4652 91975 -3924
rect 92058 -4652 92064 -3616
rect 92091 -3924 92136 -3492
rect 92091 -4640 92125 -3924
rect 91405 -4699 91452 -4652
rect 91929 -4699 91988 -4652
rect 92058 -4693 92110 -4652
rect 92063 -4699 92110 -4693
rect 91271 -4733 91452 -4699
rect 91495 -4733 92110 -4699
rect 91271 -4749 91329 -4733
rect 91344 -4746 91356 -4739
rect 91929 -4749 91987 -4733
rect 91271 -4764 91286 -4749
rect 92058 -4801 92064 -4739
rect 92205 -4801 92239 -3492
rect 92388 -3524 92390 -3512
rect 92400 -3572 92402 -3524
rect 88783 -4835 92239 -4801
rect 44808 -6642 44928 -6622
rect 45114 -6640 45354 -6088
rect 45114 -6642 45404 -6640
rect 44802 -6670 44956 -6650
rect 45114 -6668 45354 -6642
rect 45114 -6670 45432 -6668
rect 45114 -6726 45354 -6670
rect 91169 -7393 91203 -4835
rect 92599 -5844 92633 -3492
rect 93037 -5655 93071 -3492
rect 93151 -3768 93196 -3492
rect 93151 -3924 93226 -3768
rect 93151 -5494 93185 -3924
rect 93195 -5124 93226 -3924
rect 93191 -5170 93226 -5124
rect 93251 -5180 93254 -3740
rect 93191 -5198 93254 -5180
rect 93257 -3924 93302 -3492
rect 93257 -5506 93291 -3924
rect 93513 -5506 93547 -3492
rect 93627 -3924 93672 -3492
rect 93627 -5494 93661 -3924
rect 93722 -4676 97101 -3492
rect 97162 -4626 97196 -1062
rect 97230 -1450 97692 -1032
rect 97706 -1450 98168 -1032
rect 98222 -1036 98267 -1032
rect 98222 -1046 98322 -1036
rect 98222 -1062 98267 -1046
rect 98328 -1062 98373 -618
rect 98378 -838 98400 -756
rect 98222 -1318 98256 -1062
rect 97276 -1500 97310 -1450
rect 97276 -1534 97638 -1500
rect 97276 -2014 97322 -1534
rect 97480 -1602 97518 -1564
rect 97446 -1636 97518 -1602
rect 97391 -1686 97436 -1675
rect 97479 -1686 97524 -1675
rect 97402 -1862 97436 -1686
rect 97490 -1862 97524 -1686
rect 97480 -1912 97518 -1874
rect 97446 -1946 97518 -1912
rect 97604 -2014 97638 -1534
rect 97670 -2008 97672 -1466
rect 98108 -1500 98142 -1450
rect 97764 -1534 98142 -1500
rect 97276 -2048 97638 -2014
rect 97764 -2014 97798 -1534
rect 97956 -1602 97994 -1564
rect 97922 -1636 97994 -1602
rect 97867 -1686 97912 -1675
rect 97955 -1686 98000 -1675
rect 97878 -1862 97912 -1686
rect 97966 -1862 98000 -1686
rect 97956 -1912 97994 -1874
rect 97922 -1946 97994 -1912
rect 98080 -2014 98142 -1534
rect 97764 -2048 98142 -2014
rect 97134 -4676 97172 -4638
rect 93722 -4710 97172 -4676
rect 93722 -4778 97101 -4710
rect 97276 -4778 97310 -2048
rect 98108 -3434 98142 -2048
rect 98222 -1630 98262 -1318
rect 98280 -1432 98290 -1374
rect 98278 -1518 98290 -1432
rect 98280 -1574 98290 -1518
rect 98222 -2008 98256 -1630
rect 98316 -1648 98322 -1622
rect 98260 -1678 98262 -1648
rect 98260 -1704 98322 -1678
rect 98328 -2008 98362 -1062
rect 98222 -2226 98267 -2008
rect 98328 -2080 98373 -2008
rect 98328 -2166 98442 -2080
rect 98328 -2226 98373 -2166
rect 98222 -2282 98262 -2226
rect 98222 -3280 98256 -2282
rect 98328 -3280 98362 -2226
rect 98222 -3434 98267 -3280
rect 98328 -3434 98373 -3280
rect 98584 -3434 98618 -618
rect 98698 -1062 98743 -618
rect 97694 -4072 98156 -3434
rect 98170 -4072 98632 -3434
rect 97748 -4156 98098 -4122
rect 97748 -4636 97782 -4156
rect 97940 -4224 97978 -4186
rect 97906 -4258 97978 -4224
rect 97851 -4308 97896 -4297
rect 97939 -4308 97984 -4297
rect 97862 -4484 97896 -4308
rect 97950 -4484 97984 -4308
rect 97940 -4534 97978 -4496
rect 97906 -4568 97978 -4534
rect 98064 -4636 98098 -4156
rect 97748 -4670 98098 -4636
rect 93722 -4812 97310 -4778
rect 93722 -4848 97101 -4812
rect 93809 -5494 93854 -4848
rect 93915 -5506 93960 -4848
rect 94285 -5494 94330 -4848
rect 94467 -5494 94512 -4848
rect 94573 -5506 94618 -4848
rect 93245 -5553 93304 -5506
rect 93513 -5553 93560 -5506
rect 93756 -5553 94619 -5506
rect 94687 -5553 94721 -4848
rect 94943 -5494 94988 -4848
rect 95008 -5180 95036 -4848
rect 95064 -5180 95092 -4848
rect 95125 -5494 95170 -4848
rect 95601 -5494 95646 -4848
rect 95678 -5180 95706 -4848
rect 95734 -5180 95762 -4848
rect 95783 -5494 95828 -4848
rect 96204 -5553 97101 -4848
rect 93213 -5587 97101 -5553
rect 93245 -5603 93303 -5587
rect 93257 -5655 93291 -5621
rect 93513 -5655 93547 -5587
rect 93903 -5603 93961 -5587
rect 94561 -5603 94619 -5587
rect 94573 -5618 94619 -5603
rect 93915 -5655 93949 -5621
rect 94573 -5655 94607 -5618
rect 94687 -5655 94721 -5587
rect 96204 -5655 97101 -5587
rect 93037 -5689 97101 -5655
rect 98108 -5632 98142 -4072
rect 98222 -4122 98256 -4072
rect 98328 -4122 98362 -4072
rect 98222 -4156 98574 -4122
rect 98222 -4200 98267 -4156
rect 98222 -4218 98294 -4200
rect 98222 -4574 98258 -4218
rect 98266 -4300 98294 -4218
rect 98328 -4292 98362 -4156
rect 98416 -4224 98454 -4186
rect 98366 -4258 98454 -4224
rect 98328 -4308 98373 -4292
rect 98415 -4308 98460 -4297
rect 98328 -4484 98372 -4308
rect 98426 -4484 98460 -4308
rect 98266 -4574 98294 -4494
rect 98222 -4636 98294 -4574
rect 98328 -4500 98373 -4484
rect 98328 -4630 98362 -4500
rect 98416 -4534 98454 -4496
rect 98366 -4568 98454 -4534
rect 98540 -4630 98574 -4156
rect 98328 -4636 98373 -4630
rect 98540 -4636 98578 -4630
rect 98222 -4670 98578 -4636
rect 98222 -4848 98294 -4670
rect 98222 -5468 98256 -4848
rect 98266 -5196 98294 -4848
rect 98328 -4848 98373 -4670
rect 98550 -4848 98578 -4670
rect 98222 -5480 98262 -5468
rect 98216 -5492 98262 -5480
rect 98328 -5492 98362 -4848
rect 98584 -5492 98618 -4072
rect 98698 -5480 98732 -1062
rect 98799 -4324 102172 -584
rect 102239 -1062 102284 -584
rect 102308 -590 102618 -584
rect 102308 -694 102610 -590
rect 102308 -918 102520 -694
rect 102239 -4134 102273 -1062
rect 102239 -4324 102284 -4134
rect 102353 -4324 102387 -918
rect 102565 -1062 102610 -694
rect 102682 -1020 102706 -724
rect 102565 -4134 102599 -1062
rect 102565 -4324 102610 -4134
rect 102620 -4324 102632 -4106
rect 102682 -4134 102688 -1020
rect 102648 -4324 102688 -4134
rect 102715 -1062 102760 -584
rect 102715 -4134 102749 -1062
rect 102715 -4324 102760 -4134
rect 102829 -4324 102863 -584
rect 103544 -586 107249 -560
rect 103661 -610 103695 -586
rect 103775 -610 103820 -586
rect 103832 -610 103843 -586
rect 103870 -610 107249 -586
rect 103050 -1230 103472 -610
rect 103526 -1230 107249 -610
rect 103661 -2176 103695 -1230
rect 103737 -1312 103764 -1230
rect 103775 -1372 103822 -1230
rect 103870 -1344 107249 -1230
rect 107310 -1098 107355 746
rect 107310 -1344 107344 -1098
rect 107424 -1344 107458 746
rect 103775 -2176 103809 -1372
rect 103870 -1792 107458 -1344
rect 103870 -2176 107249 -1792
rect 103070 -2202 107249 -2176
rect 103661 -2232 103695 -2202
rect 103775 -2232 103809 -2202
rect 103870 -2232 107249 -2202
rect 103014 -2258 107249 -2232
rect 103154 -3774 103217 -3752
rect 103263 -3774 103290 -3752
rect 103182 -3802 103217 -3780
rect 103263 -3802 103290 -3780
rect 103202 -4324 103276 -4124
rect 98799 -4358 102470 -4324
rect 98799 -4699 102172 -4358
rect 102239 -4392 102273 -4358
rect 102222 -4426 102273 -4392
rect 102294 -4426 102341 -4379
rect 102239 -4460 102341 -4426
rect 102205 -4508 102228 -4503
rect 102183 -4519 102228 -4508
rect 102194 -4699 102228 -4519
rect 102239 -4640 102273 -4460
rect 102353 -4508 102387 -4358
rect 102311 -4519 102387 -4508
rect 102239 -4656 102262 -4640
rect 102322 -4699 102387 -4519
rect 102436 -4652 102470 -4358
rect 102556 -4358 102946 -4324
rect 102556 -4652 102599 -4358
rect 102620 -4512 102632 -4358
rect 102648 -4503 102688 -4358
rect 102715 -4392 102749 -4358
rect 102698 -4426 102749 -4392
rect 102770 -4426 102817 -4379
rect 102715 -4460 102817 -4426
rect 102648 -4512 102704 -4503
rect 102659 -4519 102704 -4512
rect 102670 -4652 102704 -4519
rect 102715 -4640 102749 -4460
rect 102829 -4508 102863 -4358
rect 102787 -4519 102863 -4508
rect 102715 -4652 102738 -4640
rect 102436 -4699 102483 -4652
rect 102553 -4699 102611 -4652
rect 102670 -4656 102738 -4652
rect 102670 -4699 102734 -4656
rect 102798 -4695 102863 -4519
rect 98799 -4733 102734 -4699
rect 98799 -4801 102172 -4733
rect 102294 -4754 102341 -4733
rect 102240 -4788 102341 -4754
rect 102353 -4801 102387 -4733
rect 102436 -4801 102470 -4733
rect 102553 -4749 102611 -4733
rect 102556 -4801 102590 -4749
rect 102682 -4801 102688 -4739
rect 102770 -4754 102817 -4707
rect 102716 -4788 102817 -4754
rect 102829 -4801 102863 -4695
rect 98799 -4835 102863 -4801
rect 98799 -4856 102172 -4835
rect 102436 -4856 102470 -4835
rect 98799 -4871 102470 -4856
rect 98880 -5480 98914 -4871
rect 98986 -5492 99020 -4871
rect 99356 -5480 99390 -4871
rect 99538 -5480 99572 -4871
rect 99644 -5492 99678 -4871
rect 98216 -5524 98244 -5492
rect 98316 -5530 98374 -5492
rect 98584 -5530 98622 -5492
rect 98974 -5530 99032 -5492
rect 99632 -5530 99690 -5492
rect 98284 -5564 99690 -5530
rect 98216 -5626 98244 -5570
rect 98316 -5580 98374 -5564
rect 98328 -5632 98362 -5598
rect 98584 -5632 98618 -5564
rect 98974 -5580 99032 -5564
rect 99632 -5580 99690 -5564
rect 99644 -5595 99690 -5580
rect 99758 -5530 99792 -4871
rect 100014 -5480 100048 -4871
rect 100084 -5180 100112 -4871
rect 100140 -5180 100168 -4871
rect 100196 -5480 100230 -4871
rect 100672 -5480 100706 -4871
rect 100748 -5180 100776 -4871
rect 100804 -5180 100832 -4871
rect 100854 -5480 100888 -4871
rect 101330 -5480 101364 -4871
rect 101400 -5180 101428 -4871
rect 101456 -5180 101484 -4871
rect 101512 -5480 101546 -4871
rect 101626 -5530 101660 -4871
rect 101757 -4890 102470 -4871
rect 102556 -4856 102590 -4835
rect 102912 -4856 102946 -4358
rect 102556 -4890 102946 -4856
rect 103032 -4358 103422 -4324
rect 103032 -4856 103066 -4358
rect 103112 -4512 103130 -4479
rect 103202 -4503 103276 -4358
rect 103202 -4507 103291 -4503
rect 103140 -4508 103158 -4507
rect 103202 -4508 103304 -4507
rect 103135 -4519 103180 -4508
rect 103146 -4695 103180 -4519
rect 103202 -4695 103308 -4508
rect 103202 -4707 103304 -4695
rect 103154 -4708 103180 -4707
rect 103182 -4711 103291 -4707
rect 103182 -4736 103276 -4711
rect 103202 -4764 103276 -4736
rect 103182 -4778 103276 -4764
rect 103182 -4828 103272 -4778
rect 103166 -4842 103182 -4840
rect 103223 -4856 103257 -4828
rect 103388 -4856 103422 -4358
rect 103032 -4890 103422 -4856
rect 101757 -4940 102172 -4890
rect 101757 -5506 102484 -4940
rect 102538 -5506 102960 -4940
rect 103014 -5506 103436 -4940
rect 101757 -5530 103436 -5506
rect 99758 -5553 103436 -5530
rect 103661 -5506 103695 -2258
rect 103775 -5494 103809 -2258
rect 103819 -4778 103850 -3768
rect 103847 -4862 103850 -4778
rect 103870 -4676 107249 -2258
rect 107310 -4626 107344 -1792
rect 107424 -4676 107458 -1792
rect 107636 -1098 107681 746
rect 107762 -1028 107784 188
rect 107636 -3280 107670 -1098
rect 107732 -1392 107758 -1042
rect 107786 -1098 107831 746
rect 107900 -812 107934 746
rect 108260 740 108278 746
rect 108288 712 108334 746
rect 108344 746 112320 780
rect 108344 740 108362 746
rect 108294 -812 108328 712
rect 107732 -1866 107758 -1578
rect 107786 -3280 107820 -1098
rect 107854 -1450 108328 -812
rect 107888 -1500 108100 -1450
rect 107888 -1534 108262 -1500
rect 107888 -1570 108100 -1534
rect 108104 -1570 108142 -1564
rect 107888 -1636 108142 -1570
rect 107888 -1796 108100 -1636
rect 108103 -1686 108148 -1675
rect 107900 -2014 107946 -1796
rect 108026 -1862 108060 -1796
rect 108114 -1862 108148 -1686
rect 108104 -1912 108142 -1874
rect 108070 -1946 108142 -1912
rect 108228 -2014 108262 -1534
rect 107900 -2048 108262 -2014
rect 107598 -3460 107632 -3378
rect 107636 -3502 107681 -3280
rect 107786 -3502 107831 -3280
rect 107900 -3434 107934 -2048
rect 108294 -3434 108328 -1450
rect 108536 -1492 108538 -1404
rect 108732 -3434 108766 746
rect 108834 740 108936 746
rect 108834 708 108892 740
rect 108946 712 112320 746
rect 108846 170 108880 708
rect 108846 -1046 108886 170
rect 108912 -990 108914 114
rect 108947 -462 112320 712
rect 108947 -910 112348 -462
rect 108846 -3280 108880 -1046
rect 108884 -1448 108886 -1392
rect 108884 -1704 108886 -1648
rect 108884 -1848 108886 -1792
rect 108884 -2104 108886 -2048
rect 108846 -3434 108891 -3280
rect 108947 -3434 112320 -910
rect 107636 -4630 107670 -3502
rect 107786 -3940 107820 -3502
rect 107762 -3996 107820 -3940
rect 107786 -4140 107820 -3996
rect 107842 -4072 108780 -3434
rect 108794 -4072 112320 -3434
rect 107900 -4122 107934 -4072
rect 108196 -4122 108210 -4072
rect 107762 -4252 107820 -4140
rect 107786 -4626 107820 -4252
rect 107896 -4156 108246 -4122
rect 107636 -4638 107681 -4630
rect 107896 -4636 107934 -4156
rect 108088 -4224 108126 -4186
rect 108054 -4258 108126 -4224
rect 107999 -4308 108044 -4297
rect 108087 -4308 108132 -4297
rect 108196 -4300 108210 -4156
rect 108010 -4484 108044 -4308
rect 108098 -4484 108132 -4308
rect 108088 -4534 108126 -4496
rect 108054 -4568 108126 -4534
rect 108212 -4636 108246 -4156
rect 107512 -4676 107796 -4638
rect 107896 -4670 108246 -4636
rect 103870 -4710 107796 -4676
rect 103870 -4778 107249 -4710
rect 107424 -4778 107458 -4710
rect 107568 -4726 107682 -4710
rect 107568 -4778 107670 -4726
rect 107900 -4778 107934 -4670
rect 103870 -4812 107934 -4778
rect 103870 -4848 107249 -4812
rect 103875 -4862 103878 -4848
rect 103847 -5124 103850 -5062
rect 103815 -5170 103850 -5124
rect 103875 -5180 103878 -5062
rect 103815 -5198 103878 -5180
rect 103881 -5506 103926 -4848
rect 104433 -5494 104478 -4848
rect 104539 -5506 104584 -4848
rect 104610 -5506 104611 -5302
rect 105048 -5506 105052 -5302
rect 105086 -5506 105090 -5302
rect 105091 -5494 105136 -4848
rect 105191 -5180 105242 -4848
rect 105197 -5506 105242 -5180
rect 103661 -5553 103708 -5506
rect 103868 -5553 105243 -5506
rect 105311 -5553 105345 -4848
rect 106828 -5492 107249 -4848
rect 107636 -5124 107670 -4812
rect 107630 -5408 107670 -5124
rect 107636 -5492 107670 -5408
rect 108294 -5492 108328 -4072
rect 108372 -4156 108722 -4122
rect 108372 -4636 108406 -4156
rect 108564 -4224 108602 -4186
rect 108530 -4258 108602 -4224
rect 108475 -4308 108520 -4297
rect 108563 -4308 108608 -4297
rect 108486 -4484 108520 -4308
rect 108574 -4484 108608 -4308
rect 108564 -4534 108602 -4496
rect 108530 -4568 108602 -4534
rect 108688 -4636 108722 -4156
rect 108372 -4670 108722 -4636
rect 106828 -5530 107948 -5492
rect 108266 -5496 108328 -5492
rect 108732 -5492 108766 -4072
rect 108846 -4122 108880 -4072
rect 108947 -4122 112320 -4072
rect 108846 -4156 112320 -4122
rect 108846 -4200 108891 -4156
rect 108947 -4200 112320 -4156
rect 108846 -4218 108918 -4200
rect 108846 -4574 108882 -4218
rect 108890 -4300 108918 -4218
rect 108946 -4300 112320 -4200
rect 108890 -4574 108918 -4494
rect 108846 -4636 108918 -4574
rect 108947 -4636 112320 -4300
rect 108846 -4670 112320 -4636
rect 112387 -4134 112421 3336
rect 112501 3042 112535 3395
rect 113913 3361 113940 3463
rect 113941 3389 113968 3435
rect 112501 1690 112538 3042
rect 112387 -4356 112432 -4134
rect 112387 -4640 112421 -4356
rect 108846 -4802 108918 -4670
rect 108947 -4699 112320 -4670
rect 112501 -4699 112535 1690
rect 113212 -28 113602 6
rect 113212 -526 113246 -28
rect 113426 -96 113473 -49
rect 113388 -130 113473 -96
rect 113315 -189 113360 -178
rect 113443 -189 113488 -178
rect 113326 -365 113360 -189
rect 113454 -365 113488 -189
rect 113426 -424 113473 -377
rect 113388 -458 113473 -424
rect 113446 -462 113452 -458
rect 113458 -498 113464 -462
rect 113568 -526 113602 -28
rect 113212 -560 113602 -526
rect 113198 -1230 113620 -610
rect 113891 -1226 113925 3336
rect 113968 1696 113970 3048
rect 113968 -378 113986 196
rect 114018 -504 115391 3497
rect 116874 3434 116908 3481
rect 117572 3450 117583 3461
rect 117595 3450 117606 3461
rect 117572 3434 117606 3450
rect 116874 3400 117606 3434
rect 116058 2392 116194 2502
rect 116058 2366 116210 2392
rect 116118 1934 116210 2366
rect 115996 -496 116458 42
rect 114018 -760 115400 -504
rect 115414 -732 115456 -532
rect 115996 -562 116606 -496
rect 115996 -596 116668 -562
rect 116116 -646 116142 -612
rect 116394 -638 116668 -596
rect 116394 -646 116606 -638
rect 116054 -680 116606 -646
rect 113826 -1312 113925 -1226
rect 113776 -2176 113802 -1372
rect 113804 -2176 113830 -1372
rect 113891 -2176 113925 -1312
rect 113968 -1372 113970 -824
rect 114018 -2176 115391 -760
rect 116054 -1160 116088 -680
rect 116142 -786 116176 -680
rect 116246 -748 116284 -710
rect 116196 -782 116210 -748
rect 116212 -782 116284 -748
rect 116142 -818 116182 -786
rect 116192 -790 116210 -786
rect 116246 -790 116268 -786
rect 116274 -818 116296 -786
rect 116142 -832 116176 -818
rect 116188 -832 116202 -821
rect 116245 -832 116290 -821
rect 116142 -1008 116202 -832
rect 116256 -1008 116290 -832
rect 116370 -944 116606 -680
rect 116766 -720 116770 -520
rect 116794 -748 116798 -492
rect 116142 -1022 116176 -1008
rect 116246 -1022 116284 -1020
rect 116142 -1126 116182 -1022
rect 116196 -1108 116210 -1050
rect 116246 -1058 116290 -1022
rect 116212 -1092 116290 -1058
rect 116246 -1108 116262 -1092
rect 116116 -1136 116182 -1126
rect 116274 -1136 116290 -1092
rect 116116 -1160 116176 -1136
rect 116370 -1160 116404 -944
rect 116054 -1194 116404 -1160
rect 116766 -1372 116790 -824
rect 116794 -1120 116818 -796
rect 116794 -1400 116822 -1120
rect 116800 -1406 116822 -1400
rect 116246 -2174 116248 -1974
rect 113218 -2202 115391 -2176
rect 116274 -2202 116276 -1946
rect 113212 -3600 113286 -3270
rect 113212 -3754 113418 -3600
rect 113212 -3924 113286 -3754
rect 113242 -4324 113267 -4290
rect 108947 -4733 112535 -4699
rect 108947 -4801 112320 -4733
rect 112501 -4749 112535 -4733
rect 112501 -4760 112512 -4749
rect 112524 -4760 112535 -4749
rect 112704 -4358 113094 -4324
rect 112704 -4749 112738 -4358
rect 112918 -4426 112965 -4379
rect 112880 -4460 112965 -4426
rect 112807 -4519 112852 -4508
rect 112935 -4519 112980 -4508
rect 112818 -4652 112852 -4519
rect 112946 -4652 112980 -4519
rect 112806 -4699 112864 -4652
rect 112934 -4699 112992 -4652
rect 112780 -4707 113018 -4699
rect 112780 -4716 112890 -4707
rect 112908 -4716 113018 -4707
rect 112780 -4733 113018 -4716
rect 112704 -4760 112715 -4749
rect 112727 -4760 112738 -4749
rect 113060 -4749 113094 -4358
rect 113180 -4358 113570 -4324
rect 113180 -4665 113214 -4358
rect 113233 -4656 113248 -4358
rect 113394 -4426 113441 -4379
rect 113356 -4460 113441 -4426
rect 113260 -4479 113267 -4469
rect 113260 -4481 113273 -4479
rect 113256 -4512 113273 -4481
rect 113294 -4507 113301 -4503
rect 113288 -4508 113301 -4507
rect 113326 -4508 113334 -4507
rect 113256 -4640 113267 -4512
rect 113283 -4519 113334 -4508
rect 113260 -4656 113267 -4640
rect 113294 -4652 113334 -4519
rect 113180 -4733 113239 -4665
rect 113282 -4699 113340 -4652
rect 113354 -4693 113362 -4479
rect 113411 -4519 113456 -4508
rect 113422 -4652 113456 -4519
rect 113410 -4699 113468 -4652
rect 113282 -4707 113494 -4699
rect 113295 -4716 113366 -4707
rect 113384 -4716 113494 -4707
rect 113295 -4718 113494 -4716
rect 113286 -4733 113494 -4718
rect 112704 -4794 112738 -4767
rect 112864 -4788 112934 -4754
rect 113060 -4760 113071 -4749
rect 113083 -4760 113094 -4749
rect 113126 -4762 113140 -4739
rect 113060 -4794 113094 -4767
rect 113154 -4790 113168 -4739
rect 113180 -4749 113214 -4733
rect 113286 -4739 113354 -4733
rect 113180 -4760 113191 -4749
rect 113203 -4760 113214 -4749
rect 113314 -4754 113354 -4746
rect 113536 -4749 113570 -4358
rect 113776 -4693 113802 -2202
rect 113804 -4693 113830 -2202
rect 113891 -4640 113925 -2202
rect 113776 -4746 113802 -4739
rect 113314 -4767 113410 -4754
rect 113536 -4760 113547 -4749
rect 113559 -4760 113570 -4749
rect 113180 -4794 113214 -4767
rect 113340 -4788 113410 -4767
rect 113536 -4794 113570 -4767
rect 113804 -4774 113830 -4739
rect 114018 -4778 115391 -2202
rect 115442 -4336 115456 -2934
rect 116246 -3774 116258 -3574
rect 116274 -3802 116286 -3546
rect 116736 -4400 116762 -2942
rect 116764 -4372 116790 -2970
rect 116870 -4372 116872 -2970
rect 116874 -4676 116908 3400
rect 116977 3350 117022 3361
rect 117447 3350 117492 3361
rect 116988 -4626 117022 3350
rect 117232 -508 117444 -490
rect 117038 -938 117444 -508
rect 117038 -956 117250 -938
rect 117458 -4626 117492 3350
rect 117572 2786 117606 3400
rect 117572 1682 117624 2786
rect 163643 2229 163677 7372
rect 165511 3967 165545 10465
rect 165987 10444 166021 10465
rect 166101 10462 166146 10465
rect 166101 10444 166135 10462
rect 165625 10428 165672 10444
rect 165613 10397 165672 10428
rect 165703 10403 165750 10444
rect 165686 10397 165750 10403
rect 165987 10397 166034 10444
rect 166101 10397 166148 10444
rect 166162 10416 166190 10465
rect 166283 10462 166328 10465
rect 166759 10462 166804 10465
rect 166283 10444 166317 10462
rect 166759 10444 166793 10462
rect 166283 10397 166330 10444
rect 166361 10397 166408 10444
rect 166759 10397 166806 10444
rect 166820 10416 166848 10465
rect 166876 10416 166904 10465
rect 166941 10462 166986 10465
rect 166941 10444 166975 10462
rect 166941 10397 166988 10444
rect 167019 10397 167066 10444
rect 165613 10363 165750 10397
rect 165793 10363 166408 10397
rect 166451 10363 167066 10397
rect 165613 10357 165715 10363
rect 165613 10316 165671 10357
rect 165742 10329 165743 10363
rect 165625 10072 165659 10316
rect 165720 10304 165765 10315
rect 165625 8608 165665 10072
rect 165682 8664 165693 10016
rect 165625 4128 165659 8608
rect 165669 4452 165700 5854
rect 165725 4424 165728 5882
rect 165731 4116 165765 10304
rect 165987 4116 166021 10363
rect 166101 4128 166135 10363
rect 166283 4128 166317 10363
rect 166378 10304 166423 10315
rect 166389 8306 166423 10304
rect 166320 8298 166532 8306
rect 166320 7858 166732 8298
rect 166389 4116 166423 7858
rect 166520 7850 166732 7858
rect 166759 4128 166793 10363
rect 166941 4128 166975 10363
rect 167036 10304 167081 10315
rect 167047 8298 167081 10304
rect 167161 8306 167195 10465
rect 167383 10462 167398 11568
rect 167161 8298 167378 8306
rect 166996 7858 167378 8298
rect 166996 7850 167208 7858
rect 167047 4116 167081 7850
rect 165719 4069 165778 4116
rect 165987 4069 166034 4116
rect 166377 4069 166436 4116
rect 167035 4069 167093 4116
rect 165687 4035 167093 4069
rect 165619 3973 165642 4029
rect 165719 4019 165777 4035
rect 165731 3967 165765 4001
rect 165987 3967 166021 4035
rect 166324 4022 166435 4035
rect 166377 4020 166435 4022
rect 166352 4019 166435 4020
rect 167035 4019 167093 4035
rect 166352 3967 166383 4019
rect 167078 4004 167093 4019
rect 167161 4069 167195 7850
rect 167417 4128 167451 12104
rect 167482 6430 167510 11780
rect 167538 6430 167566 11780
rect 167482 4075 167510 6244
rect 167538 4075 167566 6244
rect 167599 4128 167633 12104
rect 167850 8298 167854 8306
rect 167862 7858 167866 8298
rect 168075 7164 168109 12104
rect 168075 6974 168120 7164
rect 168152 6974 168180 11780
rect 168208 6974 168236 11780
rect 168257 7164 168291 12104
rect 168733 10540 168767 12104
rect 168860 10540 168888 11780
rect 168915 10540 168949 12104
rect 169029 10540 169063 12163
rect 168678 10504 169575 10540
rect 170582 10504 170616 12208
rect 171058 12202 171092 12249
rect 172558 12208 172586 12228
rect 172614 12208 172642 12240
rect 173222 12208 173250 12228
rect 173278 12208 173306 12228
rect 173930 12208 173958 12228
rect 174100 12218 174111 12229
rect 174123 12218 174134 12229
rect 174100 12202 174134 12218
rect 171058 12168 174134 12202
rect 171058 10504 171092 12168
rect 171161 12118 171206 12129
rect 171343 12118 171388 12129
rect 171819 12118 171864 12129
rect 172001 12118 172046 12129
rect 172477 12118 172522 12129
rect 171172 10504 171206 12118
rect 171248 10504 171276 11780
rect 171354 10504 171388 12118
rect 171830 10504 171864 12118
rect 171900 10504 171928 11780
rect 171956 10504 171984 11780
rect 172012 10504 172046 12118
rect 168678 10470 172266 10504
rect 168678 8298 169575 10470
rect 170582 8810 170616 10470
rect 171058 10440 171092 10470
rect 171172 10440 171206 10470
rect 170696 10433 170734 10440
rect 170684 10418 170734 10433
rect 170774 10436 170812 10440
rect 170684 10402 170742 10418
rect 170774 10408 170814 10436
rect 170750 10402 170814 10408
rect 171058 10402 171096 10440
rect 171172 10402 171210 10440
rect 171248 10428 171276 10470
rect 171354 10440 171388 10470
rect 171830 10440 171864 10470
rect 171354 10402 171392 10440
rect 171432 10402 171470 10440
rect 171830 10402 171868 10440
rect 171900 10434 171928 10470
rect 171956 10434 171984 10470
rect 172012 10440 172046 10470
rect 172012 10402 172050 10440
rect 172090 10402 172128 10440
rect 170684 10368 170814 10402
rect 170864 10368 171470 10402
rect 171522 10368 172128 10402
rect 170684 10362 170786 10368
rect 170684 10330 170742 10362
rect 170806 10334 170814 10368
rect 170696 9792 170730 10330
rect 170791 10318 170836 10329
rect 170696 8964 170736 9792
rect 168338 7850 169575 8298
rect 169704 8172 170166 8810
rect 170180 8172 170642 8810
rect 170696 8742 170741 8964
rect 170696 8586 170736 8742
rect 170762 8642 170764 9736
rect 170802 8964 170836 10318
rect 170802 8742 170847 8964
rect 170852 8784 170874 8866
rect 170762 8632 170796 8642
rect 170696 8576 170796 8586
rect 170696 8304 170730 8576
rect 168257 6974 168302 7164
rect 167872 6942 168302 6974
rect 167872 6940 168291 6942
rect 167872 6442 167906 6940
rect 168075 6919 168109 6940
rect 168075 6872 168122 6919
rect 168048 6838 168122 6872
rect 168075 6790 168109 6838
rect 168114 6790 168143 6795
rect 167975 6779 168020 6790
rect 167986 6603 168020 6779
rect 168075 6779 168148 6790
rect 168152 6786 168180 6940
rect 168208 6786 168291 6940
rect 168075 6591 168109 6779
rect 168114 6603 168148 6779
rect 168114 6591 168143 6603
rect 168075 6587 168143 6591
rect 168228 6590 168291 6786
rect 168075 6544 168122 6587
rect 168048 6510 168122 6544
rect 168075 6442 168109 6510
rect 168152 6442 168180 6590
rect 168208 6442 168291 6590
rect 167872 6408 168291 6442
rect 168075 6358 168109 6408
rect 168152 6358 168180 6408
rect 168208 6358 168236 6408
rect 168257 6358 168291 6408
rect 167858 5814 168291 6358
rect 167858 5738 168302 5814
rect 168075 5596 168120 5738
rect 168075 4128 168109 5596
rect 168152 4075 168180 5738
rect 168208 4075 168236 5738
rect 168257 5596 168302 5738
rect 168257 4128 168291 5596
rect 168678 4069 169575 7850
rect 169762 8088 170112 8122
rect 169762 7608 169796 8088
rect 169954 8020 169992 8058
rect 169920 7986 169992 8020
rect 169865 7936 169910 7947
rect 169953 7936 169998 7947
rect 169876 7760 169910 7936
rect 169964 7760 169998 7936
rect 169954 7710 169992 7748
rect 169920 7676 169992 7710
rect 170078 7608 170112 8088
rect 170144 7614 170146 8156
rect 170582 8122 170616 8172
rect 170238 8088 170616 8122
rect 169762 7574 170112 7608
rect 170238 7608 170272 8088
rect 170430 8020 170468 8058
rect 170396 7986 170468 8020
rect 170341 7936 170386 7947
rect 170429 7936 170474 7947
rect 170352 7760 170386 7936
rect 170440 7760 170474 7936
rect 170430 7710 170468 7748
rect 170396 7676 170468 7710
rect 170554 7608 170616 8088
rect 170238 7574 170616 7608
rect 167161 4035 169575 4069
rect 166389 3967 166423 4001
rect 167047 3967 167081 4001
rect 167161 3967 167195 4035
rect 167482 4022 167510 4029
rect 167538 4022 167566 4029
rect 168152 4022 168180 4029
rect 168208 4022 168236 4029
rect 168678 3967 169575 4035
rect 165511 3933 169575 3967
rect 170582 3990 170616 7574
rect 170696 7992 170736 8304
rect 170754 8190 170764 8248
rect 170752 8104 170764 8190
rect 170754 8048 170764 8104
rect 170696 7614 170730 7992
rect 170790 7974 170796 8000
rect 170734 7944 170736 7974
rect 170734 7918 170796 7944
rect 170802 7614 170836 8742
rect 170696 7396 170741 7614
rect 170802 7542 170847 7614
rect 170802 7456 170916 7542
rect 170802 7396 170847 7456
rect 170696 7340 170736 7396
rect 170696 4142 170730 7340
rect 170740 4426 170768 5828
rect 170802 4130 170836 7396
rect 171058 4130 171092 10368
rect 171172 4142 171206 10368
rect 171354 4142 171388 10368
rect 171449 10318 171494 10329
rect 171460 8278 171494 10318
rect 171416 8274 171628 8278
rect 171416 7830 171818 8274
rect 171460 4130 171494 7830
rect 171606 7826 171818 7830
rect 171830 4142 171864 10368
rect 172012 4142 172046 10368
rect 172107 10318 172152 10329
rect 172118 8274 172152 10318
rect 172232 8278 172266 10470
rect 172232 8274 172466 8278
rect 172082 7830 172466 8274
rect 172082 7826 172294 7830
rect 172118 4130 172152 7826
rect 170790 4092 170848 4130
rect 171058 4092 171096 4130
rect 171448 4092 171506 4130
rect 172106 4098 172164 4130
rect 172034 4092 172164 4098
rect 172232 4092 172266 7826
rect 172488 4142 172522 12118
rect 172558 4098 172586 12162
rect 172614 4142 172642 12162
rect 172659 12118 172704 12129
rect 173135 12118 173180 12129
rect 172670 4142 172704 12118
rect 172730 8272 172942 8278
rect 172730 7830 173134 8272
rect 172922 7824 173134 7830
rect 173146 4142 173180 12118
rect 173222 4098 173250 12162
rect 173278 4098 173306 12162
rect 173317 12118 173362 12129
rect 173793 12118 173838 12129
rect 173328 4142 173362 12118
rect 173398 8260 173610 8272
rect 173398 7824 173778 8260
rect 173566 7812 173778 7824
rect 173804 4142 173838 12118
rect 173874 10378 173902 11594
rect 173874 4218 173902 5910
rect 173930 4098 173958 12162
rect 173975 12118 174020 12129
rect 173986 4142 174020 12118
rect 174100 4092 174134 12168
rect 174231 10499 174646 12265
rect 176135 12197 176169 12235
rect 177785 12213 177796 12224
rect 177808 12213 177819 12224
rect 177785 12197 177819 12213
rect 175759 12163 178195 12197
rect 174996 10499 175002 11594
rect 175039 10499 175073 10533
rect 175697 10499 175731 10533
rect 176135 10499 176169 12163
rect 176238 12104 176294 12115
rect 176344 12104 176400 12115
rect 176896 12104 176952 12115
rect 177002 12104 177058 12115
rect 177554 12104 177610 12115
rect 177660 12104 177716 12115
rect 176249 10499 176294 12104
rect 176306 10499 176317 11780
rect 176355 10499 176400 12104
rect 176907 10499 176952 12104
rect 177013 11780 177058 12104
rect 176979 10499 176992 11780
rect 177007 10499 177058 11780
rect 177565 10499 177610 12104
rect 177628 10499 177633 11780
rect 177671 10499 177716 12104
rect 177785 10499 177819 12163
rect 174231 10465 177819 10499
rect 174231 10397 174646 10465
rect 174996 10458 175002 10465
rect 175039 10444 175073 10465
rect 175697 10444 175731 10465
rect 175011 10431 175073 10444
rect 175669 10431 175731 10444
rect 175011 10403 175079 10431
rect 175669 10403 175737 10431
rect 175005 10397 175079 10403
rect 175089 10397 175107 10403
rect 175663 10397 175737 10403
rect 175747 10397 175765 10403
rect 176135 10397 176169 10465
rect 176249 10462 176294 10465
rect 176306 10464 176317 10465
rect 176355 10462 176400 10465
rect 176907 10462 176952 10465
rect 176249 10444 176289 10462
rect 176355 10444 176389 10462
rect 176249 10413 176296 10444
rect 176237 10403 176296 10413
rect 176327 10403 176389 10444
rect 176907 10444 176941 10462
rect 176979 10458 176992 10465
rect 177007 10462 177058 10465
rect 177565 10462 177610 10465
rect 177007 10444 177048 10462
rect 176907 10413 176954 10444
rect 176237 10402 176389 10403
rect 176237 10397 176296 10402
rect 176321 10397 176389 10402
rect 176895 10403 176954 10413
rect 176985 10403 177048 10444
rect 177565 10444 177599 10462
rect 177600 10444 177605 10462
rect 177565 10413 177612 10444
rect 177628 10434 177633 10465
rect 177671 10462 177716 10465
rect 177671 10444 177705 10462
rect 176895 10402 177048 10403
rect 176895 10397 176954 10402
rect 176979 10397 177047 10402
rect 177553 10397 177612 10413
rect 177643 10403 177705 10444
rect 177637 10397 177705 10403
rect 174231 10363 175079 10397
rect 175085 10363 175737 10397
rect 175743 10363 176389 10397
rect 176401 10363 177047 10397
rect 177059 10363 177705 10397
rect 174231 5298 174646 10363
rect 175005 10357 175023 10363
rect 175033 10329 175079 10363
rect 175089 10357 175107 10363
rect 175663 10357 175681 10363
rect 175691 10329 175737 10363
rect 175747 10357 175765 10363
rect 175039 5298 175073 10329
rect 175697 5498 175731 10329
rect 175676 5298 175750 5498
rect 174231 5264 174944 5298
rect 174231 4766 174646 5264
rect 174768 5196 174815 5243
rect 174730 5162 174815 5196
rect 174657 5103 174702 5114
rect 174785 5103 174830 5114
rect 174668 4927 174702 5103
rect 174796 4927 174830 5103
rect 174768 4868 174815 4915
rect 174730 4834 174815 4868
rect 174910 4766 174944 5264
rect 174231 4732 174944 4766
rect 175030 5264 175420 5298
rect 175030 5202 175073 5264
rect 175030 4766 175064 5202
rect 175244 5196 175291 5243
rect 175206 5162 175291 5196
rect 175133 5103 175178 5114
rect 175261 5103 175306 5114
rect 175144 4927 175178 5103
rect 175272 4927 175306 5103
rect 175244 4868 175291 4915
rect 175206 4834 175291 4868
rect 175386 4766 175420 5264
rect 175030 4732 175420 4766
rect 175506 5264 175896 5298
rect 175506 4766 175540 5264
rect 175586 5110 175604 5143
rect 175676 5119 175750 5264
rect 175676 5115 175765 5119
rect 175614 5114 175632 5115
rect 175676 5114 175778 5115
rect 175609 5103 175654 5114
rect 175620 4927 175654 5103
rect 175676 4927 175782 5114
rect 175676 4915 175778 4927
rect 175628 4914 175654 4915
rect 175656 4911 175765 4915
rect 175656 4886 175750 4911
rect 175676 4858 175750 4886
rect 175656 4844 175750 4858
rect 175656 4794 175746 4844
rect 175640 4780 175656 4782
rect 175697 4766 175731 4794
rect 175862 4766 175896 5264
rect 175506 4732 175896 4766
rect 174231 4682 174646 4732
rect 174231 4116 174958 4682
rect 175012 4116 175434 4682
rect 175488 4116 175910 4682
rect 174231 4092 175910 4116
rect 170758 4069 175910 4092
rect 176135 4116 176169 10363
rect 176237 10316 176295 10363
rect 176321 10357 176339 10363
rect 176349 10329 176389 10363
rect 176249 10072 176283 10316
rect 176249 8608 176289 10072
rect 176306 8664 176317 10016
rect 176249 4128 176283 8608
rect 176321 4760 176324 5854
rect 176349 4760 176352 5882
rect 176321 4452 176324 4560
rect 176349 4424 176352 4560
rect 176355 4116 176389 10329
rect 176895 10316 176953 10363
rect 176979 10357 176997 10363
rect 177007 10329 177047 10363
rect 176468 8298 176680 8306
rect 176468 7858 176830 8298
rect 176618 7850 176830 7858
rect 176907 5876 176941 10316
rect 176907 4362 176947 5876
rect 176907 4128 176941 4362
rect 177013 4116 177047 10329
rect 177553 10316 177611 10363
rect 177637 10357 177655 10363
rect 177665 10329 177705 10363
rect 177144 7850 177476 8298
rect 177565 4128 177599 10316
rect 177600 8606 177605 10014
rect 177628 8634 177633 9986
rect 177671 5898 177705 10329
rect 177665 4384 177705 5898
rect 177671 4116 177705 4384
rect 177785 8306 177819 10465
rect 179302 10504 179723 12265
rect 181206 12202 181240 12249
rect 182856 12218 182867 12229
rect 182879 12218 182890 12229
rect 182856 12202 182890 12218
rect 181206 12168 182890 12202
rect 180110 10504 180144 10538
rect 180768 10504 180802 10538
rect 181206 10504 181240 12168
rect 181309 12118 181354 12129
rect 181415 12118 181460 12129
rect 181967 12118 182012 12129
rect 182073 12118 182118 12129
rect 182625 12118 182670 12129
rect 182731 12118 182776 12129
rect 181320 11592 181354 12118
rect 181320 10504 181360 11592
rect 181386 10504 181388 11536
rect 181426 10504 181460 12118
rect 181978 10504 182012 12118
rect 182084 11610 182118 12118
rect 182050 10504 182070 11554
rect 182078 10504 182126 11610
rect 182636 11566 182670 12118
rect 182636 10504 182676 11566
rect 182694 10504 182704 11538
rect 182742 10504 182776 12118
rect 182856 10504 182890 12168
rect 179302 10470 182890 10504
rect 179302 10402 179723 10470
rect 180110 10440 180144 10470
rect 180768 10440 180802 10470
rect 180082 10436 180144 10440
rect 180740 10436 180802 10440
rect 180082 10408 180150 10436
rect 180740 10408 180808 10436
rect 180076 10402 180150 10408
rect 180160 10402 180178 10408
rect 180734 10402 180808 10408
rect 180818 10402 180836 10408
rect 181206 10402 181240 10470
rect 181320 10418 181360 10470
rect 181386 10436 181388 10470
rect 181426 10440 181460 10470
rect 181398 10436 181460 10440
rect 181386 10432 181460 10436
rect 181308 10408 181366 10418
rect 181398 10408 181460 10432
rect 181978 10440 182012 10470
rect 182050 10450 182070 10470
rect 182078 10440 182126 10470
rect 181978 10418 182016 10440
rect 181308 10402 181460 10408
rect 181966 10408 182024 10418
rect 182056 10408 182126 10440
rect 182636 10418 182676 10470
rect 182694 10436 182704 10470
rect 182742 10440 182776 10470
rect 182714 10436 182776 10440
rect 182694 10434 182776 10436
rect 181966 10402 182126 10408
rect 182624 10408 182682 10418
rect 182714 10408 182776 10434
rect 182624 10406 182776 10408
rect 182624 10402 182682 10406
rect 182708 10402 182776 10406
rect 179302 10368 180150 10402
rect 180156 10368 180808 10402
rect 180814 10368 181460 10402
rect 181472 10368 182118 10402
rect 182130 10368 182776 10402
rect 178496 8740 178886 8774
rect 177785 8206 178002 8306
rect 178496 8298 178530 8740
rect 178710 8672 178757 8719
rect 178672 8638 178757 8672
rect 178599 8579 178644 8590
rect 178727 8579 178772 8590
rect 178610 8403 178644 8579
rect 178738 8403 178772 8579
rect 178710 8344 178757 8391
rect 178672 8334 178757 8344
rect 178646 8310 178757 8334
rect 178646 8298 178736 8310
rect 178486 8270 178736 8298
rect 178486 8242 178698 8270
rect 178852 8242 178886 8740
rect 179302 8298 179723 10368
rect 180076 10362 180094 10368
rect 180104 10334 180150 10368
rect 180160 10362 180178 10368
rect 180734 10362 180752 10368
rect 180762 10334 180808 10368
rect 180818 10362 180836 10368
rect 178486 8208 178886 8242
rect 179132 8278 179723 8298
rect 177785 8074 178038 8206
rect 178486 8158 178698 8208
rect 179132 8206 179908 8278
rect 177785 7858 178002 8074
rect 176135 4069 176182 4116
rect 176343 4069 176402 4116
rect 177001 4069 177060 4116
rect 177659 4069 177717 4116
rect 170758 4062 177717 4069
rect 170758 4058 175079 4062
rect 170690 3996 170718 4052
rect 170790 4042 170848 4058
rect 170802 3990 170836 4024
rect 171058 3990 171092 4058
rect 171448 4042 171506 4058
rect 172106 4042 172164 4058
rect 172118 4027 172164 4042
rect 171424 3990 171454 3998
rect 171460 3990 171494 4024
rect 171500 3990 171532 3998
rect 172118 3990 172152 4027
rect 172232 3990 172266 4058
rect 172558 4046 172586 4052
rect 173222 4040 173250 4052
rect 173278 4046 173306 4052
rect 173930 4040 173958 4052
rect 174100 4042 174134 4058
rect 174100 4031 174111 4042
rect 174123 4031 174134 4042
rect 174231 4035 175079 4058
rect 174231 3990 174646 4035
rect 175005 4029 175023 4035
rect 175033 4001 175079 4035
rect 175089 4035 175716 4062
rect 175719 4057 175737 4062
rect 175747 4057 177717 4062
rect 175719 4042 177717 4057
rect 175089 4029 175107 4035
rect 170582 3967 174646 3990
rect 175039 3967 175073 4001
rect 175697 3997 175707 4035
rect 175721 3997 175731 4042
rect 175759 4035 177717 4042
rect 176135 3967 176169 4035
rect 176343 4019 176401 4035
rect 176948 4029 177059 4035
rect 177001 4020 177059 4029
rect 176976 4019 177059 4020
rect 177659 4019 177717 4035
rect 176976 4001 177007 4019
rect 177702 4004 177717 4019
rect 177785 3967 177819 7858
rect 178482 7538 178904 8158
rect 179060 8130 179908 8206
rect 179132 7850 179908 8130
rect 179302 7830 179908 7850
rect 178496 6940 178886 6974
rect 178496 6442 178530 6940
rect 178710 6872 178757 6919
rect 178672 6838 178757 6872
rect 178852 6912 178886 6940
rect 178599 6779 178644 6790
rect 178727 6779 178772 6790
rect 178610 6603 178644 6779
rect 178738 6603 178772 6779
rect 178710 6582 178757 6591
rect 178580 6566 178658 6582
rect 178710 6566 178790 6582
rect 178710 6554 178757 6566
rect 178608 6538 178658 6554
rect 178710 6544 178762 6554
rect 178672 6538 178762 6544
rect 178672 6510 178757 6538
rect 178852 6504 178920 6912
rect 178852 6442 178886 6504
rect 178496 6408 178886 6442
rect 178482 5738 178904 6358
rect 179302 4092 179723 7830
rect 180110 4130 180144 10334
rect 180768 8810 180802 10334
rect 180328 8172 180802 8810
rect 180362 8122 180574 8172
rect 180362 8088 180736 8122
rect 180362 8052 180574 8088
rect 180578 8052 180616 8058
rect 180362 7986 180616 8052
rect 180362 7826 180574 7986
rect 180577 7936 180622 7947
rect 180386 7608 180420 7826
rect 180500 7760 180534 7826
rect 180588 7760 180622 7936
rect 180578 7710 180616 7748
rect 180544 7676 180616 7710
rect 180702 7608 180736 8088
rect 180386 7574 180736 7608
rect 180768 4130 180802 8172
rect 181010 8130 181012 8218
rect 180082 4126 180144 4130
rect 180740 4126 180802 4130
rect 181206 4130 181240 10368
rect 181308 10330 181366 10368
rect 181392 10362 181410 10368
rect 181420 10334 181460 10368
rect 181320 9792 181354 10330
rect 181320 8576 181360 9792
rect 181386 8632 181388 9736
rect 181320 4142 181354 8576
rect 181426 4130 181460 10334
rect 181966 10330 182024 10368
rect 182050 10362 182068 10368
rect 182078 10334 182118 10368
rect 181564 8272 181776 8278
rect 181564 7830 181890 8272
rect 181678 7824 181890 7830
rect 181978 5854 182012 10330
rect 181978 4340 182018 5854
rect 181978 4142 182012 4340
rect 182084 4130 182118 10334
rect 182624 10330 182682 10368
rect 182708 10362 182726 10368
rect 182736 10334 182776 10368
rect 182636 9766 182670 10330
rect 182636 8606 182676 9766
rect 182694 8634 182704 9738
rect 182230 8260 182442 8274
rect 182230 7826 182534 8260
rect 182322 7812 182534 7826
rect 182636 4142 182670 8606
rect 182742 5890 182776 10334
rect 182736 4376 182776 5890
rect 182742 4130 182776 4376
rect 180082 4098 180150 4126
rect 180740 4098 180808 4126
rect 180076 4092 180150 4098
rect 180160 4092 180178 4098
rect 180734 4092 180808 4098
rect 180818 4092 180836 4098
rect 181206 4092 181244 4130
rect 181414 4092 181472 4130
rect 182072 4092 182130 4130
rect 182730 4092 182788 4130
rect 182856 4092 182890 10470
rect 183934 5334 184008 5478
rect 183274 4696 183736 5334
rect 183750 4696 184212 5334
rect 185312 4780 185426 4800
rect 185306 4752 185426 4772
rect 183328 4612 183678 4646
rect 183328 4584 183362 4612
rect 183294 4550 183362 4584
rect 183328 4132 183362 4550
rect 183520 4544 183558 4582
rect 183486 4510 183558 4544
rect 183431 4460 183476 4471
rect 183519 4460 183564 4471
rect 183442 4284 183476 4460
rect 183530 4284 183564 4460
rect 183520 4234 183558 4272
rect 183486 4200 183558 4234
rect 183644 4132 183678 4612
rect 183328 4098 183678 4132
rect 183804 4612 184154 4646
rect 183804 4132 183838 4612
rect 183928 4560 183952 4578
rect 183996 4560 184034 4582
rect 183928 4544 184034 4560
rect 183946 4510 184034 4544
rect 183946 4494 183998 4510
rect 183952 4472 183994 4494
rect 184006 4472 184020 4476
rect 183907 4460 183940 4471
rect 183952 4460 183986 4472
rect 183918 4396 183986 4460
rect 183998 4471 184036 4472
rect 183918 4284 183992 4396
rect 183952 4272 183992 4284
rect 183998 4284 184040 4471
rect 183998 4272 184036 4284
rect 183952 4268 183994 4272
rect 183928 4250 183994 4268
rect 183996 4250 184034 4272
rect 183928 4234 184034 4250
rect 183946 4200 184034 4234
rect 183946 4184 183998 4200
rect 183952 4142 183986 4166
rect 184120 4132 184154 4612
rect 183804 4098 184154 4132
rect 179302 4058 180150 4092
rect 180156 4058 180808 4092
rect 180814 4058 183266 4092
rect 183356 4058 183924 4092
rect 179302 3990 179723 4058
rect 180076 4052 180094 4058
rect 180104 4024 180150 4058
rect 180160 4052 180178 4058
rect 180698 4052 180752 4058
rect 180762 4034 180808 4058
rect 180818 4052 180862 4058
rect 180726 4024 180834 4034
rect 180110 3990 180144 4024
rect 180768 3990 180802 4024
rect 181206 3990 181240 4058
rect 181414 4042 181472 4058
rect 182072 4042 182130 4058
rect 182730 4042 182788 4058
rect 182773 4027 182788 4042
rect 182856 3990 182890 4058
rect 179302 3967 184662 3990
rect 170582 3956 184662 3967
rect 165073 3778 165107 3812
rect 164406 3744 164796 3778
rect 164406 3716 164440 3744
rect 164406 3308 164474 3716
rect 164620 3676 164667 3723
rect 164582 3642 164667 3676
rect 164509 3583 164554 3594
rect 164637 3583 164682 3594
rect 164520 3407 164554 3583
rect 164648 3407 164682 3583
rect 164620 3348 164667 3395
rect 164582 3314 164667 3348
rect 164406 3246 164440 3308
rect 164762 3246 164796 3744
rect 164406 3212 164796 3246
rect 164882 3744 165272 3778
rect 164882 3246 164916 3744
rect 165073 3710 165120 3723
rect 165073 3698 165130 3710
rect 165052 3642 165130 3698
rect 164962 3590 164980 3623
rect 165052 3599 165126 3642
rect 165052 3595 165141 3599
rect 164990 3594 165008 3595
rect 165052 3594 165154 3595
rect 164985 3583 165030 3594
rect 164996 3407 165030 3583
rect 165052 3588 165158 3594
rect 165052 3584 165164 3588
rect 165052 3407 165158 3584
rect 165052 3404 165154 3407
rect 165052 3395 165164 3404
rect 165004 3394 165030 3395
rect 165032 3391 165141 3395
rect 165032 3382 165126 3391
rect 165032 3366 165130 3382
rect 165052 3338 165130 3366
rect 165032 3314 165130 3338
rect 165032 3274 165126 3314
rect 165016 3260 165032 3262
rect 165052 3246 165126 3274
rect 165138 3246 165140 3391
rect 165238 3246 165272 3744
rect 164882 3212 165272 3246
rect 165052 3162 165126 3212
rect 163723 2578 163746 2652
rect 163751 2550 163774 2652
rect 164388 2542 164810 3162
rect 164864 2542 165286 3162
rect 167161 2229 167195 3933
rect 168678 3897 169575 3933
rect 171460 2342 171494 3956
rect 171724 3146 171728 3466
rect 171762 3146 171766 3466
rect 172118 2342 172152 3956
rect 172232 2252 172266 3956
rect 174231 3933 179723 3956
rect 174231 3920 174646 3933
rect 173126 3102 173366 3534
rect 172906 3082 172950 3102
rect 173126 3082 173426 3102
rect 173126 3068 173366 3082
rect 172906 3048 172916 3068
rect 173126 3048 173392 3068
rect 173126 2896 173366 3048
rect 177785 2229 177819 3933
rect 179302 3897 179723 3933
rect 180110 2342 180144 3956
rect 182084 2342 182118 3956
rect 182856 2252 182890 3956
rect 183750 3102 183990 3534
rect 183436 3082 183574 3102
rect 183750 3082 184050 3102
rect 183750 3068 183990 3082
rect 183470 3048 183540 3068
rect 183750 3048 184016 3068
rect 183750 2896 183990 3048
rect 164022 1800 164222 1844
rect 163994 1772 164250 1788
rect 117572 -4676 117606 1682
rect 117656 -3498 117680 -3340
rect 117694 -3460 117718 -3378
rect 117990 -4072 118452 -3434
rect 118466 -4072 118928 -3434
rect 118304 -4122 118332 -4088
rect 118044 -4156 118394 -4122
rect 117680 -4630 117694 -4608
rect 118044 -4636 118078 -4156
rect 118236 -4224 118274 -4186
rect 118202 -4258 118274 -4224
rect 118234 -4266 118256 -4262
rect 118147 -4308 118192 -4297
rect 118212 -4300 118220 -4270
rect 118262 -4294 118284 -4262
rect 118304 -4270 118314 -4258
rect 118240 -4297 118248 -4296
rect 118270 -4297 118280 -4294
rect 118235 -4308 118280 -4297
rect 118158 -4484 118192 -4308
rect 118246 -4484 118280 -4308
rect 118270 -4496 118280 -4484
rect 118236 -4500 118280 -4496
rect 118236 -4534 118274 -4500
rect 118304 -4522 118318 -4270
rect 118304 -4534 118314 -4522
rect 118202 -4568 118274 -4534
rect 118326 -4602 118338 -4156
rect 118304 -4626 118338 -4602
rect 118326 -4630 118338 -4626
rect 118360 -4636 118394 -4156
rect 117642 -4670 117658 -4642
rect 116874 -4710 117606 -4676
rect 117614 -4676 117630 -4670
rect 117614 -4698 117634 -4676
rect 117626 -4710 117634 -4698
rect 116874 -4726 116908 -4710
rect 116874 -4737 116885 -4726
rect 116897 -4737 116908 -4726
rect 117572 -4726 117606 -4710
rect 117572 -4737 117583 -4726
rect 117595 -4737 117606 -4726
rect 117660 -4744 117668 -4642
rect 118044 -4670 118394 -4636
rect 118520 -4156 118870 -4122
rect 118520 -4636 118554 -4156
rect 118712 -4224 118750 -4186
rect 118678 -4258 118750 -4224
rect 118623 -4308 118668 -4297
rect 118711 -4308 118756 -4297
rect 118634 -4484 118668 -4308
rect 118722 -4484 118756 -4308
rect 118712 -4534 118750 -4496
rect 118678 -4568 118750 -4534
rect 118836 -4636 118870 -4156
rect 118520 -4670 118870 -4636
rect 117708 -4702 118276 -4676
rect 117708 -4710 118278 -4702
rect 118326 -4744 118342 -4670
rect 118354 -4716 118370 -4670
rect 114018 -4801 120330 -4778
rect 108846 -4848 108891 -4802
rect 108947 -4812 120330 -4801
rect 108947 -4835 115391 -4812
rect 108846 -5468 108880 -4848
rect 108947 -4871 112320 -4835
rect 112838 -4842 112958 -4835
rect 113314 -4842 113434 -4840
rect 114018 -4848 115391 -4835
rect 112832 -4856 112986 -4850
rect 112738 -4869 113060 -4856
rect 113214 -4869 113536 -4856
rect 112832 -4870 112986 -4869
rect 113286 -4870 113462 -4869
rect 108846 -5480 108886 -5468
rect 108868 -5492 108886 -5480
rect 108952 -5492 108986 -4871
rect 109504 -5180 109544 -4871
rect 109504 -5480 109538 -5180
rect 109610 -5492 109644 -4871
rect 110162 -5480 110196 -4871
rect 110206 -5180 110228 -5098
rect 110262 -5180 110302 -4871
rect 110314 -5022 110336 -4871
rect 110268 -5492 110302 -5180
rect 108266 -5524 108334 -5496
rect 108260 -5530 108334 -5524
rect 108344 -5530 108362 -5524
rect 108732 -5530 108770 -5492
rect 108830 -5524 108868 -5492
rect 108886 -5524 108896 -5492
rect 108940 -5530 108998 -5492
rect 109598 -5530 109656 -5492
rect 110256 -5530 110314 -5492
rect 110382 -5530 110416 -4871
rect 110800 -4926 111262 -4871
rect 111276 -4926 111738 -4871
rect 113144 -4926 113384 -4871
rect 110662 -4976 111124 -4954
rect 110662 -5010 111204 -4976
rect 110662 -5490 111124 -5010
rect 111170 -5490 111204 -5010
rect 110662 -5524 111204 -5490
rect 111330 -5010 111680 -4976
rect 111330 -5490 111364 -5010
rect 111454 -5062 111478 -5044
rect 111522 -5062 111560 -5040
rect 111454 -5078 111560 -5062
rect 111472 -5112 111560 -5078
rect 111472 -5128 111524 -5112
rect 111478 -5150 111520 -5128
rect 111532 -5150 111546 -5146
rect 111433 -5162 111466 -5151
rect 111478 -5162 111512 -5150
rect 111444 -5338 111512 -5162
rect 111478 -5350 111512 -5338
rect 111524 -5151 111562 -5150
rect 111524 -5338 111566 -5151
rect 111604 -5160 111628 -5094
rect 111524 -5350 111562 -5338
rect 111478 -5354 111520 -5350
rect 111454 -5372 111520 -5354
rect 111522 -5372 111560 -5350
rect 111454 -5388 111560 -5372
rect 111472 -5422 111560 -5388
rect 111472 -5438 111524 -5422
rect 111478 -5480 111512 -5456
rect 111646 -5490 111680 -5010
rect 112320 -5124 112520 -5098
rect 112876 -5120 112918 -5098
rect 120048 -5132 120120 -5124
rect 120048 -5134 120116 -5132
rect 113394 -5180 113408 -5154
rect 120130 -5352 120150 -5173
rect 120130 -5373 120160 -5352
rect 111330 -5524 111680 -5490
rect 110662 -5530 111124 -5524
rect 99758 -5560 105721 -5553
rect 99758 -5564 102599 -5560
rect 98986 -5632 99020 -5598
rect 99644 -5632 99678 -5595
rect 99758 -5632 99792 -5564
rect 101626 -5580 101660 -5564
rect 101626 -5591 101637 -5580
rect 101649 -5591 101660 -5580
rect 101757 -5587 102599 -5564
rect 102627 -5587 103242 -5560
rect 101757 -5632 102172 -5587
rect 98108 -5655 102172 -5632
rect 102565 -5655 102599 -5587
rect 103223 -5625 103233 -5587
rect 103247 -5625 103257 -5560
rect 103285 -5587 105721 -5560
rect 106828 -5564 107670 -5530
rect 107698 -5564 108334 -5530
rect 108340 -5558 111450 -5530
rect 108340 -5564 110314 -5558
rect 103661 -5655 103695 -5587
rect 103869 -5603 103927 -5587
rect 104527 -5603 104585 -5587
rect 104572 -5655 104573 -5603
rect 104610 -5622 104611 -5587
rect 105048 -5622 105052 -5587
rect 105086 -5622 105090 -5587
rect 105185 -5603 105243 -5587
rect 105197 -5618 105243 -5603
rect 105197 -5655 105231 -5618
rect 105311 -5655 105345 -5587
rect 106828 -5632 107249 -5564
rect 107636 -5618 107670 -5564
rect 108224 -5570 108278 -5564
rect 108288 -5588 108334 -5564
rect 108344 -5570 108388 -5564
rect 108252 -5598 108360 -5588
rect 107602 -5632 107612 -5618
rect 107630 -5632 107670 -5618
rect 108294 -5632 108328 -5598
rect 108732 -5632 108766 -5564
rect 108830 -5632 108868 -5570
rect 108886 -5632 108896 -5570
rect 108940 -5580 108998 -5564
rect 109598 -5580 109656 -5564
rect 110256 -5580 110314 -5564
rect 110299 -5595 110314 -5580
rect 110382 -5564 111450 -5558
rect 110382 -5632 110416 -5564
rect 110662 -5592 111124 -5564
rect 106828 -5655 112188 -5632
rect 98108 -5666 112188 -5655
rect 91932 -5878 92322 -5844
rect 91932 -5906 91966 -5878
rect 91932 -6314 92000 -5906
rect 92146 -5946 92193 -5899
rect 92108 -5980 92193 -5946
rect 92035 -6039 92080 -6028
rect 92163 -6039 92208 -6028
rect 92046 -6215 92080 -6039
rect 92174 -6215 92208 -6039
rect 92146 -6274 92193 -6227
rect 92108 -6308 92193 -6274
rect 91932 -6376 91966 -6314
rect 92288 -6376 92322 -5878
rect 91932 -6410 92322 -6376
rect 92408 -5878 92798 -5844
rect 92408 -6376 92442 -5878
rect 92599 -5899 92633 -5878
rect 92599 -5912 92646 -5899
rect 92599 -5924 92656 -5912
rect 92578 -5980 92656 -5924
rect 92578 -6023 92652 -5980
rect 92578 -6027 92667 -6023
rect 92578 -6028 92680 -6027
rect 92511 -6039 92556 -6028
rect 92522 -6215 92556 -6039
rect 92578 -6215 92684 -6028
rect 92578 -6227 92680 -6215
rect 92578 -6231 92667 -6227
rect 92578 -6240 92652 -6231
rect 92578 -6284 92656 -6240
rect 92558 -6308 92656 -6284
rect 92558 -6348 92652 -6308
rect 92506 -6368 92558 -6360
rect 92578 -6376 92652 -6348
rect 92666 -6368 92720 -6332
rect 92664 -6376 92666 -6368
rect 92764 -6376 92798 -5878
rect 92408 -6410 92798 -6376
rect 92506 -6424 92558 -6410
rect 92578 -6460 92652 -6410
rect 92666 -6424 92720 -6410
rect 91249 -7044 91272 -6970
rect 91277 -7072 91300 -6970
rect 91914 -7080 92336 -6460
rect 92390 -7080 92812 -6460
rect 94573 -7294 94607 -5689
rect 94687 -7393 94721 -5689
rect 96204 -5725 97101 -5689
rect 96978 -5726 96988 -5725
rect 97006 -5726 97044 -5725
rect 97628 -6034 97642 -5726
rect 98986 -7280 99020 -5666
rect 99250 -6476 99254 -6156
rect 99288 -6476 99292 -6156
rect 99644 -7280 99678 -5666
rect 99758 -7370 99792 -5666
rect 101757 -5689 107249 -5666
rect 101757 -5702 102172 -5689
rect 100652 -6520 100892 -6088
rect 100432 -6540 100476 -6520
rect 100652 -6540 100952 -6520
rect 100652 -6554 100892 -6540
rect 100432 -6574 100442 -6554
rect 100652 -6574 100918 -6554
rect 100652 -6726 100892 -6574
rect 105197 -7294 105231 -5689
rect 105311 -7393 105345 -5689
rect 106828 -5725 107249 -5689
rect 107602 -5726 107612 -5666
rect 107630 -5726 107670 -5666
rect 107636 -7280 107670 -5726
rect 108252 -6034 108266 -5726
rect 108830 -6034 108868 -5666
rect 108886 -6034 108896 -5666
rect 109610 -7280 109644 -5666
rect 110382 -7370 110416 -5666
rect 110812 -5676 110970 -5666
rect 120096 -5712 120154 -5710
rect 120070 -5746 120120 -5744
rect 110874 -6088 110908 -6086
rect 110800 -6226 111102 -6088
rect 111276 -6520 111516 -6088
rect 110962 -6540 111100 -6520
rect 111276 -6540 111576 -6520
rect 111276 -6554 111516 -6540
rect 110996 -6574 111066 -6554
rect 111276 -6574 111542 -6554
rect 111276 -6726 111516 -6574
rect 28650 -7455 34962 -7432
rect 23711 -7466 34962 -7455
rect 23711 -7489 30023 -7466
rect 25040 -7525 26010 -7489
rect 28650 -7502 30023 -7489
rect -32992 -7822 -32792 -7778
rect -27400 -7822 -27200 -7778
rect -16066 -7822 -15866 -7778
rect 91548 -7822 91748 -7778
rect -33020 -7850 -32764 -7834
rect -27428 -7850 -27172 -7834
rect -16094 -7850 -15838 -7834
rect 91520 -7850 91776 -7834
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
rect 0 -2400 200 -2200
rect 0 -2800 200 -2600
rect 0 -3200 200 -3000
rect 0 -3600 200 -3400
rect 0 -4000 200 -3800
rect 0 -4400 200 -4200
rect 0 -4800 200 -4600
rect 0 -5200 200 -5000
rect 0 -5600 200 -5400
rect 0 -6000 200 -5800
use buffer  buffer_0
timestamp 1695461801
transform 1 0 76460 0 1 1400
box -6068 -1844 19288 10814
use buffer  buffer_1
timestamp 1695461801
transform 1 0 -27400 0 1 -5568
box -6068 -1844 19288 10814
use buffer  buffer_2
timestamp 1695461801
transform 1 0 -21332 0 1 -7178
box -6068 -1844 19288 10814
use diffamp  diffamp_0
timestamp 1695461801
transform 1 0 -27400 0 1 32314
box 0 -31714 61184 4684
use diffamp  diffamp_1
timestamp 1695461801
transform 1 0 0 0 1 32314
box 0 -31714 61184 4684
use integrator  integrator_0
timestamp 1695461801
transform 1 0 19202 0 1 11168
box 0 -10568 126198 37774
use integrator  integrator_1
timestamp 1695461801
transform 1 0 -27400 0 1 4200
box 0 -10568 126198 37774
use integrator  integrator_2
timestamp 1695461801
transform 1 0 -27400 0 1 1546
box 0 -10568 126198 37774
use mux2_1  mux2_1_0
timestamp 1695461801
transform 1 0 91548 0 1 -7822
box -476 -1200 22640 33492
use mux2_1  mux2_1_1
timestamp 1695461801
transform 1 0 -27400 0 1 -5168
box -476 -1200 22640 33492
use mux2_1  mux2_1_2
timestamp 1695461801
transform 1 0 -32992 0 1 -7822
box -476 -1200 22640 33492
use diffamp  x1
timestamp 1695461801
transform 1 0 0 0 1 28570
box 0 -31714 61184 4684
use integrator  x2
timestamp 1695461801
transform 1 0 57968 0 1 4200
box 0 -10568 126198 37774
use mux2_1  x3
timestamp 1695461801
transform 1 0 164022 0 1 1800
box -476 -1200 22640 33492
use buffer  x7
timestamp 1695461801
transform 1 0 145216 0 1 1400
box -6068 -1844 19288 10814
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 GROUND
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 AIn0
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 AOut
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 AIn1
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 AIn2
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 256 0 0 0 AIn3
port 6 nsew
flabel metal1 0 -2800 200 -2600 0 FreeSans 256 0 0 0 AIn4
port 7 nsew
flabel metal1 0 -3200 200 -3000 0 FreeSans 256 0 0 0 AIn5
port 8 nsew
flabel metal1 0 -3600 200 -3400 0 FreeSans 256 0 0 0 REG0
port 9 nsew
flabel metal1 0 -4000 200 -3800 0 FreeSans 256 0 0 0 REG1
port 10 nsew
flabel metal1 0 -4400 200 -4200 0 FreeSans 256 0 0 0 REG2
port 11 nsew
flabel metal1 0 -4800 200 -4600 0 FreeSans 256 0 0 0 REG3
port 12 nsew
flabel metal1 0 -5200 200 -5000 0 FreeSans 256 0 0 0 REG4
port 13 nsew
flabel metal1 0 -5600 200 -5400 0 FreeSans 256 0 0 0 REG5
port 14 nsew
flabel metal1 0 -6000 200 -5800 0 FreeSans 256 0 0 0 REG6
port 15 nsew
<< end >>
