magic
tech sky130A
timestamp 1695908076
<< pwell >>
rect -906 -2105 906 2105
<< nmoslvt >>
rect -808 -2000 -508 2000
rect -479 -2000 -179 2000
rect -150 -2000 150 2000
rect 179 -2000 479 2000
rect 508 -2000 808 2000
<< ndiff >>
rect -837 1994 -808 2000
rect -837 -1994 -831 1994
rect -814 -1994 -808 1994
rect -837 -2000 -808 -1994
rect -508 1994 -479 2000
rect -508 -1994 -502 1994
rect -485 -1994 -479 1994
rect -508 -2000 -479 -1994
rect -179 1994 -150 2000
rect -179 -1994 -173 1994
rect -156 -1994 -150 1994
rect -179 -2000 -150 -1994
rect 150 1994 179 2000
rect 150 -1994 156 1994
rect 173 -1994 179 1994
rect 150 -2000 179 -1994
rect 479 1994 508 2000
rect 479 -1994 485 1994
rect 502 -1994 508 1994
rect 479 -2000 508 -1994
rect 808 1994 837 2000
rect 808 -1994 814 1994
rect 831 -1994 837 1994
rect 808 -2000 837 -1994
<< ndiffc >>
rect -831 -1994 -814 1994
rect -502 -1994 -485 1994
rect -173 -1994 -156 1994
rect 156 -1994 173 1994
rect 485 -1994 502 1994
rect 814 -1994 831 1994
<< psubdiff >>
rect -888 2070 -840 2087
rect 840 2070 888 2087
rect -888 2039 -871 2070
rect 871 2039 888 2070
rect -888 -2070 -871 -2039
rect 871 -2070 888 -2039
rect -888 -2087 -840 -2070
rect 840 -2087 888 -2070
<< psubdiffcont >>
rect -840 2070 840 2087
rect -888 -2039 -871 2039
rect 871 -2039 888 2039
rect -840 -2087 840 -2070
<< poly >>
rect -808 2036 -508 2044
rect -808 2019 -800 2036
rect -516 2019 -508 2036
rect -808 2000 -508 2019
rect -479 2036 -179 2044
rect -479 2019 -471 2036
rect -187 2019 -179 2036
rect -479 2000 -179 2019
rect -150 2036 150 2044
rect -150 2019 -142 2036
rect 142 2019 150 2036
rect -150 2000 150 2019
rect 179 2036 479 2044
rect 179 2019 187 2036
rect 471 2019 479 2036
rect 179 2000 479 2019
rect 508 2036 808 2044
rect 508 2019 516 2036
rect 800 2019 808 2036
rect 508 2000 808 2019
rect -808 -2019 -508 -2000
rect -808 -2036 -800 -2019
rect -516 -2036 -508 -2019
rect -808 -2044 -508 -2036
rect -479 -2019 -179 -2000
rect -479 -2036 -471 -2019
rect -187 -2036 -179 -2019
rect -479 -2044 -179 -2036
rect -150 -2019 150 -2000
rect -150 -2036 -142 -2019
rect 142 -2036 150 -2019
rect -150 -2044 150 -2036
rect 179 -2019 479 -2000
rect 179 -2036 187 -2019
rect 471 -2036 479 -2019
rect 179 -2044 479 -2036
rect 508 -2019 808 -2000
rect 508 -2036 516 -2019
rect 800 -2036 808 -2019
rect 508 -2044 808 -2036
<< polycont >>
rect -800 2019 -516 2036
rect -471 2019 -187 2036
rect -142 2019 142 2036
rect 187 2019 471 2036
rect 516 2019 800 2036
rect -800 -2036 -516 -2019
rect -471 -2036 -187 -2019
rect -142 -2036 142 -2019
rect 187 -2036 471 -2019
rect 516 -2036 800 -2019
<< locali >>
rect -888 2070 -840 2087
rect 840 2070 888 2087
rect -888 2039 -871 2070
rect 871 2039 888 2070
rect -808 2019 -800 2036
rect -516 2019 -508 2036
rect -479 2019 -471 2036
rect -187 2019 -179 2036
rect -150 2019 -142 2036
rect 142 2019 150 2036
rect 179 2019 187 2036
rect 471 2019 479 2036
rect 508 2019 516 2036
rect 800 2019 808 2036
rect -831 1994 -814 2002
rect -831 -2002 -814 -1994
rect -502 1994 -485 2002
rect -502 -2002 -485 -1994
rect -173 1994 -156 2002
rect -173 -2002 -156 -1994
rect 156 1994 173 2002
rect 156 -2002 173 -1994
rect 485 1994 502 2002
rect 485 -2002 502 -1994
rect 814 1994 831 2002
rect 814 -2002 831 -1994
rect -808 -2036 -800 -2019
rect -516 -2036 -508 -2019
rect -479 -2036 -471 -2019
rect -187 -2036 -179 -2019
rect -150 -2036 -142 -2019
rect 142 -2036 150 -2019
rect 179 -2036 187 -2019
rect 471 -2036 479 -2019
rect 508 -2036 516 -2019
rect 800 -2036 808 -2019
rect -888 -2070 -871 -2039
rect 871 -2070 888 -2039
rect -888 -2087 -840 -2070
rect 840 -2087 888 -2070
<< viali >>
rect -800 2019 -516 2036
rect -471 2019 -187 2036
rect -142 2019 142 2036
rect 187 2019 471 2036
rect 516 2019 800 2036
rect -831 -1994 -814 1994
rect -502 -1994 -485 1994
rect -173 -1994 -156 1994
rect 156 -1994 173 1994
rect 485 -1994 502 1994
rect 814 -1994 831 1994
rect -800 -2036 -516 -2019
rect -471 -2036 -187 -2019
rect -142 -2036 142 -2019
rect 187 -2036 471 -2019
rect 516 -2036 800 -2019
<< metal1 >>
rect -806 2036 -510 2039
rect -806 2019 -800 2036
rect -516 2019 -510 2036
rect -806 2016 -510 2019
rect -477 2036 -181 2039
rect -477 2019 -471 2036
rect -187 2019 -181 2036
rect -477 2016 -181 2019
rect -148 2036 148 2039
rect -148 2019 -142 2036
rect 142 2019 148 2036
rect -148 2016 148 2019
rect 181 2036 477 2039
rect 181 2019 187 2036
rect 471 2019 477 2036
rect 181 2016 477 2019
rect 510 2036 806 2039
rect 510 2019 516 2036
rect 800 2019 806 2036
rect 510 2016 806 2019
rect -834 1994 -811 2000
rect -834 -1994 -831 1994
rect -814 -1994 -811 1994
rect -834 -2000 -811 -1994
rect -505 1994 -482 2000
rect -505 -1994 -502 1994
rect -485 -1994 -482 1994
rect -505 -2000 -482 -1994
rect -176 1994 -153 2000
rect -176 -1994 -173 1994
rect -156 -1994 -153 1994
rect -176 -2000 -153 -1994
rect 153 1994 176 2000
rect 153 -1994 156 1994
rect 173 -1994 176 1994
rect 153 -2000 176 -1994
rect 482 1994 505 2000
rect 482 -1994 485 1994
rect 502 -1994 505 1994
rect 482 -2000 505 -1994
rect 811 1994 834 2000
rect 811 -1994 814 1994
rect 831 -1994 834 1994
rect 811 -2000 834 -1994
rect -806 -2019 -510 -2016
rect -806 -2036 -800 -2019
rect -516 -2036 -510 -2019
rect -806 -2039 -510 -2036
rect -477 -2019 -181 -2016
rect -477 -2036 -471 -2019
rect -187 -2036 -181 -2019
rect -477 -2039 -181 -2036
rect -148 -2019 148 -2016
rect -148 -2036 -142 -2019
rect 142 -2036 148 -2019
rect -148 -2039 148 -2036
rect 181 -2019 477 -2016
rect 181 -2036 187 -2019
rect 471 -2036 477 -2019
rect 181 -2039 477 -2036
rect 510 -2019 806 -2016
rect 510 -2036 516 -2019
rect 800 -2036 806 -2019
rect 510 -2039 806 -2036
<< labels >>
rlabel poly -150 2000 150 2019 1 G
rlabel locali -831 1994 -814 2002 1 D
rlabel psubdiffcont -840 2070 840 2087 1 B
rlabel locali 814 1994 831 2002 1 S
<< properties >>
string FIXED_BBOX -879 -2078 879 2078
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 40.0 l 3.0 m 1 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
