magic
tech sky130A
magscale 1 2
timestamp 1696133064
<< nwell >>
rect -4754 -3219 4754 3219
<< pmoslvt >>
rect -4558 -3000 -1558 3000
rect -1500 -3000 1500 3000
rect 1558 -3000 4558 3000
<< pdiff >>
rect -4616 2988 -4558 3000
rect -4616 -2988 -4604 2988
rect -4570 -2988 -4558 2988
rect -4616 -3000 -4558 -2988
rect -1558 2988 -1500 3000
rect -1558 -2988 -1546 2988
rect -1512 -2988 -1500 2988
rect -1558 -3000 -1500 -2988
rect 1500 2988 1558 3000
rect 1500 -2988 1512 2988
rect 1546 -2988 1558 2988
rect 1500 -3000 1558 -2988
rect 4558 2988 4616 3000
rect 4558 -2988 4570 2988
rect 4604 -2988 4616 2988
rect 4558 -3000 4616 -2988
<< pdiffc >>
rect -4604 -2988 -4570 2988
rect -1546 -2988 -1512 2988
rect 1512 -2988 1546 2988
rect 4570 -2988 4604 2988
<< nsubdiff >>
rect -4718 3149 -4622 3183
rect 4622 3149 4718 3183
rect -4718 3087 -4684 3149
rect 4684 3087 4718 3149
rect -4718 -3149 -4684 -3087
rect 4684 -3149 4718 -3087
rect -4718 -3183 -4622 -3149
rect 4622 -3183 4718 -3149
<< nsubdiffcont >>
rect -4622 3149 4622 3183
rect -4718 -3087 -4684 3087
rect 4684 -3087 4718 3087
rect -4622 -3183 4622 -3149
<< poly >>
rect -4558 3081 -1558 3097
rect -4558 3047 -4542 3081
rect -1574 3047 -1558 3081
rect -4558 3000 -1558 3047
rect -1500 3081 1500 3097
rect -1500 3047 -1484 3081
rect 1484 3047 1500 3081
rect -1500 3000 1500 3047
rect 1558 3081 4558 3097
rect 1558 3047 1574 3081
rect 4542 3047 4558 3081
rect 1558 3000 4558 3047
rect -4558 -3047 -1558 -3000
rect -4558 -3081 -4542 -3047
rect -1574 -3081 -1558 -3047
rect -4558 -3097 -1558 -3081
rect -1500 -3047 1500 -3000
rect -1500 -3081 -1484 -3047
rect 1484 -3081 1500 -3047
rect -1500 -3097 1500 -3081
rect 1558 -3047 4558 -3000
rect 1558 -3081 1574 -3047
rect 4542 -3081 4558 -3047
rect 1558 -3097 4558 -3081
<< polycont >>
rect -4542 3047 -1574 3081
rect -1484 3047 1484 3081
rect 1574 3047 4542 3081
rect -4542 -3081 -1574 -3047
rect -1484 -3081 1484 -3047
rect 1574 -3081 4542 -3047
<< locali >>
rect -4718 3149 -4622 3183
rect 4622 3149 4718 3183
rect -4718 3087 -4684 3149
rect 4684 3087 4718 3149
rect -4558 3047 -4542 3081
rect -1574 3047 -1558 3081
rect -1500 3047 -1484 3081
rect 1484 3047 1500 3081
rect 1558 3047 1574 3081
rect 4542 3047 4558 3081
rect -4604 2988 -4570 3004
rect -4604 -3004 -4570 -2988
rect -1546 2988 -1512 3004
rect -1546 -3004 -1512 -2988
rect 1512 2988 1546 3004
rect 1512 -3004 1546 -2988
rect 4570 2988 4604 3004
rect 4570 -3004 4604 -2988
rect -4558 -3081 -4542 -3047
rect -1574 -3081 -1558 -3047
rect -1500 -3081 -1484 -3047
rect 1484 -3081 1500 -3047
rect 1558 -3081 1574 -3047
rect 4542 -3081 4558 -3047
rect -4718 -3149 -4684 -3087
rect 4684 -3149 4718 -3087
rect -4718 -3183 -4622 -3149
rect 4622 -3183 4718 -3149
<< viali >>
rect -4542 3047 -1574 3081
rect -1484 3047 1484 3081
rect 1574 3047 4542 3081
rect -4604 -2988 -4570 2988
rect -1546 -2988 -1512 2988
rect 1512 -2988 1546 2988
rect 4570 -2988 4604 2988
rect -4542 -3081 -1574 -3047
rect -1484 -3081 1484 -3047
rect 1574 -3081 4542 -3047
<< metal1 >>
rect -4554 3081 -1562 3087
rect -4554 3047 -4542 3081
rect -1574 3047 -1562 3081
rect -4554 3041 -1562 3047
rect -1496 3081 1496 3087
rect -1496 3047 -1484 3081
rect 1484 3047 1496 3081
rect -1496 3041 1496 3047
rect 1562 3081 4554 3087
rect 1562 3047 1574 3081
rect 4542 3047 4554 3081
rect 1562 3041 4554 3047
rect -4610 2988 -4564 3000
rect -4610 -2988 -4604 2988
rect -4570 -2988 -4564 2988
rect -4610 -3000 -4564 -2988
rect -1552 2988 -1506 3000
rect -1552 -2988 -1546 2988
rect -1512 -2988 -1506 2988
rect -1552 -3000 -1506 -2988
rect 1506 2988 1552 3000
rect 1506 -2988 1512 2988
rect 1546 -2988 1552 2988
rect 1506 -3000 1552 -2988
rect 4564 2988 4610 3000
rect 4564 -2988 4570 2988
rect 4604 -2988 4610 2988
rect 4564 -3000 4610 -2988
rect -4554 -3047 -1562 -3041
rect -4554 -3081 -4542 -3047
rect -1574 -3081 -1562 -3047
rect -4554 -3087 -1562 -3081
rect -1496 -3047 1496 -3041
rect -1496 -3081 -1484 -3047
rect 1484 -3081 1496 -3047
rect -1496 -3087 1496 -3081
rect 1562 -3047 4554 -3041
rect 1562 -3081 1574 -3047
rect 4542 -3081 4554 -3047
rect 1562 -3087 4554 -3081
<< properties >>
string FIXED_BBOX -4701 -3166 4701 3166
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 30.0 l 15.0 m 1 nf 3 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
