magic
tech sky130A
magscale 1 2
timestamp 1694848836
<< pwell >>
rect -6747 -260 6747 260
<< nmoslvt >>
rect -6551 -50 -5951 50
rect -5893 -50 -5293 50
rect -5235 -50 -4635 50
rect -4577 -50 -3977 50
rect -3919 -50 -3319 50
rect -3261 -50 -2661 50
rect -2603 -50 -2003 50
rect -1945 -50 -1345 50
rect -1287 -50 -687 50
rect -629 -50 -29 50
rect 29 -50 629 50
rect 687 -50 1287 50
rect 1345 -50 1945 50
rect 2003 -50 2603 50
rect 2661 -50 3261 50
rect 3319 -50 3919 50
rect 3977 -50 4577 50
rect 4635 -50 5235 50
rect 5293 -50 5893 50
rect 5951 -50 6551 50
<< ndiff >>
rect -6609 38 -6551 50
rect -6609 -38 -6597 38
rect -6563 -38 -6551 38
rect -6609 -50 -6551 -38
rect -5951 38 -5893 50
rect -5951 -38 -5939 38
rect -5905 -38 -5893 38
rect -5951 -50 -5893 -38
rect -5293 38 -5235 50
rect -5293 -38 -5281 38
rect -5247 -38 -5235 38
rect -5293 -50 -5235 -38
rect -4635 38 -4577 50
rect -4635 -38 -4623 38
rect -4589 -38 -4577 38
rect -4635 -50 -4577 -38
rect -3977 38 -3919 50
rect -3977 -38 -3965 38
rect -3931 -38 -3919 38
rect -3977 -50 -3919 -38
rect -3319 38 -3261 50
rect -3319 -38 -3307 38
rect -3273 -38 -3261 38
rect -3319 -50 -3261 -38
rect -2661 38 -2603 50
rect -2661 -38 -2649 38
rect -2615 -38 -2603 38
rect -2661 -50 -2603 -38
rect -2003 38 -1945 50
rect -2003 -38 -1991 38
rect -1957 -38 -1945 38
rect -2003 -50 -1945 -38
rect -1345 38 -1287 50
rect -1345 -38 -1333 38
rect -1299 -38 -1287 38
rect -1345 -50 -1287 -38
rect -687 38 -629 50
rect -687 -38 -675 38
rect -641 -38 -629 38
rect -687 -50 -629 -38
rect -29 38 29 50
rect -29 -38 -17 38
rect 17 -38 29 38
rect -29 -50 29 -38
rect 629 38 687 50
rect 629 -38 641 38
rect 675 -38 687 38
rect 629 -50 687 -38
rect 1287 38 1345 50
rect 1287 -38 1299 38
rect 1333 -38 1345 38
rect 1287 -50 1345 -38
rect 1945 38 2003 50
rect 1945 -38 1957 38
rect 1991 -38 2003 38
rect 1945 -50 2003 -38
rect 2603 38 2661 50
rect 2603 -38 2615 38
rect 2649 -38 2661 38
rect 2603 -50 2661 -38
rect 3261 38 3319 50
rect 3261 -38 3273 38
rect 3307 -38 3319 38
rect 3261 -50 3319 -38
rect 3919 38 3977 50
rect 3919 -38 3931 38
rect 3965 -38 3977 38
rect 3919 -50 3977 -38
rect 4577 38 4635 50
rect 4577 -38 4589 38
rect 4623 -38 4635 38
rect 4577 -50 4635 -38
rect 5235 38 5293 50
rect 5235 -38 5247 38
rect 5281 -38 5293 38
rect 5235 -50 5293 -38
rect 5893 38 5951 50
rect 5893 -38 5905 38
rect 5939 -38 5951 38
rect 5893 -50 5951 -38
rect 6551 38 6609 50
rect 6551 -38 6563 38
rect 6597 -38 6609 38
rect 6551 -50 6609 -38
<< ndiffc >>
rect -6597 -38 -6563 38
rect -5939 -38 -5905 38
rect -5281 -38 -5247 38
rect -4623 -38 -4589 38
rect -3965 -38 -3931 38
rect -3307 -38 -3273 38
rect -2649 -38 -2615 38
rect -1991 -38 -1957 38
rect -1333 -38 -1299 38
rect -675 -38 -641 38
rect -17 -38 17 38
rect 641 -38 675 38
rect 1299 -38 1333 38
rect 1957 -38 1991 38
rect 2615 -38 2649 38
rect 3273 -38 3307 38
rect 3931 -38 3965 38
rect 4589 -38 4623 38
rect 5247 -38 5281 38
rect 5905 -38 5939 38
rect 6563 -38 6597 38
<< psubdiff >>
rect -6711 190 -6615 224
rect 6615 190 6711 224
rect -6711 128 -6677 190
rect 6677 128 6711 190
rect -6711 -190 -6677 -128
rect 6677 -190 6711 -128
rect -6711 -224 -6615 -190
rect 6615 -224 6711 -190
<< psubdiffcont >>
rect -6615 190 6615 224
rect -6711 -128 -6677 128
rect 6677 -128 6711 128
rect -6615 -224 6615 -190
<< poly >>
rect -6551 122 -5951 138
rect -6551 88 -6535 122
rect -5967 88 -5951 122
rect -6551 50 -5951 88
rect -5893 122 -5293 138
rect -5893 88 -5877 122
rect -5309 88 -5293 122
rect -5893 50 -5293 88
rect -5235 122 -4635 138
rect -5235 88 -5219 122
rect -4651 88 -4635 122
rect -5235 50 -4635 88
rect -4577 122 -3977 138
rect -4577 88 -4561 122
rect -3993 88 -3977 122
rect -4577 50 -3977 88
rect -3919 122 -3319 138
rect -3919 88 -3903 122
rect -3335 88 -3319 122
rect -3919 50 -3319 88
rect -3261 122 -2661 138
rect -3261 88 -3245 122
rect -2677 88 -2661 122
rect -3261 50 -2661 88
rect -2603 122 -2003 138
rect -2603 88 -2587 122
rect -2019 88 -2003 122
rect -2603 50 -2003 88
rect -1945 122 -1345 138
rect -1945 88 -1929 122
rect -1361 88 -1345 122
rect -1945 50 -1345 88
rect -1287 122 -687 138
rect -1287 88 -1271 122
rect -703 88 -687 122
rect -1287 50 -687 88
rect -629 122 -29 138
rect -629 88 -613 122
rect -45 88 -29 122
rect -629 50 -29 88
rect 29 122 629 138
rect 29 88 45 122
rect 613 88 629 122
rect 29 50 629 88
rect 687 122 1287 138
rect 687 88 703 122
rect 1271 88 1287 122
rect 687 50 1287 88
rect 1345 122 1945 138
rect 1345 88 1361 122
rect 1929 88 1945 122
rect 1345 50 1945 88
rect 2003 122 2603 138
rect 2003 88 2019 122
rect 2587 88 2603 122
rect 2003 50 2603 88
rect 2661 122 3261 138
rect 2661 88 2677 122
rect 3245 88 3261 122
rect 2661 50 3261 88
rect 3319 122 3919 138
rect 3319 88 3335 122
rect 3903 88 3919 122
rect 3319 50 3919 88
rect 3977 122 4577 138
rect 3977 88 3993 122
rect 4561 88 4577 122
rect 3977 50 4577 88
rect 4635 122 5235 138
rect 4635 88 4651 122
rect 5219 88 5235 122
rect 4635 50 5235 88
rect 5293 122 5893 138
rect 5293 88 5309 122
rect 5877 88 5893 122
rect 5293 50 5893 88
rect 5951 122 6551 138
rect 5951 88 5967 122
rect 6535 88 6551 122
rect 5951 50 6551 88
rect -6551 -88 -5951 -50
rect -6551 -122 -6535 -88
rect -5967 -122 -5951 -88
rect -6551 -138 -5951 -122
rect -5893 -88 -5293 -50
rect -5893 -122 -5877 -88
rect -5309 -122 -5293 -88
rect -5893 -138 -5293 -122
rect -5235 -88 -4635 -50
rect -5235 -122 -5219 -88
rect -4651 -122 -4635 -88
rect -5235 -138 -4635 -122
rect -4577 -88 -3977 -50
rect -4577 -122 -4561 -88
rect -3993 -122 -3977 -88
rect -4577 -138 -3977 -122
rect -3919 -88 -3319 -50
rect -3919 -122 -3903 -88
rect -3335 -122 -3319 -88
rect -3919 -138 -3319 -122
rect -3261 -88 -2661 -50
rect -3261 -122 -3245 -88
rect -2677 -122 -2661 -88
rect -3261 -138 -2661 -122
rect -2603 -88 -2003 -50
rect -2603 -122 -2587 -88
rect -2019 -122 -2003 -88
rect -2603 -138 -2003 -122
rect -1945 -88 -1345 -50
rect -1945 -122 -1929 -88
rect -1361 -122 -1345 -88
rect -1945 -138 -1345 -122
rect -1287 -88 -687 -50
rect -1287 -122 -1271 -88
rect -703 -122 -687 -88
rect -1287 -138 -687 -122
rect -629 -88 -29 -50
rect -629 -122 -613 -88
rect -45 -122 -29 -88
rect -629 -138 -29 -122
rect 29 -88 629 -50
rect 29 -122 45 -88
rect 613 -122 629 -88
rect 29 -138 629 -122
rect 687 -88 1287 -50
rect 687 -122 703 -88
rect 1271 -122 1287 -88
rect 687 -138 1287 -122
rect 1345 -88 1945 -50
rect 1345 -122 1361 -88
rect 1929 -122 1945 -88
rect 1345 -138 1945 -122
rect 2003 -88 2603 -50
rect 2003 -122 2019 -88
rect 2587 -122 2603 -88
rect 2003 -138 2603 -122
rect 2661 -88 3261 -50
rect 2661 -122 2677 -88
rect 3245 -122 3261 -88
rect 2661 -138 3261 -122
rect 3319 -88 3919 -50
rect 3319 -122 3335 -88
rect 3903 -122 3919 -88
rect 3319 -138 3919 -122
rect 3977 -88 4577 -50
rect 3977 -122 3993 -88
rect 4561 -122 4577 -88
rect 3977 -138 4577 -122
rect 4635 -88 5235 -50
rect 4635 -122 4651 -88
rect 5219 -122 5235 -88
rect 4635 -138 5235 -122
rect 5293 -88 5893 -50
rect 5293 -122 5309 -88
rect 5877 -122 5893 -88
rect 5293 -138 5893 -122
rect 5951 -88 6551 -50
rect 5951 -122 5967 -88
rect 6535 -122 6551 -88
rect 5951 -138 6551 -122
<< polycont >>
rect -6535 88 -5967 122
rect -5877 88 -5309 122
rect -5219 88 -4651 122
rect -4561 88 -3993 122
rect -3903 88 -3335 122
rect -3245 88 -2677 122
rect -2587 88 -2019 122
rect -1929 88 -1361 122
rect -1271 88 -703 122
rect -613 88 -45 122
rect 45 88 613 122
rect 703 88 1271 122
rect 1361 88 1929 122
rect 2019 88 2587 122
rect 2677 88 3245 122
rect 3335 88 3903 122
rect 3993 88 4561 122
rect 4651 88 5219 122
rect 5309 88 5877 122
rect 5967 88 6535 122
rect -6535 -122 -5967 -88
rect -5877 -122 -5309 -88
rect -5219 -122 -4651 -88
rect -4561 -122 -3993 -88
rect -3903 -122 -3335 -88
rect -3245 -122 -2677 -88
rect -2587 -122 -2019 -88
rect -1929 -122 -1361 -88
rect -1271 -122 -703 -88
rect -613 -122 -45 -88
rect 45 -122 613 -88
rect 703 -122 1271 -88
rect 1361 -122 1929 -88
rect 2019 -122 2587 -88
rect 2677 -122 3245 -88
rect 3335 -122 3903 -88
rect 3993 -122 4561 -88
rect 4651 -122 5219 -88
rect 5309 -122 5877 -88
rect 5967 -122 6535 -88
<< locali >>
rect -6711 190 -6615 224
rect 6615 190 6711 224
rect -6711 128 -6677 190
rect 6677 128 6711 190
rect -6551 88 -6535 122
rect -5967 88 -5951 122
rect -5893 88 -5877 122
rect -5309 88 -5293 122
rect -5235 88 -5219 122
rect -4651 88 -4635 122
rect -4577 88 -4561 122
rect -3993 88 -3977 122
rect -3919 88 -3903 122
rect -3335 88 -3319 122
rect -3261 88 -3245 122
rect -2677 88 -2661 122
rect -2603 88 -2587 122
rect -2019 88 -2003 122
rect -1945 88 -1929 122
rect -1361 88 -1345 122
rect -1287 88 -1271 122
rect -703 88 -687 122
rect -629 88 -613 122
rect -45 88 -29 122
rect 29 88 45 122
rect 613 88 629 122
rect 687 88 703 122
rect 1271 88 1287 122
rect 1345 88 1361 122
rect 1929 88 1945 122
rect 2003 88 2019 122
rect 2587 88 2603 122
rect 2661 88 2677 122
rect 3245 88 3261 122
rect 3319 88 3335 122
rect 3903 88 3919 122
rect 3977 88 3993 122
rect 4561 88 4577 122
rect 4635 88 4651 122
rect 5219 88 5235 122
rect 5293 88 5309 122
rect 5877 88 5893 122
rect 5951 88 5967 122
rect 6535 88 6551 122
rect -6597 38 -6563 54
rect -6597 -54 -6563 -38
rect -5939 38 -5905 54
rect -5939 -54 -5905 -38
rect -5281 38 -5247 54
rect -5281 -54 -5247 -38
rect -4623 38 -4589 54
rect -4623 -54 -4589 -38
rect -3965 38 -3931 54
rect -3965 -54 -3931 -38
rect -3307 38 -3273 54
rect -3307 -54 -3273 -38
rect -2649 38 -2615 54
rect -2649 -54 -2615 -38
rect -1991 38 -1957 54
rect -1991 -54 -1957 -38
rect -1333 38 -1299 54
rect -1333 -54 -1299 -38
rect -675 38 -641 54
rect -675 -54 -641 -38
rect -17 38 17 54
rect -17 -54 17 -38
rect 641 38 675 54
rect 641 -54 675 -38
rect 1299 38 1333 54
rect 1299 -54 1333 -38
rect 1957 38 1991 54
rect 1957 -54 1991 -38
rect 2615 38 2649 54
rect 2615 -54 2649 -38
rect 3273 38 3307 54
rect 3273 -54 3307 -38
rect 3931 38 3965 54
rect 3931 -54 3965 -38
rect 4589 38 4623 54
rect 4589 -54 4623 -38
rect 5247 38 5281 54
rect 5247 -54 5281 -38
rect 5905 38 5939 54
rect 5905 -54 5939 -38
rect 6563 38 6597 54
rect 6563 -54 6597 -38
rect -6551 -122 -6535 -88
rect -5967 -122 -5951 -88
rect -5893 -122 -5877 -88
rect -5309 -122 -5293 -88
rect -5235 -122 -5219 -88
rect -4651 -122 -4635 -88
rect -4577 -122 -4561 -88
rect -3993 -122 -3977 -88
rect -3919 -122 -3903 -88
rect -3335 -122 -3319 -88
rect -3261 -122 -3245 -88
rect -2677 -122 -2661 -88
rect -2603 -122 -2587 -88
rect -2019 -122 -2003 -88
rect -1945 -122 -1929 -88
rect -1361 -122 -1345 -88
rect -1287 -122 -1271 -88
rect -703 -122 -687 -88
rect -629 -122 -613 -88
rect -45 -122 -29 -88
rect 29 -122 45 -88
rect 613 -122 629 -88
rect 687 -122 703 -88
rect 1271 -122 1287 -88
rect 1345 -122 1361 -88
rect 1929 -122 1945 -88
rect 2003 -122 2019 -88
rect 2587 -122 2603 -88
rect 2661 -122 2677 -88
rect 3245 -122 3261 -88
rect 3319 -122 3335 -88
rect 3903 -122 3919 -88
rect 3977 -122 3993 -88
rect 4561 -122 4577 -88
rect 4635 -122 4651 -88
rect 5219 -122 5235 -88
rect 5293 -122 5309 -88
rect 5877 -122 5893 -88
rect 5951 -122 5967 -88
rect 6535 -122 6551 -88
rect -6711 -190 -6677 -128
rect 6677 -190 6711 -128
rect -6711 -224 -6615 -190
rect 6615 -224 6711 -190
<< viali >>
rect -6535 88 -5967 122
rect -5877 88 -5309 122
rect -5219 88 -4651 122
rect -4561 88 -3993 122
rect -3903 88 -3335 122
rect -3245 88 -2677 122
rect -2587 88 -2019 122
rect -1929 88 -1361 122
rect -1271 88 -703 122
rect -613 88 -45 122
rect 45 88 613 122
rect 703 88 1271 122
rect 1361 88 1929 122
rect 2019 88 2587 122
rect 2677 88 3245 122
rect 3335 88 3903 122
rect 3993 88 4561 122
rect 4651 88 5219 122
rect 5309 88 5877 122
rect 5967 88 6535 122
rect -6597 -38 -6563 38
rect -5939 -38 -5905 38
rect -5281 -38 -5247 38
rect -4623 -38 -4589 38
rect -3965 -38 -3931 38
rect -3307 -38 -3273 38
rect -2649 -38 -2615 38
rect -1991 -38 -1957 38
rect -1333 -38 -1299 38
rect -675 -38 -641 38
rect -17 -38 17 38
rect 641 -38 675 38
rect 1299 -38 1333 38
rect 1957 -38 1991 38
rect 2615 -38 2649 38
rect 3273 -38 3307 38
rect 3931 -38 3965 38
rect 4589 -38 4623 38
rect 5247 -38 5281 38
rect 5905 -38 5939 38
rect 6563 -38 6597 38
rect -6535 -122 -5967 -88
rect -5877 -122 -5309 -88
rect -5219 -122 -4651 -88
rect -4561 -122 -3993 -88
rect -3903 -122 -3335 -88
rect -3245 -122 -2677 -88
rect -2587 -122 -2019 -88
rect -1929 -122 -1361 -88
rect -1271 -122 -703 -88
rect -613 -122 -45 -88
rect 45 -122 613 -88
rect 703 -122 1271 -88
rect 1361 -122 1929 -88
rect 2019 -122 2587 -88
rect 2677 -122 3245 -88
rect 3335 -122 3903 -88
rect 3993 -122 4561 -88
rect 4651 -122 5219 -88
rect 5309 -122 5877 -88
rect 5967 -122 6535 -88
<< metal1 >>
rect -6547 122 -5955 128
rect -6547 88 -6535 122
rect -5967 88 -5955 122
rect -6547 82 -5955 88
rect -5889 122 -5297 128
rect -5889 88 -5877 122
rect -5309 88 -5297 122
rect -5889 82 -5297 88
rect -5231 122 -4639 128
rect -5231 88 -5219 122
rect -4651 88 -4639 122
rect -5231 82 -4639 88
rect -4573 122 -3981 128
rect -4573 88 -4561 122
rect -3993 88 -3981 122
rect -4573 82 -3981 88
rect -3915 122 -3323 128
rect -3915 88 -3903 122
rect -3335 88 -3323 122
rect -3915 82 -3323 88
rect -3257 122 -2665 128
rect -3257 88 -3245 122
rect -2677 88 -2665 122
rect -3257 82 -2665 88
rect -2599 122 -2007 128
rect -2599 88 -2587 122
rect -2019 88 -2007 122
rect -2599 82 -2007 88
rect -1941 122 -1349 128
rect -1941 88 -1929 122
rect -1361 88 -1349 122
rect -1941 82 -1349 88
rect -1283 122 -691 128
rect -1283 88 -1271 122
rect -703 88 -691 122
rect -1283 82 -691 88
rect -625 122 -33 128
rect -625 88 -613 122
rect -45 88 -33 122
rect -625 82 -33 88
rect 33 122 625 128
rect 33 88 45 122
rect 613 88 625 122
rect 33 82 625 88
rect 691 122 1283 128
rect 691 88 703 122
rect 1271 88 1283 122
rect 691 82 1283 88
rect 1349 122 1941 128
rect 1349 88 1361 122
rect 1929 88 1941 122
rect 1349 82 1941 88
rect 2007 122 2599 128
rect 2007 88 2019 122
rect 2587 88 2599 122
rect 2007 82 2599 88
rect 2665 122 3257 128
rect 2665 88 2677 122
rect 3245 88 3257 122
rect 2665 82 3257 88
rect 3323 122 3915 128
rect 3323 88 3335 122
rect 3903 88 3915 122
rect 3323 82 3915 88
rect 3981 122 4573 128
rect 3981 88 3993 122
rect 4561 88 4573 122
rect 3981 82 4573 88
rect 4639 122 5231 128
rect 4639 88 4651 122
rect 5219 88 5231 122
rect 4639 82 5231 88
rect 5297 122 5889 128
rect 5297 88 5309 122
rect 5877 88 5889 122
rect 5297 82 5889 88
rect 5955 122 6547 128
rect 5955 88 5967 122
rect 6535 88 6547 122
rect 5955 82 6547 88
rect -6603 38 -6557 50
rect -6603 -38 -6597 38
rect -6563 -38 -6557 38
rect -6603 -50 -6557 -38
rect -5945 38 -5899 50
rect -5945 -38 -5939 38
rect -5905 -38 -5899 38
rect -5945 -50 -5899 -38
rect -5287 38 -5241 50
rect -5287 -38 -5281 38
rect -5247 -38 -5241 38
rect -5287 -50 -5241 -38
rect -4629 38 -4583 50
rect -4629 -38 -4623 38
rect -4589 -38 -4583 38
rect -4629 -50 -4583 -38
rect -3971 38 -3925 50
rect -3971 -38 -3965 38
rect -3931 -38 -3925 38
rect -3971 -50 -3925 -38
rect -3313 38 -3267 50
rect -3313 -38 -3307 38
rect -3273 -38 -3267 38
rect -3313 -50 -3267 -38
rect -2655 38 -2609 50
rect -2655 -38 -2649 38
rect -2615 -38 -2609 38
rect -2655 -50 -2609 -38
rect -1997 38 -1951 50
rect -1997 -38 -1991 38
rect -1957 -38 -1951 38
rect -1997 -50 -1951 -38
rect -1339 38 -1293 50
rect -1339 -38 -1333 38
rect -1299 -38 -1293 38
rect -1339 -50 -1293 -38
rect -681 38 -635 50
rect -681 -38 -675 38
rect -641 -38 -635 38
rect -681 -50 -635 -38
rect -23 38 23 50
rect -23 -38 -17 38
rect 17 -38 23 38
rect -23 -50 23 -38
rect 635 38 681 50
rect 635 -38 641 38
rect 675 -38 681 38
rect 635 -50 681 -38
rect 1293 38 1339 50
rect 1293 -38 1299 38
rect 1333 -38 1339 38
rect 1293 -50 1339 -38
rect 1951 38 1997 50
rect 1951 -38 1957 38
rect 1991 -38 1997 38
rect 1951 -50 1997 -38
rect 2609 38 2655 50
rect 2609 -38 2615 38
rect 2649 -38 2655 38
rect 2609 -50 2655 -38
rect 3267 38 3313 50
rect 3267 -38 3273 38
rect 3307 -38 3313 38
rect 3267 -50 3313 -38
rect 3925 38 3971 50
rect 3925 -38 3931 38
rect 3965 -38 3971 38
rect 3925 -50 3971 -38
rect 4583 38 4629 50
rect 4583 -38 4589 38
rect 4623 -38 4629 38
rect 4583 -50 4629 -38
rect 5241 38 5287 50
rect 5241 -38 5247 38
rect 5281 -38 5287 38
rect 5241 -50 5287 -38
rect 5899 38 5945 50
rect 5899 -38 5905 38
rect 5939 -38 5945 38
rect 5899 -50 5945 -38
rect 6557 38 6603 50
rect 6557 -38 6563 38
rect 6597 -38 6603 38
rect 6557 -50 6603 -38
rect -6547 -88 -5955 -82
rect -6547 -122 -6535 -88
rect -5967 -122 -5955 -88
rect -6547 -128 -5955 -122
rect -5889 -88 -5297 -82
rect -5889 -122 -5877 -88
rect -5309 -122 -5297 -88
rect -5889 -128 -5297 -122
rect -5231 -88 -4639 -82
rect -5231 -122 -5219 -88
rect -4651 -122 -4639 -88
rect -5231 -128 -4639 -122
rect -4573 -88 -3981 -82
rect -4573 -122 -4561 -88
rect -3993 -122 -3981 -88
rect -4573 -128 -3981 -122
rect -3915 -88 -3323 -82
rect -3915 -122 -3903 -88
rect -3335 -122 -3323 -88
rect -3915 -128 -3323 -122
rect -3257 -88 -2665 -82
rect -3257 -122 -3245 -88
rect -2677 -122 -2665 -88
rect -3257 -128 -2665 -122
rect -2599 -88 -2007 -82
rect -2599 -122 -2587 -88
rect -2019 -122 -2007 -88
rect -2599 -128 -2007 -122
rect -1941 -88 -1349 -82
rect -1941 -122 -1929 -88
rect -1361 -122 -1349 -88
rect -1941 -128 -1349 -122
rect -1283 -88 -691 -82
rect -1283 -122 -1271 -88
rect -703 -122 -691 -88
rect -1283 -128 -691 -122
rect -625 -88 -33 -82
rect -625 -122 -613 -88
rect -45 -122 -33 -88
rect -625 -128 -33 -122
rect 33 -88 625 -82
rect 33 -122 45 -88
rect 613 -122 625 -88
rect 33 -128 625 -122
rect 691 -88 1283 -82
rect 691 -122 703 -88
rect 1271 -122 1283 -88
rect 691 -128 1283 -122
rect 1349 -88 1941 -82
rect 1349 -122 1361 -88
rect 1929 -122 1941 -88
rect 1349 -128 1941 -122
rect 2007 -88 2599 -82
rect 2007 -122 2019 -88
rect 2587 -122 2599 -88
rect 2007 -128 2599 -122
rect 2665 -88 3257 -82
rect 2665 -122 2677 -88
rect 3245 -122 3257 -88
rect 2665 -128 3257 -122
rect 3323 -88 3915 -82
rect 3323 -122 3335 -88
rect 3903 -122 3915 -88
rect 3323 -128 3915 -122
rect 3981 -88 4573 -82
rect 3981 -122 3993 -88
rect 4561 -122 4573 -88
rect 3981 -128 4573 -122
rect 4639 -88 5231 -82
rect 4639 -122 4651 -88
rect 5219 -122 5231 -88
rect 4639 -128 5231 -122
rect 5297 -88 5889 -82
rect 5297 -122 5309 -88
rect 5877 -122 5889 -88
rect 5297 -128 5889 -122
rect 5955 -88 6547 -82
rect 5955 -122 5967 -88
rect 6535 -122 6547 -88
rect 5955 -128 6547 -122
<< properties >>
string FIXED_BBOX -6694 -207 6694 207
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 0.5 l 3.0 m 1 nf 20 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
