magic
tech sky130A
magscale 1 2
timestamp 1695195202
<< nwell >>
rect -1154 -3219 1154 3219
<< pmoslvt >>
rect -958 -3000 -358 3000
rect -300 -3000 300 3000
rect 358 -3000 958 3000
<< pdiff >>
rect -1016 2988 -958 3000
rect -1016 -2988 -1004 2988
rect -970 -2988 -958 2988
rect -1016 -3000 -958 -2988
rect -358 2988 -300 3000
rect -358 -2988 -346 2988
rect -312 -2988 -300 2988
rect -358 -3000 -300 -2988
rect 300 2988 358 3000
rect 300 -2988 312 2988
rect 346 -2988 358 2988
rect 300 -3000 358 -2988
rect 958 2988 1016 3000
rect 958 -2988 970 2988
rect 1004 -2988 1016 2988
rect 958 -3000 1016 -2988
<< pdiffc >>
rect -1004 -2988 -970 2988
rect -346 -2988 -312 2988
rect 312 -2988 346 2988
rect 970 -2988 1004 2988
<< nsubdiff >>
rect -1118 3149 -1022 3183
rect 1022 3149 1118 3183
rect -1118 3087 -1084 3149
rect 1084 3087 1118 3149
rect -1118 -3149 -1084 -3087
rect 1084 -3149 1118 -3087
rect -1118 -3183 -1022 -3149
rect 1022 -3183 1118 -3149
<< nsubdiffcont >>
rect -1022 3149 1022 3183
rect -1118 -3087 -1084 3087
rect 1084 -3087 1118 3087
rect -1022 -3183 1022 -3149
<< poly >>
rect -958 3081 -358 3097
rect -958 3047 -942 3081
rect -374 3047 -358 3081
rect -958 3000 -358 3047
rect -300 3081 300 3097
rect -300 3047 -284 3081
rect 284 3047 300 3081
rect -300 3000 300 3047
rect 358 3081 958 3097
rect 358 3047 374 3081
rect 942 3047 958 3081
rect 358 3000 958 3047
rect -958 -3047 -358 -3000
rect -958 -3081 -942 -3047
rect -374 -3081 -358 -3047
rect -958 -3097 -358 -3081
rect -300 -3047 300 -3000
rect -300 -3081 -284 -3047
rect 284 -3081 300 -3047
rect -300 -3097 300 -3081
rect 358 -3047 958 -3000
rect 358 -3081 374 -3047
rect 942 -3081 958 -3047
rect 358 -3097 958 -3081
<< polycont >>
rect -942 3047 -374 3081
rect -284 3047 284 3081
rect 374 3047 942 3081
rect -942 -3081 -374 -3047
rect -284 -3081 284 -3047
rect 374 -3081 942 -3047
<< locali >>
rect -1118 3149 -1022 3183
rect 1022 3149 1118 3183
rect -1118 3087 -1084 3149
rect 1084 3087 1118 3149
rect -958 3047 -942 3081
rect -374 3047 -358 3081
rect -300 3047 -284 3081
rect 284 3047 300 3081
rect 358 3047 374 3081
rect 942 3047 958 3081
rect -1004 2988 -970 3004
rect -1004 -3004 -970 -2988
rect -346 2988 -312 3004
rect -346 -3004 -312 -2988
rect 312 2988 346 3004
rect 312 -3004 346 -2988
rect 970 2988 1004 3004
rect 970 -3004 1004 -2988
rect -958 -3081 -942 -3047
rect -374 -3081 -358 -3047
rect -300 -3081 -284 -3047
rect 284 -3081 300 -3047
rect 358 -3081 374 -3047
rect 942 -3081 958 -3047
rect -1118 -3149 -1084 -3087
rect 1084 -3149 1118 -3087
rect -1118 -3183 -1022 -3149
rect 1022 -3183 1118 -3149
<< viali >>
rect -942 3047 -374 3081
rect -284 3047 284 3081
rect 374 3047 942 3081
rect -1004 -2988 -970 2988
rect -346 -2988 -312 2988
rect 312 -2988 346 2988
rect 970 -2988 1004 2988
rect -942 -3081 -374 -3047
rect -284 -3081 284 -3047
rect 374 -3081 942 -3047
<< metal1 >>
rect -954 3081 -362 3087
rect -954 3047 -942 3081
rect -374 3047 -362 3081
rect -954 3041 -362 3047
rect -296 3081 296 3087
rect -296 3047 -284 3081
rect 284 3047 296 3081
rect -296 3041 296 3047
rect 362 3081 954 3087
rect 362 3047 374 3081
rect 942 3047 954 3081
rect 362 3041 954 3047
rect -1010 2988 -964 3000
rect -1010 -2988 -1004 2988
rect -970 -2988 -964 2988
rect -1010 -3000 -964 -2988
rect -352 2988 -306 3000
rect -352 -2988 -346 2988
rect -312 -2988 -306 2988
rect -352 -3000 -306 -2988
rect 306 2988 352 3000
rect 306 -2988 312 2988
rect 346 -2988 352 2988
rect 306 -3000 352 -2988
rect 964 2988 1010 3000
rect 964 -2988 970 2988
rect 1004 -2988 1010 2988
rect 964 -3000 1010 -2988
rect -954 -3047 -362 -3041
rect -954 -3081 -942 -3047
rect -374 -3081 -362 -3047
rect -954 -3087 -362 -3081
rect -296 -3047 296 -3041
rect -296 -3081 -284 -3047
rect 284 -3081 296 -3047
rect -296 -3087 296 -3081
rect 362 -3047 954 -3041
rect 362 -3081 374 -3047
rect 942 -3081 954 -3047
rect 362 -3087 954 -3081
<< properties >>
string FIXED_BBOX -1101 -3166 1101 3166
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 30.0 l 3.0 m 1 nf 3 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
