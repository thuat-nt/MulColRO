magic
tech sky130A
timestamp 1695441144
<< pwell >>
rect -906 -905 906 905
<< nmoslvt >>
rect -808 -800 -508 800
rect -479 -800 -179 800
rect -150 -800 150 800
rect 179 -800 479 800
rect 508 -800 808 800
<< ndiff >>
rect -837 794 -808 800
rect -837 -794 -831 794
rect -814 -794 -808 794
rect -837 -800 -808 -794
rect -508 794 -479 800
rect -508 -794 -502 794
rect -485 -794 -479 794
rect -508 -800 -479 -794
rect -179 794 -150 800
rect -179 -794 -173 794
rect -156 -794 -150 794
rect -179 -800 -150 -794
rect 150 794 179 800
rect 150 -794 156 794
rect 173 -794 179 794
rect 150 -800 179 -794
rect 479 794 508 800
rect 479 -794 485 794
rect 502 -794 508 794
rect 479 -800 508 -794
rect 808 794 837 800
rect 808 -794 814 794
rect 831 -794 837 794
rect 808 -800 837 -794
<< ndiffc >>
rect -831 -794 -814 794
rect -502 -794 -485 794
rect -173 -794 -156 794
rect 156 -794 173 794
rect 485 -794 502 794
rect 814 -794 831 794
<< psubdiff >>
rect -888 870 -840 887
rect 840 870 888 887
rect -888 839 -871 870
rect 871 839 888 870
rect -888 -870 -871 -839
rect 871 -870 888 -839
rect -888 -887 -840 -870
rect 840 -887 888 -870
<< psubdiffcont >>
rect -840 870 840 887
rect -888 -839 -871 839
rect 871 -839 888 839
rect -840 -887 840 -870
<< poly >>
rect -808 836 -508 844
rect -808 819 -800 836
rect -516 819 -508 836
rect -808 800 -508 819
rect -479 836 -179 844
rect -479 819 -471 836
rect -187 819 -179 836
rect -479 800 -179 819
rect -150 836 150 844
rect -150 819 -142 836
rect 142 819 150 836
rect -150 800 150 819
rect 179 836 479 844
rect 179 819 187 836
rect 471 819 479 836
rect 179 800 479 819
rect 508 836 808 844
rect 508 819 516 836
rect 800 819 808 836
rect 508 800 808 819
rect -808 -819 -508 -800
rect -808 -836 -800 -819
rect -516 -836 -508 -819
rect -808 -844 -508 -836
rect -479 -819 -179 -800
rect -479 -836 -471 -819
rect -187 -836 -179 -819
rect -479 -844 -179 -836
rect -150 -819 150 -800
rect -150 -836 -142 -819
rect 142 -836 150 -819
rect -150 -844 150 -836
rect 179 -819 479 -800
rect 179 -836 187 -819
rect 471 -836 479 -819
rect 179 -844 479 -836
rect 508 -819 808 -800
rect 508 -836 516 -819
rect 800 -836 808 -819
rect 508 -844 808 -836
<< polycont >>
rect -800 819 -516 836
rect -471 819 -187 836
rect -142 819 142 836
rect 187 819 471 836
rect 516 819 800 836
rect -800 -836 -516 -819
rect -471 -836 -187 -819
rect -142 -836 142 -819
rect 187 -836 471 -819
rect 516 -836 800 -819
<< locali >>
rect -888 870 -840 887
rect 840 870 888 887
rect -888 839 -871 870
rect 871 839 888 870
rect -808 819 -800 836
rect -516 819 -508 836
rect -479 819 -471 836
rect -187 819 -179 836
rect -150 819 -142 836
rect 142 819 150 836
rect 179 819 187 836
rect 471 819 479 836
rect 508 819 516 836
rect 800 819 808 836
rect -831 794 -814 802
rect -831 -802 -814 -794
rect -502 794 -485 802
rect -502 -802 -485 -794
rect -173 794 -156 802
rect -173 -802 -156 -794
rect 156 794 173 802
rect 156 -802 173 -794
rect 485 794 502 802
rect 485 -802 502 -794
rect 814 794 831 802
rect 814 -802 831 -794
rect -808 -836 -800 -819
rect -516 -836 -508 -819
rect -479 -836 -471 -819
rect -187 -836 -179 -819
rect -150 -836 -142 -819
rect 142 -836 150 -819
rect 179 -836 187 -819
rect 471 -836 479 -819
rect 508 -836 516 -819
rect 800 -836 808 -819
rect -888 -870 -871 -839
rect 871 -870 888 -839
rect -888 -887 -840 -870
rect 840 -887 888 -870
<< viali >>
rect -800 819 -516 836
rect -471 819 -187 836
rect -142 819 142 836
rect 187 819 471 836
rect 516 819 800 836
rect -831 -794 -814 794
rect -502 -794 -485 794
rect -173 -794 -156 794
rect 156 -794 173 794
rect 485 -794 502 794
rect 814 -794 831 794
rect -800 -836 -516 -819
rect -471 -836 -187 -819
rect -142 -836 142 -819
rect 187 -836 471 -819
rect 516 -836 800 -819
<< metal1 >>
rect -806 836 -510 839
rect -806 819 -800 836
rect -516 819 -510 836
rect -806 816 -510 819
rect -477 836 -181 839
rect -477 819 -471 836
rect -187 819 -181 836
rect -477 816 -181 819
rect -148 836 148 839
rect -148 819 -142 836
rect 142 819 148 836
rect -148 816 148 819
rect 181 836 477 839
rect 181 819 187 836
rect 471 819 477 836
rect 181 816 477 819
rect 510 836 806 839
rect 510 819 516 836
rect 800 819 806 836
rect 510 816 806 819
rect -834 794 -811 800
rect -834 -794 -831 794
rect -814 -794 -811 794
rect -834 -800 -811 -794
rect -505 794 -482 800
rect -505 -794 -502 794
rect -485 -794 -482 794
rect -505 -800 -482 -794
rect -176 794 -153 800
rect -176 -794 -173 794
rect -156 -794 -153 794
rect -176 -800 -153 -794
rect 153 794 176 800
rect 153 -794 156 794
rect 173 -794 176 794
rect 153 -800 176 -794
rect 482 794 505 800
rect 482 -794 485 794
rect 502 -794 505 794
rect 482 -800 505 -794
rect 811 794 834 800
rect 811 -794 814 794
rect 831 -794 834 794
rect 811 -800 834 -794
rect -806 -819 -510 -816
rect -806 -836 -800 -819
rect -516 -836 -510 -819
rect -806 -839 -510 -836
rect -477 -819 -181 -816
rect -477 -836 -471 -819
rect -187 -836 -181 -819
rect -477 -839 -181 -836
rect -148 -819 148 -816
rect -148 -836 -142 -819
rect 142 -836 148 -819
rect -148 -839 148 -836
rect 181 -819 477 -816
rect 181 -836 187 -819
rect 471 -836 477 -819
rect 181 -839 477 -836
rect 510 -819 806 -816
rect 510 -836 516 -819
rect 800 -836 806 -819
rect 510 -839 806 -836
<< labels >>
rlabel locali -831 794 -814 802 1 D
rlabel poly -808 800 -508 819 1 G
rlabel locali -502 794 -485 802 1 S
rlabel psubdiffcont -840 -887 840 -870 1 B
<< properties >>
string FIXED_BBOX -879 -878 879 878
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 16.0 l 3.0 m 1 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
