magic
tech sky130A
magscale 1 2
timestamp 1698976668
<< locali >>
rect 472 946 1284 1034
rect 476 892 614 946
rect 476 810 528 892
rect 476 768 614 810
rect 494 -420 1232 -360
rect 494 -530 542 -420
rect 650 -530 1232 -420
rect 494 -578 1232 -530
<< viali >>
rect 528 810 614 892
rect 542 -530 650 -420
<< metal1 >>
rect 476 892 662 990
rect 476 814 528 892
rect 474 810 528 814
rect 614 814 662 892
rect 1020 848 1096 914
rect 614 810 1012 814
rect 1310 810 1412 818
rect 474 708 1012 810
rect 474 706 996 708
rect 474 656 1004 706
rect 474 414 1012 656
rect 1100 428 1412 810
rect 994 360 1114 378
rect 994 296 1010 360
rect 1100 296 1114 360
rect 994 282 1114 296
rect 512 232 712 274
rect 512 156 614 232
rect 686 216 712 232
rect 1308 256 1412 428
rect 1668 256 1868 262
rect 686 156 714 216
rect 512 130 714 156
rect 512 74 712 130
rect 1006 78 1112 98
rect 1006 26 1030 78
rect 1086 26 1112 78
rect 1006 8 1112 26
rect 1308 70 1868 256
rect 1308 -34 1412 70
rect 1668 62 1868 70
rect 492 -212 1004 -34
rect 1106 -36 1412 -34
rect 1106 -210 1410 -36
rect 492 -420 700 -212
rect 1308 -220 1410 -210
rect 1020 -314 1086 -256
rect 492 -530 542 -420
rect 650 -530 700 -420
rect 492 -578 700 -530
<< via1 >>
rect 1010 296 1100 360
rect 614 156 686 232
rect 1030 26 1086 78
<< metal2 >>
rect 1024 380 1088 408
rect 984 360 1138 380
rect 984 296 1010 360
rect 1100 296 1138 360
rect 984 278 1138 296
rect 1024 250 1088 278
rect 584 232 1088 250
rect 584 156 614 232
rect 686 156 1088 232
rect 584 142 1088 156
rect 1024 88 1088 142
rect 1018 78 1098 88
rect 1018 26 1030 78
rect 1086 26 1098 78
rect 1018 14 1098 26
use sky130_fd_pr__nfet_01v8_lvt_6LX62X  XM1
timestamp 1696652587
transform 1 0 1055 0 1 -122
box -231 -310 231 310
use sky130_fd_pr__pfet_01v8_lvt_4QFWD3  XM10
timestamp 1696652587
transform 1 0 1055 0 1 617
box -231 -419 231 419
<< labels >>
flabel metal1 512 74 712 274 0 FreeSans 256 0 0 0 in
port 1 nsew
flabel metal1 1668 62 1868 262 0 FreeSans 256 0 0 0 out
port 0 nsew
rlabel locali 472 946 1284 1034 1 VDD
port 4 nsew
rlabel locali 494 -578 1232 -360 1 VSS
port 5 nsew
<< end >>
