magic
tech sky130A
magscale 1 2
timestamp 1696348358
<< pwell >>
rect 10708 4824 10888 4998
<< nmoslvt >>
rect 10708 4824 10888 4998
<< locali >>
rect 7334 8992 18966 9014
rect 7334 8778 14840 8992
rect 15112 8778 18966 8992
rect 7334 8482 18966 8778
rect 6154 7224 11066 7710
rect 6154 7210 14704 7224
rect 6154 6780 15260 7210
rect 6164 5406 6532 6780
rect 11268 5404 11636 6780
rect 6476 3696 7476 3942
rect 6476 3424 6788 3696
rect 7146 3424 7476 3696
rect 6476 1756 7476 3424
rect 7674 3692 8674 3930
rect 7674 3454 7972 3692
rect 8354 3454 8674 3692
rect 7674 1756 8674 3454
rect 8968 3290 9980 3344
rect 8968 3136 9340 3290
rect 9610 3136 9980 3290
rect 8968 1756 9980 3136
rect 10140 3258 11152 3348
rect 10140 3080 10484 3258
rect 10818 3080 11152 3258
rect 10140 1756 11152 3080
rect 6276 1644 15318 1756
rect 6276 1370 12950 1644
rect 13302 1370 15318 1644
rect 6276 1244 15318 1370
<< viali >>
rect 14840 8778 15112 8992
rect 6788 3424 7146 3696
rect 7972 3454 8354 3692
rect 9340 3136 9610 3290
rect 10484 3080 10818 3258
rect 12950 1370 13302 1644
<< metal1 >>
rect 14824 8998 15122 9002
rect 14824 8992 15124 8998
rect 14824 8778 14840 8992
rect 15112 8778 15124 8992
rect 14824 8772 15124 8778
rect 14824 8768 15122 8772
rect 7118 8164 7318 8178
rect 7118 7994 7132 8164
rect 7300 7994 7318 8164
rect 7718 8096 8220 8432
rect 8254 8344 8350 8346
rect 8254 8168 8272 8344
rect 8336 8168 8350 8344
rect 8254 8154 8350 8168
rect 7718 8042 7738 8096
rect 8208 8042 8220 8096
rect 7118 7978 7318 7994
rect 7502 7994 7666 8002
rect 7502 7846 7514 7994
rect 7662 7846 7672 7994
rect 7502 7840 7666 7846
rect 7718 7772 8220 8042
rect 8380 8094 8882 8432
rect 8380 8032 8466 8094
rect 8762 8032 8882 8094
rect 8380 7772 8882 8032
rect 9038 8094 9540 8432
rect 9580 8326 9664 8348
rect 9580 8184 9590 8326
rect 9656 8184 9664 8326
rect 9580 8162 9664 8184
rect 9038 8032 9126 8094
rect 9422 8032 9540 8094
rect 8928 7988 9000 7998
rect 8924 7858 8934 7988
rect 8994 7858 9004 7988
rect 8928 7856 9000 7858
rect 9038 7772 9540 8032
rect 9694 8094 10196 8432
rect 9694 8032 9810 8094
rect 10106 8032 10196 8094
rect 9694 7772 10196 8032
rect 11240 8002 11738 8436
rect 11772 8346 11862 8350
rect 11772 8096 11788 8346
rect 11842 8096 11862 8346
rect 11772 8082 11862 8096
rect 10248 7988 10310 7998
rect 10242 7862 10252 7988
rect 10304 7862 10314 7988
rect 10248 7858 10310 7862
rect 11240 7848 11358 8002
rect 11602 7848 11738 8002
rect 11080 7580 11206 7598
rect 11080 7368 11100 7580
rect 11192 7368 11206 7580
rect 11080 7358 11206 7368
rect 11240 7274 11738 7848
rect 11892 7998 12390 8436
rect 11892 7852 12040 7998
rect 12290 7852 12390 7998
rect 11892 7274 12390 7852
rect 13326 8002 13824 8434
rect 13862 8344 13950 8348
rect 13862 8186 13878 8344
rect 13934 8186 13950 8344
rect 13862 8172 13950 8186
rect 13326 7848 13452 8002
rect 13696 7848 13824 8002
rect 12422 7676 12530 7706
rect 12422 7368 12432 7676
rect 12514 7368 12530 7676
rect 12422 7358 12530 7368
rect 13178 7596 13294 7614
rect 13178 7362 13188 7596
rect 13280 7362 13294 7596
rect 13178 7358 13294 7362
rect 13326 7272 13824 7848
rect 13980 7998 14478 8434
rect 13980 7852 14100 7998
rect 14350 7852 14478 7998
rect 13980 7272 14478 7852
rect 14518 7610 14608 7668
rect 14516 7364 14526 7610
rect 14600 7364 14610 7610
rect 14518 7356 14608 7364
rect 15432 7012 15928 8436
rect 15962 8348 16054 8350
rect 15962 8188 15978 8348
rect 16038 8188 16054 8348
rect 15962 8164 16054 8188
rect 15432 6848 15488 7012
rect 15876 6848 15928 7012
rect 6068 6304 6268 6320
rect 6068 6134 6084 6304
rect 6252 6134 6268 6304
rect 6068 6120 6268 6134
rect 6710 6270 7206 6724
rect 7236 6636 7330 6640
rect 7236 6372 7246 6636
rect 7320 6372 7330 6636
rect 7236 6354 7330 6372
rect 6710 6166 6760 6270
rect 7174 6166 7206 6270
rect 6570 5886 6672 5926
rect 6570 5654 6588 5886
rect 6664 5654 6674 5886
rect 6570 5648 6672 5654
rect 6710 5562 7206 6166
rect 7362 6272 7858 6724
rect 7362 6166 7496 6272
rect 7782 6166 7858 6272
rect 7362 5562 7858 6166
rect 8022 6274 8518 6724
rect 8562 6628 8652 6640
rect 8558 6440 8568 6628
rect 8646 6440 8656 6628
rect 8562 6432 8652 6440
rect 8022 6168 8154 6274
rect 8440 6168 8518 6274
rect 7888 5918 7990 5926
rect 7888 5666 7902 5918
rect 7982 5666 7992 5918
rect 7888 5654 7990 5666
rect 8022 5562 8518 6168
rect 9288 6254 9780 6730
rect 9812 6642 9910 6644
rect 9812 6438 9824 6642
rect 9900 6438 9910 6642
rect 9812 6434 9910 6438
rect 9288 6186 9302 6254
rect 9756 6186 9780 6254
rect 9288 6038 9780 6186
rect 9150 5930 9254 5952
rect 9150 5666 9160 5930
rect 9242 5666 9254 5930
rect 9150 5656 9254 5666
rect 9284 5568 9780 6038
rect 9944 6254 10440 6730
rect 9944 6192 10046 6254
rect 10342 6192 10440 6254
rect 9944 5568 10440 6192
rect 10606 6254 11102 6730
rect 11136 6636 11218 6644
rect 11134 6452 11144 6636
rect 11206 6452 11218 6636
rect 11136 6440 11218 6452
rect 10606 6192 10708 6254
rect 11004 6192 11102 6254
rect 10468 5920 10574 5932
rect 10468 5656 10474 5920
rect 10564 5656 10574 5920
rect 10468 5650 10574 5656
rect 10606 5568 11102 6192
rect 11534 6296 11734 6314
rect 11534 6126 11546 6296
rect 11714 6126 11734 6296
rect 11534 6114 11734 6126
rect 6572 5060 6684 5064
rect 6572 4898 6598 5060
rect 6676 4898 6686 5060
rect 6572 4878 6684 4898
rect 6734 4646 7230 5138
rect 7762 5058 7882 5062
rect 7762 4790 7776 5058
rect 7862 4790 7882 5058
rect 7762 4780 7882 4790
rect 6734 4522 6774 4646
rect 7202 4522 7230 4646
rect 6734 3994 7230 4522
rect 7918 4642 8414 5138
rect 9084 5068 9188 5070
rect 9084 4856 9098 5068
rect 9176 4856 9188 5068
rect 9084 4840 9188 4856
rect 7918 4518 7948 4642
rect 8376 4518 8414 4642
rect 7268 4322 7392 4356
rect 7266 4082 7276 4322
rect 7380 4082 7392 4322
rect 7268 4074 7392 4082
rect 7918 3994 8414 4518
rect 9226 4412 9730 5146
rect 10254 5074 10358 5076
rect 10254 4882 10270 5074
rect 10346 4882 10358 5074
rect 10254 4862 10358 4882
rect 8444 4386 8578 4400
rect 8444 4118 8470 4386
rect 8556 4118 8578 4386
rect 8444 4090 8578 4118
rect 9226 4336 9412 4412
rect 9562 4336 9730 4412
rect 6756 3696 7174 3726
rect 6756 3424 6788 3696
rect 7146 3424 7174 3696
rect 6756 3406 7174 3424
rect 7908 3692 8402 3756
rect 7908 3454 7972 3692
rect 8354 3454 8402 3692
rect 7908 3418 8402 3454
rect 9226 3402 9730 4336
rect 10386 4416 10890 5154
rect 11420 4770 11526 5080
rect 11420 4684 11428 4770
rect 11518 4684 11526 4770
rect 11420 4674 11526 4684
rect 10386 4348 10626 4416
rect 10748 4348 10890 4416
rect 9760 3664 9884 3686
rect 9760 3482 9770 3664
rect 9856 3482 9884 3664
rect 9760 3480 9884 3482
rect 10386 3410 10890 4348
rect 11556 3778 12054 5158
rect 10922 3692 11046 3742
rect 10922 3492 10936 3692
rect 11026 3492 11046 3692
rect 10922 3486 11046 3492
rect 11556 3654 11828 3778
rect 11980 3654 12054 3778
rect 9318 3290 9632 3304
rect 9318 3136 9340 3290
rect 9610 3136 9632 3290
rect 9318 3122 9632 3136
rect 10466 3258 10832 3280
rect 10466 3080 10484 3258
rect 10818 3080 10832 3258
rect 10466 3054 10832 3080
rect 11556 1814 12054 3654
rect 12206 3782 12704 5158
rect 12738 5046 12840 5062
rect 12738 4748 12752 5046
rect 12830 4748 12840 5046
rect 12738 4734 12840 4748
rect 12206 3668 12366 3782
rect 12558 3668 12704 3782
rect 12084 2104 12176 2152
rect 12084 1892 12094 2104
rect 12168 1892 12176 2104
rect 12084 1890 12176 1892
rect 12206 1814 12704 3668
rect 12870 3782 13368 5158
rect 12870 3668 13050 3782
rect 13242 3668 13368 3782
rect 12870 1814 13368 3668
rect 13528 3774 14026 5158
rect 14056 5078 14158 5080
rect 14056 4792 14062 5078
rect 14148 4792 14158 5078
rect 14056 4782 14158 4792
rect 13528 3660 13678 3774
rect 13870 3660 14026 3774
rect 13398 2126 13500 2192
rect 13398 1896 13408 2126
rect 13488 1896 13500 2126
rect 13398 1890 13500 1896
rect 13528 1814 14026 3660
rect 14192 3790 14690 5158
rect 15286 4708 15396 4760
rect 15286 4366 15294 4708
rect 15384 4366 15396 4708
rect 15286 4352 15396 4366
rect 15432 4274 15928 6848
rect 16082 6996 16578 8436
rect 16082 6882 16262 6996
rect 16454 6882 16578 6996
rect 16082 4274 16578 6882
rect 16738 7002 17234 8436
rect 17272 8344 17374 8366
rect 17272 8156 17282 8344
rect 17360 8156 17374 8344
rect 17272 8144 17374 8156
rect 16738 6888 16906 7002
rect 17098 6888 17234 7002
rect 16612 4560 16706 4570
rect 16612 4364 16622 4560
rect 16694 4364 16706 4560
rect 16612 4358 16706 4364
rect 16738 4274 17234 6888
rect 17410 6996 17906 8436
rect 17410 6882 17562 6996
rect 17754 6882 17906 6996
rect 17410 4274 17906 6882
rect 18060 6986 18556 8436
rect 18590 8354 18686 8364
rect 18590 8176 18600 8354
rect 18674 8176 18686 8354
rect 18590 8168 18686 8176
rect 18060 6872 18202 6986
rect 18394 6872 18556 6986
rect 17936 4556 18032 4568
rect 17936 4364 17946 4556
rect 18020 4364 18032 4556
rect 17936 4360 18032 4364
rect 18060 4274 18556 6872
rect 14192 3676 14300 3790
rect 14492 3676 14690 3790
rect 14192 1814 14690 3676
rect 16658 2568 16858 2576
rect 16658 2384 16692 2568
rect 16844 2384 16858 2568
rect 16658 2376 16858 2384
rect 14720 2182 14836 2200
rect 14720 1898 14730 2182
rect 14818 1898 14836 2182
rect 14720 1894 14836 1898
rect 12922 1644 13332 1672
rect 12922 1370 12950 1644
rect 13302 1370 13332 1644
rect 12922 1348 13332 1370
<< via1 >>
rect 14840 8778 15112 8992
rect 7132 7994 7300 8164
rect 8272 8168 8336 8344
rect 7738 8042 8208 8096
rect 7514 7846 7662 7994
rect 8466 8032 8762 8094
rect 9590 8184 9656 8326
rect 9126 8032 9422 8094
rect 8934 7858 8994 7988
rect 9810 8032 10106 8094
rect 11788 8096 11842 8346
rect 10252 7862 10304 7988
rect 11358 7848 11602 8002
rect 11100 7368 11192 7580
rect 12040 7852 12290 7998
rect 13878 8186 13934 8344
rect 13452 7848 13696 8002
rect 12432 7368 12514 7676
rect 13188 7362 13280 7596
rect 14100 7852 14350 7998
rect 14526 7364 14600 7610
rect 15978 8188 16038 8348
rect 15488 6848 15876 7012
rect 6084 6134 6252 6304
rect 7246 6372 7320 6636
rect 6760 6166 7174 6270
rect 6588 5654 6664 5886
rect 7496 6166 7782 6272
rect 8568 6440 8646 6628
rect 8154 6168 8440 6274
rect 7902 5666 7982 5918
rect 9824 6438 9900 6642
rect 9302 6186 9756 6254
rect 9160 5666 9242 5930
rect 10046 6192 10342 6254
rect 11144 6452 11206 6636
rect 10708 6192 11004 6254
rect 10474 5656 10564 5920
rect 11546 6126 11714 6296
rect 6598 4898 6676 5060
rect 7776 4790 7862 5058
rect 6774 4522 7202 4646
rect 9098 4856 9176 5068
rect 7948 4518 8376 4642
rect 7276 4082 7380 4322
rect 10270 4882 10346 5074
rect 8470 4118 8556 4386
rect 9412 4336 9562 4412
rect 6788 3424 7146 3696
rect 7972 3454 8354 3692
rect 11428 4684 11518 4770
rect 10626 4348 10748 4416
rect 9770 3482 9856 3664
rect 10936 3492 11026 3692
rect 11828 3654 11980 3778
rect 9340 3136 9610 3290
rect 10484 3080 10818 3258
rect 12752 4748 12830 5046
rect 12366 3668 12558 3782
rect 12094 1892 12168 2104
rect 13050 3668 13242 3782
rect 14062 4792 14148 5078
rect 13678 3660 13870 3774
rect 13408 1896 13488 2126
rect 15294 4366 15384 4708
rect 16262 6882 16454 6996
rect 17282 8156 17360 8344
rect 16906 6888 17098 7002
rect 16622 4364 16694 4560
rect 17562 6882 17754 6996
rect 18600 8176 18674 8354
rect 18202 6872 18394 6986
rect 17946 4364 18020 4556
rect 14300 3676 14492 3790
rect 16692 2384 16844 2568
rect 14730 1898 14818 2182
rect 12950 1370 13302 1644
<< metal2 >>
rect 14806 8992 15136 9012
rect 14806 8778 14840 8992
rect 15112 8778 15136 8992
rect 14806 8436 15136 8778
rect 7480 8354 18806 8436
rect 7480 8348 18600 8354
rect 7480 8346 15978 8348
rect 7480 8344 11788 8346
rect 7132 8164 7300 8174
rect 7480 8168 8272 8344
rect 8336 8326 11788 8344
rect 8336 8184 9590 8326
rect 9656 8184 11788 8326
rect 8336 8168 11788 8184
rect 7480 8134 11788 8168
rect 7738 8096 8208 8106
rect 11842 8344 15978 8346
rect 11842 8186 13878 8344
rect 13934 8188 15978 8344
rect 16038 8344 18600 8348
rect 16038 8188 17282 8344
rect 13934 8186 17282 8188
rect 11842 8156 17282 8186
rect 17360 8176 18600 8344
rect 18674 8176 18806 8354
rect 17360 8156 18806 8176
rect 11842 8134 18806 8156
rect 14806 8130 15136 8134
rect 7300 8042 7738 8096
rect 8208 8094 10458 8096
rect 8208 8042 8466 8094
rect 7300 8032 8466 8042
rect 8762 8032 9126 8094
rect 9422 8032 9810 8094
rect 10106 8032 10458 8094
rect 11788 8086 11842 8096
rect 7132 7984 7300 7994
rect 7480 7994 10446 8004
rect 7480 7846 7514 7994
rect 7662 7988 10446 7994
rect 7662 7858 8934 7988
rect 8994 7862 10252 7988
rect 10304 7862 10446 7988
rect 8994 7858 10446 7862
rect 7662 7846 10446 7858
rect 7480 7770 10446 7846
rect 10992 8002 14736 8014
rect 10992 7848 11358 8002
rect 11602 7998 13452 8002
rect 11602 7852 12040 7998
rect 12290 7852 13452 7998
rect 11602 7848 13452 7852
rect 13696 7998 14736 8002
rect 13696 7852 14100 7998
rect 14350 7852 14736 7998
rect 13696 7848 14736 7852
rect 10992 7836 14736 7848
rect 8794 6730 8998 7770
rect 10992 7676 12642 7758
rect 10992 7580 12432 7676
rect 10992 7368 11100 7580
rect 11192 7504 12432 7580
rect 11326 7368 12432 7504
rect 12514 7644 12642 7676
rect 12768 7644 12960 7836
rect 12514 7470 12960 7644
rect 13078 7610 14728 7756
rect 13078 7596 14526 7610
rect 12514 7368 12642 7470
rect 10992 7318 11142 7368
rect 11326 7318 12642 7368
rect 10992 7274 12642 7318
rect 13078 7362 13188 7596
rect 13280 7508 14526 7596
rect 13280 7362 13334 7508
rect 13078 7334 13334 7362
rect 13514 7364 14526 7508
rect 14600 7364 14728 7610
rect 13514 7334 14728 7364
rect 13078 7272 14728 7334
rect 18502 7032 18710 7036
rect 15182 7026 18806 7032
rect 15182 7012 18502 7026
rect 15182 6848 15488 7012
rect 15876 7002 18502 7012
rect 15876 6996 16906 7002
rect 15876 6882 16262 6996
rect 16454 6888 16906 6996
rect 17098 6996 18502 7002
rect 17098 6888 17562 6996
rect 16454 6882 17562 6888
rect 17754 6986 18502 6996
rect 17754 6882 18202 6986
rect 15876 6872 18202 6882
rect 18394 6872 18502 6986
rect 15876 6848 18502 6872
rect 15182 6834 18502 6848
rect 18710 6834 18806 7026
rect 15182 6832 18806 6834
rect 18502 6824 18710 6832
rect 6458 6728 11236 6730
rect 6458 6726 11302 6728
rect 6446 6642 11302 6726
rect 6446 6636 9824 6642
rect 6446 6438 7246 6636
rect 6458 6426 7246 6438
rect 7320 6628 9824 6636
rect 7320 6440 8568 6628
rect 8646 6440 9824 6628
rect 7320 6438 9824 6440
rect 9900 6636 11302 6642
rect 9900 6452 11144 6636
rect 11206 6452 11302 6636
rect 9900 6438 11302 6452
rect 7320 6436 11302 6438
rect 7320 6432 11206 6436
rect 7246 6362 7320 6372
rect 6084 6304 6252 6314
rect 11546 6296 11714 6306
rect 6252 6274 8766 6282
rect 6252 6272 8154 6274
rect 6252 6270 7496 6272
rect 6252 6166 6760 6270
rect 7174 6166 7496 6270
rect 7782 6168 8154 6272
rect 8440 6168 8766 6274
rect 9302 6260 9756 6264
rect 9036 6254 11546 6260
rect 9036 6186 9302 6254
rect 9756 6192 10046 6254
rect 10342 6192 10708 6254
rect 11004 6192 11546 6254
rect 9756 6186 11546 6192
rect 9036 6180 11546 6186
rect 9302 6176 9756 6180
rect 7782 6166 8766 6168
rect 6252 6152 8766 6166
rect 6084 6124 6252 6134
rect 11546 6116 11714 6126
rect 6458 5918 8766 6006
rect 6458 5886 7902 5918
rect 6458 5654 6588 5886
rect 6664 5666 7902 5886
rect 7982 5666 8766 5918
rect 6664 5654 8766 5666
rect 6458 5562 8766 5654
rect 9036 5930 11344 6010
rect 9036 5666 9160 5930
rect 9242 5920 11344 5930
rect 9242 5666 10474 5920
rect 9036 5656 10474 5666
rect 10564 5656 11344 5920
rect 9036 5566 11344 5656
rect 6700 5356 6940 5562
rect 9060 5404 9246 5566
rect 6700 5316 7602 5356
rect 6700 5138 6940 5316
rect 6482 5060 7474 5138
rect 6482 4898 6598 5060
rect 6676 4898 7474 5060
rect 6482 4768 7474 4898
rect 7548 4818 7602 5316
rect 8194 5296 9246 5404
rect 8194 5138 8460 5296
rect 7672 5058 8664 5138
rect 7520 4808 7626 4818
rect 7672 4790 7776 5058
rect 7862 4790 8664 5058
rect 7672 4770 8664 4790
rect 7520 4688 7626 4698
rect 6774 4650 7202 4656
rect 7548 4650 7602 4688
rect 7948 4650 8376 4652
rect 6478 4646 8666 4650
rect 6478 4522 6774 4646
rect 7202 4642 8666 4646
rect 7202 4522 7948 4642
rect 6478 4518 7948 4522
rect 8376 4518 8666 4642
rect 6478 4512 8666 4518
rect 7948 4508 8376 4512
rect 6482 4322 7474 4450
rect 6482 4082 7276 4322
rect 7380 4082 7474 4322
rect 6482 3994 7474 4082
rect 7672 4386 8664 4450
rect 7672 4118 8470 4386
rect 8556 4118 8664 4386
rect 7672 3994 8664 4118
rect 8804 4416 8882 5296
rect 8982 5068 9974 5146
rect 8982 4856 9098 5068
rect 9176 5038 9974 5068
rect 9176 4856 9644 5038
rect 8982 4852 9644 4856
rect 9828 4852 9974 5038
rect 8982 4708 9974 4852
rect 10150 5074 11142 5154
rect 10150 4882 10270 5074
rect 10346 5008 11142 5074
rect 10346 4882 10684 5008
rect 10150 4822 10684 4882
rect 10868 4822 11142 5008
rect 10150 4716 11142 4822
rect 11310 5084 14934 5158
rect 11310 4882 11434 5084
rect 11504 5078 14934 5084
rect 11504 5046 14062 5078
rect 11504 4882 12752 5046
rect 11310 4770 12752 4882
rect 11310 4684 11428 4770
rect 11518 4748 12752 4770
rect 12830 4792 14062 5046
rect 14148 5030 14934 5078
rect 14148 4792 14408 5030
rect 12830 4748 14408 4792
rect 11518 4684 14408 4748
rect 11310 4676 14408 4684
rect 14596 4676 14934 5030
rect 10176 4432 10282 4442
rect 8804 4412 9974 4416
rect 8804 4336 9412 4412
rect 9562 4336 9974 4412
rect 10150 4340 10176 4420
rect 8804 4334 9974 4336
rect 8804 4332 8882 4334
rect 6734 3696 7212 3994
rect 6734 3424 6788 3696
rect 7146 3424 7212 3696
rect 6734 3384 7212 3424
rect 7886 3692 8432 3994
rect 7886 3454 7972 3692
rect 8354 3454 8432 3692
rect 8804 3776 8880 4332
rect 10282 4416 11142 4420
rect 10282 4348 10626 4416
rect 10748 4348 11142 4416
rect 11310 4380 14934 4676
rect 15182 4708 18806 5950
rect 10282 4340 11142 4348
rect 15182 4366 15294 4708
rect 15384 4560 18806 4708
rect 15384 4366 16622 4560
rect 15182 4364 16622 4366
rect 16694 4556 18806 4560
rect 16694 4444 17946 4556
rect 16694 4364 17484 4444
rect 10176 4312 10282 4322
rect 15182 4272 17484 4364
rect 17806 4364 17946 4444
rect 18020 4364 18806 4556
rect 17806 4272 18806 4364
rect 17484 4200 17806 4210
rect 8804 3766 8914 3776
rect 8804 3656 8808 3766
rect 8804 3646 8914 3656
rect 8982 3664 9974 3890
rect 8804 3642 8880 3646
rect 7886 3396 8432 3454
rect 8982 3482 9770 3664
rect 9856 3482 9974 3664
rect 8982 3402 9974 3482
rect 10150 3692 11142 3896
rect 14610 3846 14932 3856
rect 10150 3492 10936 3692
rect 11026 3492 11142 3692
rect 11310 3790 14610 3802
rect 11310 3782 14300 3790
rect 11310 3778 12366 3782
rect 11310 3652 11590 3778
rect 11748 3654 11828 3778
rect 11980 3668 12366 3778
rect 12558 3668 13050 3782
rect 13242 3774 14300 3782
rect 13242 3668 13678 3774
rect 11980 3660 13678 3668
rect 13870 3676 14300 3774
rect 14492 3676 14610 3790
rect 13870 3660 14610 3676
rect 11980 3654 14610 3660
rect 11748 3652 14610 3654
rect 11310 3642 14610 3652
rect 14932 3642 14934 3802
rect 14610 3602 14932 3612
rect 10150 3408 11142 3492
rect 9308 3290 9644 3402
rect 9308 3136 9340 3290
rect 9610 3136 9644 3290
rect 9308 3118 9644 3136
rect 10412 3258 10878 3408
rect 10412 3080 10484 3258
rect 10818 3080 10878 3258
rect 10412 3040 10878 3080
rect 11310 2182 14934 2728
rect 16646 2568 16858 2596
rect 16646 2384 16692 2568
rect 16844 2384 16858 2568
rect 16646 2366 16858 2384
rect 11310 2126 14730 2182
rect 11310 2104 13408 2126
rect 11310 1892 12094 2104
rect 12168 1896 13408 2104
rect 13488 1898 14730 2126
rect 14818 1898 14934 2182
rect 13488 1896 14934 1898
rect 12168 1892 14934 1896
rect 11310 1814 14934 1892
rect 12886 1644 13352 1814
rect 12886 1370 12950 1644
rect 13302 1370 13352 1644
rect 12886 1332 13352 1370
<< via2 >>
rect 11142 7368 11192 7504
rect 11192 7368 11326 7504
rect 11142 7318 11326 7368
rect 13334 7334 13514 7508
rect 18502 6834 18710 7026
rect 7520 4698 7626 4808
rect 9644 4852 9828 5038
rect 10684 4822 10868 5008
rect 14408 4676 14596 5030
rect 10176 4322 10282 4432
rect 17484 4210 17806 4444
rect 8808 3656 8914 3766
rect 11590 3652 11748 3778
rect 14610 3612 14932 3846
rect 16692 2384 16844 2568
<< metal3 >>
rect 9584 7504 11388 7562
rect 9584 7318 11142 7504
rect 11326 7318 11388 7504
rect 9584 7282 11388 7318
rect 13310 7508 13556 7540
rect 13310 7334 13334 7508
rect 13514 7334 13556 7508
rect 9098 4856 9176 5068
rect 9594 5038 9880 7282
rect 13310 5042 13556 7334
rect 18972 7042 19272 7046
rect 18496 7031 19276 7042
rect 18492 7026 19276 7031
rect 18492 6834 18502 7026
rect 18710 6834 19276 7026
rect 18492 6829 19276 6834
rect 18496 6820 19276 6829
rect 9594 4852 9644 5038
rect 9828 4852 9880 5038
rect 7510 4808 7638 4820
rect 9594 4814 9880 4852
rect 10328 5008 13556 5042
rect 10328 4822 10684 5008
rect 10868 4822 13556 5008
rect 7510 4698 7520 4808
rect 7626 4698 7638 4808
rect 10328 4790 13556 4822
rect 14360 5030 14638 5086
rect 7510 4446 7638 4698
rect 14360 4676 14408 5030
rect 14596 4676 14638 5030
rect 14360 4604 14638 4676
rect 7510 4432 10340 4446
rect 7510 4322 10176 4432
rect 10282 4322 10340 4432
rect 7510 4308 10340 4322
rect 17442 4444 17848 4478
rect 17442 4226 17484 4444
rect 17438 4210 17484 4226
rect 17806 4226 17848 4444
rect 17806 4210 17850 4226
rect 17438 4142 17850 4210
rect 17434 3916 17856 4142
rect 14600 3846 16048 3854
rect 8804 3778 11766 3786
rect 8804 3771 11590 3778
rect 8798 3766 11590 3771
rect 8798 3656 8808 3766
rect 8914 3656 11590 3766
rect 8798 3652 11590 3656
rect 11748 3652 11766 3778
rect 8798 3651 11766 3652
rect 8804 3642 11766 3651
rect 14600 3612 14610 3846
rect 14932 3816 16048 3846
rect 14932 3612 15810 3816
rect 16024 3612 16048 3816
rect 17434 3794 17472 3916
rect 17830 3794 17856 3916
rect 17434 3784 17856 3794
rect 14600 3586 16048 3612
rect 15552 3584 16048 3586
rect 18972 3316 19272 6820
rect 18972 3286 19288 3316
rect 18972 3244 18992 3286
rect 18974 3046 18992 3244
rect 19258 3046 19288 3286
rect 18974 3008 19288 3046
rect 16614 2568 16858 2614
rect 16614 2384 16692 2568
rect 16844 2384 16858 2568
rect 16614 2342 16858 2384
<< via3 >>
rect 14408 4676 14596 5030
rect 15810 3612 16024 3816
rect 17472 3794 17830 3916
rect 18992 3046 19258 3286
rect 16692 2384 16844 2568
<< metal4 >>
rect 14312 5030 15330 5088
rect 14312 4676 14408 5030
rect 14596 4676 15330 5030
rect 14312 4594 15330 4676
rect 15046 2690 15328 4594
rect 17434 3916 17856 3930
rect 15796 3816 16048 3854
rect 15796 3612 15810 3816
rect 16024 3612 16048 3816
rect 17434 3794 17472 3916
rect 17830 3794 17856 3916
rect 15796 2932 16048 3612
rect 16688 3562 17102 3670
rect 17434 3572 17856 3794
rect 16688 2704 16866 3562
rect 17026 3286 19276 3326
rect 17026 3046 18992 3286
rect 19258 3046 19276 3286
rect 17026 3008 19276 3046
rect 15046 2310 15996 2690
rect 16084 2568 16866 2704
rect 16084 2384 16692 2568
rect 16844 2384 16866 2568
rect 16084 2380 16866 2384
rect 15046 2308 15328 2310
rect 16084 2292 16858 2380
use sky130_fd_pr__cap_mim_m3_1_ZYFHHD  XC1 ~/ColRO/mag
timestamp 1695378092
transform 0 -1 17434 1 0 3284
box -386 -440 386 440
use sky130_fd_pr__cap_mim_m3_1_ZYFHHD  XC2
timestamp 1695378092
transform 0 -1 15894 1 0 2646
box -386 -440 386 440
use sky130_fd_pr__nfet_01v8_lvt_7233E2  XM2 ~/ColRO/mag
timestamp 1695441144
transform 1 0 9478 0 1 4274
box -496 -1010 496 1010
use sky130_fd_pr__pfet_01v8_lvt_CEAZV5  XM3 ~/ColRO/mag
timestamp 1695440875
transform 1 0 11817 0 1 7855
box -825 -719 825 719
use sky130_fd_pr__pfet_01v8_lvt_CEAZV5  XM4
timestamp 1695440875
transform 1 0 13903 0 1 7853
box -825 -719 825 719
use sky130_fd_pr__nfet_01v8_lvt_7233E2  XM5
timestamp 1695441144
transform 1 0 10646 0 1 4282
box -496 -1010 496 1010
use sky130_fd_pr__pfet_01v8_lvt_LEXMNV  XM10 ~/ColRO/mag
timestamp 1695441144
transform 1 0 16994 0 1 6355
box -1812 -2219 1812 2219
use sky130_fd_pr__pfet_01v8_lvt_CEE7V5  XM14 ~/ColRO/mag
timestamp 1696133064
transform 1 0 7612 0 1 6143
box -1154 -719 1154 719
use sky130_fd_pr__pfet_01v8_lvt_CEE7V5  XM15
timestamp 1696133064
transform 1 0 10190 0 1 6149
box -1154 -719 1154 719
use sky130_fd_pr__nfet_01v8_lvt_HZEGLD  XM17 ~/ColRO/mag
timestamp 1695441144
transform 1 0 13122 0 1 3486
box -1812 -1810 1812 1810
use sky130_fd_pr__nfet_01v8_lvt_RFVHWA  XM19 ~/ColRO/mag
timestamp 1695441144
transform 1 0 6978 0 1 4566
box -496 -710 496 710
use sky130_fd_pr__nfet_01v8_lvt_RFVHWA  XM20
timestamp 1695441144
transform 1 0 8168 0 1 4566
box -496 -710 496 710
use sky130_fd_pr__pfet_01v8_lvt_8WRJS5  XM26 ~/ColRO/mag
timestamp 1695378092
transform 1 0 8963 0 1 8101
box -1483 -469 1483 469
<< labels >>
flabel metal1 7118 7978 7318 8178 0 FreeSans 256 0 0 0 opbias
port 0 nsew
flabel metal1 6068 6120 6268 6320 0 FreeSans 256 0 0 0 inn
port 2 nsew
flabel metal1 11534 6114 11734 6314 0 FreeSans 256 0 0 0 inp
port 1 nsew
flabel metal1 16658 2376 16858 2576 0 FreeSans 256 0 0 0 out
port 3 nsew
rlabel locali 6276 1244 15318 1756 1 GROUND
port 5 nsew
rlabel locali 7334 8482 18966 9014 1 VDD
port 4 nsew
<< end >>
