magic
tech sky130A
timestamp 1695195131
<< pwell >>
rect -198 -2605 198 2605
<< nmoslvt >>
rect -100 -2500 100 2500
<< ndiff >>
rect -129 2494 -100 2500
rect -129 -2494 -123 2494
rect -106 -2494 -100 2494
rect -129 -2500 -100 -2494
rect 100 2494 129 2500
rect 100 -2494 106 2494
rect 123 -2494 129 2494
rect 100 -2500 129 -2494
<< ndiffc >>
rect -123 -2494 -106 2494
rect 106 -2494 123 2494
<< psubdiff >>
rect -180 2570 -132 2587
rect 132 2570 180 2587
rect -180 2539 -163 2570
rect 163 2539 180 2570
rect -180 -2570 -163 -2539
rect 163 -2570 180 -2539
rect -180 -2587 -132 -2570
rect 132 -2587 180 -2570
<< psubdiffcont >>
rect -132 2570 132 2587
rect -180 -2539 -163 2539
rect 163 -2539 180 2539
rect -132 -2587 132 -2570
<< poly >>
rect -100 2536 100 2544
rect -100 2519 -92 2536
rect 92 2519 100 2536
rect -100 2500 100 2519
rect -100 -2519 100 -2500
rect -100 -2536 -92 -2519
rect 92 -2536 100 -2519
rect -100 -2544 100 -2536
<< polycont >>
rect -92 2519 92 2536
rect -92 -2536 92 -2519
<< locali >>
rect -180 2570 -132 2587
rect 132 2570 180 2587
rect -180 2539 -163 2570
rect 163 2539 180 2570
rect -100 2519 -92 2536
rect 92 2519 100 2536
rect -123 2494 -106 2502
rect -123 -2502 -106 -2494
rect 106 2494 123 2502
rect 106 -2502 123 -2494
rect -100 -2536 -92 -2519
rect 92 -2536 100 -2519
rect -180 -2570 -163 -2539
rect 163 -2570 180 -2539
rect -180 -2587 -132 -2570
rect 132 -2587 180 -2570
<< viali >>
rect -92 2519 92 2536
rect -123 -2494 -106 2494
rect 106 -2494 123 2494
rect -92 -2536 92 -2519
<< metal1 >>
rect -98 2536 98 2539
rect -98 2519 -92 2536
rect 92 2519 98 2536
rect -98 2516 98 2519
rect -126 2494 -103 2500
rect -126 -2494 -123 2494
rect -106 -2494 -103 2494
rect -126 -2500 -103 -2494
rect 103 2494 126 2500
rect 103 -2494 106 2494
rect 123 -2494 126 2494
rect 103 -2500 126 -2494
rect -98 -2519 98 -2516
rect -98 -2536 -92 -2519
rect 92 -2536 98 -2519
rect -98 -2539 98 -2536
<< properties >>
string FIXED_BBOX -171 -2578 171 2578
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 50.0 l 2.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
