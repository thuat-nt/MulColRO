magic
tech sky130A
magscale 1 2
timestamp 1694848836
<< nwell >>
rect -1812 -399 1812 399
<< pmoslvt >>
rect -1616 -180 -1016 180
rect -958 -180 -358 180
rect -300 -180 300 180
rect 358 -180 958 180
rect 1016 -180 1616 180
<< pdiff >>
rect -1674 168 -1616 180
rect -1674 -168 -1662 168
rect -1628 -168 -1616 168
rect -1674 -180 -1616 -168
rect -1016 168 -958 180
rect -1016 -168 -1004 168
rect -970 -168 -958 168
rect -1016 -180 -958 -168
rect -358 168 -300 180
rect -358 -168 -346 168
rect -312 -168 -300 168
rect -358 -180 -300 -168
rect 300 168 358 180
rect 300 -168 312 168
rect 346 -168 358 168
rect 300 -180 358 -168
rect 958 168 1016 180
rect 958 -168 970 168
rect 1004 -168 1016 168
rect 958 -180 1016 -168
rect 1616 168 1674 180
rect 1616 -168 1628 168
rect 1662 -168 1674 168
rect 1616 -180 1674 -168
<< pdiffc >>
rect -1662 -168 -1628 168
rect -1004 -168 -970 168
rect -346 -168 -312 168
rect 312 -168 346 168
rect 970 -168 1004 168
rect 1628 -168 1662 168
<< nsubdiff >>
rect -1776 329 -1680 363
rect 1680 329 1776 363
rect -1776 267 -1742 329
rect 1742 267 1776 329
rect -1776 -329 -1742 -267
rect 1742 -329 1776 -267
rect -1776 -363 -1680 -329
rect 1680 -363 1776 -329
<< nsubdiffcont >>
rect -1680 329 1680 363
rect -1776 -267 -1742 267
rect 1742 -267 1776 267
rect -1680 -363 1680 -329
<< poly >>
rect -1616 261 -1016 277
rect -1616 227 -1600 261
rect -1032 227 -1016 261
rect -1616 180 -1016 227
rect -958 261 -358 277
rect -958 227 -942 261
rect -374 227 -358 261
rect -958 180 -358 227
rect -300 261 300 277
rect -300 227 -284 261
rect 284 227 300 261
rect -300 180 300 227
rect 358 261 958 277
rect 358 227 374 261
rect 942 227 958 261
rect 358 180 958 227
rect 1016 261 1616 277
rect 1016 227 1032 261
rect 1600 227 1616 261
rect 1016 180 1616 227
rect -1616 -227 -1016 -180
rect -1616 -261 -1600 -227
rect -1032 -261 -1016 -227
rect -1616 -277 -1016 -261
rect -958 -227 -358 -180
rect -958 -261 -942 -227
rect -374 -261 -358 -227
rect -958 -277 -358 -261
rect -300 -227 300 -180
rect -300 -261 -284 -227
rect 284 -261 300 -227
rect -300 -277 300 -261
rect 358 -227 958 -180
rect 358 -261 374 -227
rect 942 -261 958 -227
rect 358 -277 958 -261
rect 1016 -227 1616 -180
rect 1016 -261 1032 -227
rect 1600 -261 1616 -227
rect 1016 -277 1616 -261
<< polycont >>
rect -1600 227 -1032 261
rect -942 227 -374 261
rect -284 227 284 261
rect 374 227 942 261
rect 1032 227 1600 261
rect -1600 -261 -1032 -227
rect -942 -261 -374 -227
rect -284 -261 284 -227
rect 374 -261 942 -227
rect 1032 -261 1600 -227
<< locali >>
rect -1776 329 -1680 363
rect 1680 329 1776 363
rect -1776 267 -1742 329
rect 1742 267 1776 329
rect -1616 227 -1600 261
rect -1032 227 -1016 261
rect -958 227 -942 261
rect -374 227 -358 261
rect -300 227 -284 261
rect 284 227 300 261
rect 358 227 374 261
rect 942 227 958 261
rect 1016 227 1032 261
rect 1600 227 1616 261
rect -1662 168 -1628 184
rect -1662 -184 -1628 -168
rect -1004 168 -970 184
rect -1004 -184 -970 -168
rect -346 168 -312 184
rect -346 -184 -312 -168
rect 312 168 346 184
rect 312 -184 346 -168
rect 970 168 1004 184
rect 970 -184 1004 -168
rect 1628 168 1662 184
rect 1628 -184 1662 -168
rect -1616 -261 -1600 -227
rect -1032 -261 -1016 -227
rect -958 -261 -942 -227
rect -374 -261 -358 -227
rect -300 -261 -284 -227
rect 284 -261 300 -227
rect 358 -261 374 -227
rect 942 -261 958 -227
rect 1016 -261 1032 -227
rect 1600 -261 1616 -227
rect -1776 -329 -1742 -267
rect 1742 -329 1776 -267
rect -1776 -363 -1680 -329
rect 1680 -363 1776 -329
<< viali >>
rect -1600 227 -1032 261
rect -942 227 -374 261
rect -284 227 284 261
rect 374 227 942 261
rect 1032 227 1600 261
rect -1662 -168 -1628 168
rect -1004 -168 -970 168
rect -346 -168 -312 168
rect 312 -168 346 168
rect 970 -168 1004 168
rect 1628 -168 1662 168
rect -1600 -261 -1032 -227
rect -942 -261 -374 -227
rect -284 -261 284 -227
rect 374 -261 942 -227
rect 1032 -261 1600 -227
<< metal1 >>
rect -1612 261 -1020 267
rect -1612 227 -1600 261
rect -1032 227 -1020 261
rect -1612 221 -1020 227
rect -954 261 -362 267
rect -954 227 -942 261
rect -374 227 -362 261
rect -954 221 -362 227
rect -296 261 296 267
rect -296 227 -284 261
rect 284 227 296 261
rect -296 221 296 227
rect 362 261 954 267
rect 362 227 374 261
rect 942 227 954 261
rect 362 221 954 227
rect 1020 261 1612 267
rect 1020 227 1032 261
rect 1600 227 1612 261
rect 1020 221 1612 227
rect -1668 168 -1622 180
rect -1668 -168 -1662 168
rect -1628 -168 -1622 168
rect -1668 -180 -1622 -168
rect -1010 168 -964 180
rect -1010 -168 -1004 168
rect -970 -168 -964 168
rect -1010 -180 -964 -168
rect -352 168 -306 180
rect -352 -168 -346 168
rect -312 -168 -306 168
rect -352 -180 -306 -168
rect 306 168 352 180
rect 306 -168 312 168
rect 346 -168 352 168
rect 306 -180 352 -168
rect 964 168 1010 180
rect 964 -168 970 168
rect 1004 -168 1010 168
rect 964 -180 1010 -168
rect 1622 168 1668 180
rect 1622 -168 1628 168
rect 1662 -168 1668 168
rect 1622 -180 1668 -168
rect -1612 -227 -1020 -221
rect -1612 -261 -1600 -227
rect -1032 -261 -1020 -227
rect -1612 -267 -1020 -261
rect -954 -227 -362 -221
rect -954 -261 -942 -227
rect -374 -261 -362 -227
rect -954 -267 -362 -261
rect -296 -227 296 -221
rect -296 -261 -284 -227
rect 284 -261 296 -227
rect -296 -267 296 -261
rect 362 -227 954 -221
rect 362 -261 374 -227
rect 942 -261 954 -227
rect 362 -267 954 -261
rect 1020 -227 1612 -221
rect 1020 -261 1032 -227
rect 1600 -261 1612 -227
rect 1020 -267 1612 -261
<< properties >>
string FIXED_BBOX -1759 -346 1759 346
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 1.8 l 3.0 m 1 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
