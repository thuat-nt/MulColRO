magic
tech sky130A
magscale 1 2
timestamp 1695461801
<< metal3 >>
rect -56 58 56 115
rect -56 -115 56 -58
<< rmetal3 >>
rect -56 -58 56 58
<< properties >>
string gencell sky130_fd_pr__res_generic_m3
string library sky130
string parameters w 0.56 l 0.58 m 1 nx 1 wmin 0.30 lmin 0.30 rho 0.047 val 48.678m dummy 0 dw 0.0 term 0.0 roverlap 0
<< end >>
