magic
tech sky130A
magscale 1 2
timestamp 1694848836
<< nwell >>
rect -1154 -6852 1154 6852
<< pmoslvt >>
rect -958 -6633 -358 6633
rect -300 -6633 300 6633
rect 358 -6633 958 6633
<< pdiff >>
rect -1016 6621 -958 6633
rect -1016 -6621 -1004 6621
rect -970 -6621 -958 6621
rect -1016 -6633 -958 -6621
rect -358 6621 -300 6633
rect -358 -6621 -346 6621
rect -312 -6621 -300 6621
rect -358 -6633 -300 -6621
rect 300 6621 358 6633
rect 300 -6621 312 6621
rect 346 -6621 358 6621
rect 300 -6633 358 -6621
rect 958 6621 1016 6633
rect 958 -6621 970 6621
rect 1004 -6621 1016 6621
rect 958 -6633 1016 -6621
<< pdiffc >>
rect -1004 -6621 -970 6621
rect -346 -6621 -312 6621
rect 312 -6621 346 6621
rect 970 -6621 1004 6621
<< nsubdiff >>
rect -1118 6782 -1022 6816
rect 1022 6782 1118 6816
rect -1118 6720 -1084 6782
rect 1084 6720 1118 6782
rect -1118 -6782 -1084 -6720
rect 1084 -6782 1118 -6720
rect -1118 -6816 -1022 -6782
rect 1022 -6816 1118 -6782
<< nsubdiffcont >>
rect -1022 6782 1022 6816
rect -1118 -6720 -1084 6720
rect 1084 -6720 1118 6720
rect -1022 -6816 1022 -6782
<< poly >>
rect -958 6714 -358 6730
rect -958 6680 -942 6714
rect -374 6680 -358 6714
rect -958 6633 -358 6680
rect -300 6714 300 6730
rect -300 6680 -284 6714
rect 284 6680 300 6714
rect -300 6633 300 6680
rect 358 6714 958 6730
rect 358 6680 374 6714
rect 942 6680 958 6714
rect 358 6633 958 6680
rect -958 -6680 -358 -6633
rect -958 -6714 -942 -6680
rect -374 -6714 -358 -6680
rect -958 -6730 -358 -6714
rect -300 -6680 300 -6633
rect -300 -6714 -284 -6680
rect 284 -6714 300 -6680
rect -300 -6730 300 -6714
rect 358 -6680 958 -6633
rect 358 -6714 374 -6680
rect 942 -6714 958 -6680
rect 358 -6730 958 -6714
<< polycont >>
rect -942 6680 -374 6714
rect -284 6680 284 6714
rect 374 6680 942 6714
rect -942 -6714 -374 -6680
rect -284 -6714 284 -6680
rect 374 -6714 942 -6680
<< locali >>
rect -1118 6782 -1022 6816
rect 1022 6782 1118 6816
rect -1118 6720 -1084 6782
rect 1084 6720 1118 6782
rect -958 6680 -942 6714
rect -374 6680 -358 6714
rect -300 6680 -284 6714
rect 284 6680 300 6714
rect 358 6680 374 6714
rect 942 6680 958 6714
rect -1004 6621 -970 6637
rect -1004 -6637 -970 -6621
rect -346 6621 -312 6637
rect -346 -6637 -312 -6621
rect 312 6621 346 6637
rect 312 -6637 346 -6621
rect 970 6621 1004 6637
rect 970 -6637 1004 -6621
rect -958 -6714 -942 -6680
rect -374 -6714 -358 -6680
rect -300 -6714 -284 -6680
rect 284 -6714 300 -6680
rect 358 -6714 374 -6680
rect 942 -6714 958 -6680
rect -1118 -6782 -1084 -6720
rect 1084 -6782 1118 -6720
rect -1118 -6816 -1022 -6782
rect 1022 -6816 1118 -6782
<< viali >>
rect -942 6680 -374 6714
rect -284 6680 284 6714
rect 374 6680 942 6714
rect -1004 -6621 -970 6621
rect -346 -6621 -312 6621
rect 312 -6621 346 6621
rect 970 -6621 1004 6621
rect -942 -6714 -374 -6680
rect -284 -6714 284 -6680
rect 374 -6714 942 -6680
<< metal1 >>
rect -954 6714 -362 6720
rect -954 6680 -942 6714
rect -374 6680 -362 6714
rect -954 6674 -362 6680
rect -296 6714 296 6720
rect -296 6680 -284 6714
rect 284 6680 296 6714
rect -296 6674 296 6680
rect 362 6714 954 6720
rect 362 6680 374 6714
rect 942 6680 954 6714
rect 362 6674 954 6680
rect -1010 6621 -964 6633
rect -1010 -6621 -1004 6621
rect -970 -6621 -964 6621
rect -1010 -6633 -964 -6621
rect -352 6621 -306 6633
rect -352 -6621 -346 6621
rect -312 -6621 -306 6621
rect -352 -6633 -306 -6621
rect 306 6621 352 6633
rect 306 -6621 312 6621
rect 346 -6621 352 6621
rect 306 -6633 352 -6621
rect 964 6621 1010 6633
rect 964 -6621 970 6621
rect 1004 -6621 1010 6621
rect 964 -6633 1010 -6621
rect -954 -6680 -362 -6674
rect -954 -6714 -942 -6680
rect -374 -6714 -362 -6680
rect -954 -6720 -362 -6714
rect -296 -6680 296 -6674
rect -296 -6714 -284 -6680
rect 284 -6714 296 -6680
rect -296 -6720 296 -6714
rect 362 -6680 954 -6674
rect 362 -6714 374 -6680
rect 942 -6714 954 -6680
rect 362 -6720 954 -6714
<< properties >>
string FIXED_BBOX -1101 -6799 1101 6799
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 66.33333333333333 l 3.0 m 1 nf 3 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
